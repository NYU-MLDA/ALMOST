//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G85gat), .ZN(new_n205_));
  INV_X1    g004(.A(G92gat), .ZN(new_n206_));
  NOR3_X1   g005(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT9), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G85gat), .B(G92gat), .Z(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT9), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT10), .B(G99gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n208_), .B(new_n210_), .C1(G106gat), .C2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT7), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n204_), .B1(new_n216_), .B2(KEYINPUT64), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(KEYINPUT64), .B2(new_n216_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n213_), .B1(new_n218_), .B2(new_n209_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n213_), .B(new_n209_), .C1(new_n216_), .C2(new_n204_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n212_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G43gat), .B(G50gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(G29gat), .B(G36gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT15), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n227_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n212_), .B(new_n231_), .C1(new_n221_), .C2(new_n223_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G232gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT34), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT35), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT68), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n230_), .A2(new_n232_), .A3(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n235_), .A2(new_n236_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n239_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n230_), .A2(new_n241_), .A3(new_n232_), .A4(new_n237_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G190gat), .B(G218gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G134gat), .B(G162gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT67), .B(KEYINPUT36), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n243_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n240_), .A2(KEYINPUT69), .A3(new_n242_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n246_), .B(KEYINPUT36), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n251_), .B1(new_n243_), .B2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n248_), .B1(new_n249_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n248_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT37), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n251_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n257_));
  OAI22_X1  g056(.A1(new_n254_), .A2(KEYINPUT37), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT73), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G57gat), .B(G64gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT11), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT66), .ZN(new_n262_));
  XOR2_X1   g061(.A(G71gat), .B(G78gat), .Z(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(KEYINPUT11), .B2(new_n260_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n262_), .B(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G231gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT71), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n265_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G1gat), .B(G8gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT70), .ZN(new_n270_));
  INV_X1    g069(.A(G15gat), .ZN(new_n271_));
  INV_X1    g070(.A(G22gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G15gat), .A2(G22gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G1gat), .A2(G8gat), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n273_), .A2(new_n274_), .B1(KEYINPUT14), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n270_), .B(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n268_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n268_), .A2(new_n277_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G127gat), .B(G155gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G183gat), .B(G211gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT17), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n278_), .A2(new_n279_), .A3(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n278_), .A2(new_n279_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT17), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n259_), .B(new_n286_), .C1(new_n287_), .C2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(KEYINPUT73), .A3(new_n285_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n258_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT74), .ZN(new_n295_));
  INV_X1    g094(.A(new_n265_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n224_), .A2(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n212_), .B(new_n265_), .C1(new_n221_), .C2(new_n223_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G230gat), .A2(G233gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(KEYINPUT12), .A3(new_n298_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT12), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n224_), .A2(new_n304_), .A3(new_n296_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n300_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G120gat), .B(G148gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT5), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G176gat), .B(G204gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n302_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n300_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n314_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n311_), .B1(new_n301_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT13), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n313_), .A2(KEYINPUT13), .A3(new_n316_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G127gat), .B(G134gat), .Z(new_n322_));
  XOR2_X1   g121(.A(G113gat), .B(G120gat), .Z(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT84), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT83), .B1(new_n325_), .B2(KEYINPUT31), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(KEYINPUT31), .B2(new_n325_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(G15gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT30), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n327_), .B(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT77), .A2(G169gat), .A3(G176gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT81), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT22), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G169gat), .ZN(new_n338_));
  INV_X1    g137(.A(G169gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT22), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n336_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n336_), .B1(new_n339_), .B2(KEYINPUT22), .ZN(new_n342_));
  INV_X1    g141(.A(G176gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n335_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT82), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT82), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n347_), .B(new_n335_), .C1(new_n341_), .C2(new_n344_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(G183gat), .B2(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n357_), .A2(KEYINPUT78), .A3(new_n360_), .A4(new_n332_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT25), .B(G183gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT26), .B(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT78), .B1(new_n335_), .B2(new_n357_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n355_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n360_), .A2(new_n332_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n356_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n370_), .A2(KEYINPUT79), .A3(new_n364_), .A4(new_n361_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT24), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n339_), .A3(new_n343_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT80), .B1(new_n352_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n378_));
  AND4_X1   g177(.A1(KEYINPUT80), .A2(new_n373_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n367_), .A2(new_n371_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n354_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G71gat), .B(G99gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G43gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n382_), .B(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n331_), .B(new_n385_), .Z(new_n386_));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G85gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT0), .B(G57gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(new_n389_), .Z(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT85), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(G141gat), .A3(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n395_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G141gat), .ZN(new_n400_));
  INV_X1    g199(.A(G148gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT3), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(G141gat), .B2(G148gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G155gat), .A2(G162gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G155gat), .A2(G162gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT86), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT86), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(G155gat), .A3(G162gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT88), .B1(new_n407_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(KEYINPUT88), .A3(new_n413_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n410_), .A2(new_n412_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n408_), .B1(new_n417_), .B2(KEYINPUT1), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT1), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n410_), .A2(new_n412_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n410_), .A2(new_n412_), .A3(KEYINPUT87), .A4(new_n419_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n418_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n395_), .A2(new_n397_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n415_), .A2(new_n416_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n324_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n393_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n426_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n407_), .A2(KEYINPUT88), .A3(new_n413_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n431_), .B(KEYINPUT97), .C1(new_n414_), .C2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n324_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n415_), .A2(new_n416_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n436_), .A2(KEYINPUT97), .A3(new_n431_), .A4(new_n324_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n430_), .B1(new_n438_), .B2(KEYINPUT4), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n393_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n391_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n392_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n428_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n442_), .B(new_n390_), .C1(new_n443_), .C2(new_n430_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n386_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(G228gat), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT29), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n427_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G197gat), .A2(G204gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT92), .B(G197gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n455_), .B2(G204gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G211gat), .B(G218gat), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT21), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n455_), .A2(G204gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n458_), .B1(G197gat), .B2(G204gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n457_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n456_), .A2(KEYINPUT21), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n460_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT91), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n451_), .B1(new_n453_), .B2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n466_), .A2(KEYINPUT91), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n469_), .B(new_n450_), .C1(new_n452_), .C2(new_n427_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G78gat), .B(G106gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n468_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT89), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n436_), .A2(new_n431_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(KEYINPUT29), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n427_), .A2(KEYINPUT89), .A3(new_n452_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G22gat), .B(G50gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT28), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n478_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n475_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n468_), .A2(new_n470_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n471_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n473_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n484_), .A2(new_n487_), .A3(KEYINPUT93), .A4(new_n473_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n363_), .B(KEYINPUT94), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n362_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n352_), .A2(new_n373_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n496_), .B1(new_n358_), .B2(new_n357_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n338_), .A2(new_n340_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n369_), .B1(new_n498_), .B2(new_n343_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n495_), .A2(new_n497_), .B1(new_n353_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n493_), .B1(new_n501_), .B2(new_n466_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G226gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT19), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n465_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n457_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n506_), .A2(new_n508_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n354_), .A2(new_n381_), .A3(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n502_), .A2(new_n505_), .A3(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT20), .B1(new_n501_), .B2(new_n466_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT95), .ZN(new_n513_));
  INV_X1    g312(.A(new_n353_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n514_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n371_), .A2(new_n380_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n516_), .B2(new_n367_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n513_), .B1(new_n517_), .B2(new_n509_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n382_), .A2(KEYINPUT95), .A3(new_n466_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n512_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n511_), .B1(new_n520_), .B2(new_n505_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G8gat), .B(G36gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT18), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G64gat), .B(G92gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT102), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n521_), .A2(new_n526_), .ZN(new_n527_));
  AOI211_X1 g326(.A(new_n493_), .B(new_n504_), .C1(new_n500_), .C2(new_n509_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n517_), .A2(new_n513_), .A3(new_n509_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT95), .B1(new_n382_), .B2(new_n466_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n502_), .A2(new_n510_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n504_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n533_), .A3(new_n525_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n527_), .A2(KEYINPUT27), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT27), .ZN(new_n536_));
  OAI211_X1 g335(.A(KEYINPUT20), .B(new_n505_), .C1(new_n501_), .C2(new_n466_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n505_), .B1(new_n502_), .B2(new_n510_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n525_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n525_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n536_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n535_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n492_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n446_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n445_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n489_), .A2(new_n547_), .A3(new_n490_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n525_), .A2(KEYINPUT32), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n521_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n531_), .A2(new_n533_), .A3(new_n550_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n445_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT101), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n552_), .A2(new_n445_), .A3(new_n553_), .A4(KEYINPUT101), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT33), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n391_), .A2(new_n558_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n442_), .B(new_n559_), .C1(new_n443_), .C2(new_n430_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT98), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n438_), .A2(KEYINPUT4), .ZN(new_n562_));
  INV_X1    g361(.A(new_n430_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT98), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(new_n442_), .A4(new_n559_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n438_), .A2(new_n393_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n391_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n392_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n443_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT100), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n390_), .B1(new_n438_), .B2(new_n393_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT100), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n573_), .B(new_n574_), .C1(new_n443_), .C2(new_n570_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n444_), .A2(KEYINPUT99), .A3(new_n558_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT99), .B1(new_n444_), .B2(new_n558_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n567_), .B(new_n576_), .C1(new_n577_), .C2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT96), .B1(new_n541_), .B2(new_n542_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n540_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT96), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n534_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n556_), .B(new_n557_), .C1(new_n579_), .C2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n549_), .B1(new_n585_), .B2(new_n491_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n386_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n546_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n277_), .B(new_n231_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT75), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n277_), .A2(new_n231_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n277_), .A2(new_n231_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(KEYINPUT75), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n589_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT76), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n228_), .B2(new_n277_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n589_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT76), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n598_), .B1(new_n596_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G113gat), .B(G141gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G169gat), .B(G197gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n605_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n598_), .B(new_n607_), .C1(new_n596_), .C2(new_n601_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n588_), .A2(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n295_), .A2(new_n321_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(G1gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n445_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT38), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n253_), .A2(new_n249_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n255_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n588_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n617_), .A2(KEYINPUT103), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(KEYINPUT103), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n321_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n609_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(new_n293_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n445_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n614_), .B1(new_n612_), .B2(new_n626_), .ZN(G1324gat));
  INV_X1    g426(.A(G8gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n611_), .A2(new_n628_), .A3(new_n544_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n544_), .B(new_n623_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n630_), .A2(new_n631_), .A3(G8gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n630_), .B2(G8gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(G1325gat));
  NAND3_X1  g435(.A1(new_n611_), .A2(new_n271_), .A3(new_n587_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n624_), .A2(new_n587_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n638_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT41), .B1(new_n638_), .B2(G15gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n637_), .B1(new_n639_), .B2(new_n640_), .ZN(G1326gat));
  NAND2_X1  g440(.A1(new_n492_), .A2(new_n272_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT104), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n611_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n624_), .A2(new_n492_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(G22gat), .ZN(new_n647_));
  AOI211_X1 g446(.A(KEYINPUT42), .B(new_n272_), .C1(new_n624_), .C2(new_n492_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n644_), .B1(new_n647_), .B2(new_n648_), .ZN(G1327gat));
  NOR2_X1   g448(.A1(new_n616_), .A2(new_n292_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n621_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT106), .B1(new_n610_), .B2(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n321_), .A2(new_n616_), .A3(new_n292_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n653_), .A2(new_n654_), .A3(new_n588_), .A4(new_n609_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n547_), .A2(G29gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n652_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n622_), .A2(new_n292_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n588_), .A2(new_n659_), .A3(new_n258_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n588_), .B2(new_n258_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n658_), .B(KEYINPUT44), .C1(new_n660_), .C2(new_n661_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n445_), .A3(new_n665_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n666_), .A2(KEYINPUT105), .A3(G29gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT105), .B1(new_n666_), .B2(G29gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n657_), .B1(new_n667_), .B2(new_n668_), .ZN(G1328gat));
  NAND3_X1  g468(.A1(new_n664_), .A2(new_n544_), .A3(new_n665_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G36gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n544_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(G36gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n652_), .A2(new_n655_), .A3(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT45), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT46), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT46), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT107), .B(new_n679_), .C1(new_n671_), .C2(new_n675_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1329gat));
  NAND4_X1  g480(.A1(new_n664_), .A2(G43gat), .A3(new_n587_), .A4(new_n665_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n652_), .A2(new_n587_), .A3(new_n655_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT108), .B(G43gat), .Z(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(G1330gat));
  NAND4_X1  g486(.A1(new_n664_), .A2(G50gat), .A3(new_n492_), .A4(new_n665_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n652_), .A2(new_n492_), .A3(new_n655_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(G50gat), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT110), .ZN(G1331gat));
  NOR2_X1   g490(.A1(new_n295_), .A2(new_n621_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n609_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n588_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n547_), .A2(G57gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n293_), .A2(new_n609_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n321_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n620_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G57gat), .B1(new_n701_), .B2(new_n547_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n698_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT111), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n698_), .A2(new_n702_), .A3(KEYINPUT111), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1332gat));
  OAI211_X1 g506(.A(new_n544_), .B(new_n700_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(G64gat), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G64gat), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n672_), .A2(G64gat), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n710_), .A2(new_n711_), .B1(new_n695_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT113), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(G1333gat));
  INV_X1    g514(.A(G71gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n696_), .A2(new_n716_), .A3(new_n587_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT49), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n620_), .A2(new_n700_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n587_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n718_), .B1(new_n720_), .B2(G71gat), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT49), .B(new_n716_), .C1(new_n719_), .C2(new_n587_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n717_), .B1(new_n721_), .B2(new_n722_), .ZN(G1334gat));
  OR3_X1    g522(.A1(new_n695_), .A2(G78gat), .A3(new_n491_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n719_), .A2(new_n492_), .ZN(new_n725_));
  XOR2_X1   g524(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(G78gat), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(G78gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(G1335gat));
  AND2_X1   g528(.A1(new_n650_), .A2(new_n321_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n694_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n205_), .A3(new_n445_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n660_), .A2(new_n661_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n621_), .A2(new_n292_), .A3(new_n609_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n445_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n733_), .B1(new_n738_), .B2(new_n205_), .ZN(G1336gat));
  OAI21_X1  g538(.A(new_n206_), .B1(new_n731_), .B2(new_n672_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n740_), .A2(KEYINPUT115), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(KEYINPUT115), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n672_), .A2(new_n206_), .ZN(new_n743_));
  AOI22_X1  g542(.A1(new_n741_), .A2(new_n742_), .B1(new_n736_), .B2(new_n743_), .ZN(G1337gat));
  INV_X1    g543(.A(G99gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n736_), .B2(new_n587_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n731_), .A2(new_n386_), .A3(new_n211_), .ZN(new_n747_));
  OR3_X1    g546(.A1(new_n746_), .A2(KEYINPUT51), .A3(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT51), .B1(new_n746_), .B2(new_n747_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1338gat));
  OR3_X1    g549(.A1(new_n731_), .A2(G106gat), .A3(new_n491_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n734_), .A2(new_n492_), .A3(new_n735_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G106gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G106gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n751_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1339gat));
  INV_X1    g559(.A(new_n595_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT75), .B1(new_n593_), .B2(new_n594_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n589_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n607_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n764_), .A2(KEYINPUT116), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n599_), .A2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n599_), .A2(new_n766_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n589_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n764_), .B2(KEYINPUT116), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n765_), .A2(new_n770_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n312_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n301_), .A2(new_n315_), .A3(new_n311_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT118), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n317_), .A2(new_n776_), .A3(new_n771_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n313_), .A2(new_n609_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n303_), .A2(new_n314_), .A3(new_n305_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n307_), .A2(KEYINPUT55), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n312_), .B1(new_n315_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n783_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n779_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n616_), .B1(new_n778_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n771_), .A2(new_n313_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n787_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n783_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n792_), .B(KEYINPUT58), .C1(new_n793_), .C2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT119), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n786_), .A2(new_n787_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(KEYINPUT58), .A4(new_n792_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n796_), .A2(new_n799_), .A3(new_n802_), .A4(new_n258_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT57), .B(new_n616_), .C1(new_n778_), .C2(new_n788_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n791_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n293_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n699_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT54), .B1(new_n258_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT37), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n248_), .A2(new_n257_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n616_), .B2(new_n809_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n621_), .A2(new_n811_), .A3(new_n812_), .A4(new_n699_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n808_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n806_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n545_), .A2(new_n587_), .A3(new_n445_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(KEYINPUT120), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  INV_X1    g618(.A(new_n814_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n805_), .B2(new_n293_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n821_), .B2(new_n816_), .ZN(new_n822_));
  INV_X1    g621(.A(G113gat), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n818_), .A2(new_n822_), .A3(new_n823_), .A4(new_n609_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n815_), .A2(new_n825_), .A3(new_n817_), .A4(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n826_), .B(new_n827_), .C1(new_n821_), .C2(new_n816_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n693_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n824_), .B1(new_n831_), .B2(new_n823_), .ZN(G1340gat));
  INV_X1    g631(.A(KEYINPUT60), .ZN(new_n833_));
  AOI21_X1  g632(.A(G120gat), .B1(new_n321_), .B2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n833_), .B2(G120gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n818_), .A2(new_n822_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n621_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n837_));
  INV_X1    g636(.A(G120gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(G1341gat));
  INV_X1    g638(.A(G127gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n818_), .A2(new_n292_), .A3(new_n822_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n829_), .A2(new_n830_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n292_), .A2(G127gat), .ZN(new_n843_));
  XOR2_X1   g642(.A(new_n843_), .B(KEYINPUT122), .Z(new_n844_));
  AOI22_X1  g643(.A1(new_n840_), .A2(new_n841_), .B1(new_n842_), .B2(new_n844_), .ZN(G1342gat));
  INV_X1    g644(.A(G134gat), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n818_), .A2(new_n822_), .A3(new_n846_), .A4(new_n254_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n811_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n846_), .ZN(G1343gat));
  NOR2_X1   g648(.A1(new_n587_), .A2(new_n547_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n492_), .A3(new_n672_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT123), .B1(new_n815_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n821_), .A2(new_n854_), .A3(new_n851_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n609_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G141gat), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n400_), .B(new_n609_), .C1(new_n853_), .C2(new_n855_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1344gat));
  OAI21_X1  g658(.A(new_n321_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G148gat), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n401_), .B(new_n321_), .C1(new_n853_), .C2(new_n855_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1345gat));
  OAI21_X1  g662(.A(new_n292_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n865_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n292_), .B(new_n867_), .C1(new_n853_), .C2(new_n855_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1346gat));
  INV_X1    g668(.A(G162gat), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n870_), .B(new_n254_), .C1(new_n853_), .C2(new_n855_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n815_), .A2(KEYINPUT123), .A3(new_n852_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n854_), .B1(new_n821_), .B2(new_n851_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n811_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n871_), .B1(new_n870_), .B2(new_n874_), .ZN(G1347gat));
  NOR2_X1   g674(.A1(new_n821_), .A2(new_n492_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n446_), .A2(new_n544_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(KEYINPUT62), .B(G169gat), .C1(new_n879_), .C2(new_n693_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n821_), .A2(new_n492_), .A3(new_n693_), .A4(new_n877_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n339_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n498_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(new_n883_), .A3(new_n884_), .ZN(G1348gat));
  XNOR2_X1  g684(.A(new_n876_), .B(KEYINPUT124), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n621_), .A2(new_n343_), .A3(new_n877_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n876_), .A2(new_n321_), .A3(new_n878_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n886_), .A2(new_n887_), .B1(new_n343_), .B2(new_n888_), .ZN(G1349gat));
  NAND2_X1  g688(.A1(new_n815_), .A2(new_n491_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n890_), .A2(new_n362_), .A3(new_n293_), .A4(new_n877_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(KEYINPUT124), .ZN(new_n892_));
  OR3_X1    g691(.A1(new_n821_), .A2(KEYINPUT124), .A3(new_n492_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(new_n292_), .A4(new_n878_), .ZN(new_n894_));
  INV_X1    g693(.A(G183gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n891_), .B1(new_n894_), .B2(new_n895_), .ZN(G1350gat));
  OAI21_X1  g695(.A(G190gat), .B1(new_n879_), .B2(new_n811_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n254_), .A2(new_n494_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT125), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n879_), .B2(new_n899_), .ZN(G1351gat));
  NOR3_X1   g699(.A1(new_n587_), .A2(new_n548_), .A3(new_n672_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n815_), .A2(KEYINPUT126), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903_));
  INV_X1    g702(.A(new_n901_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n821_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G197gat), .B1(new_n906_), .B2(new_n609_), .ZN(new_n907_));
  INV_X1    g706(.A(G197gat), .ZN(new_n908_));
  AOI211_X1 g707(.A(new_n908_), .B(new_n693_), .C1(new_n902_), .C2(new_n905_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1352gat));
  AOI21_X1  g709(.A(KEYINPUT126), .B1(new_n815_), .B2(new_n901_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n821_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n321_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G204gat), .ZN(new_n914_));
  INV_X1    g713(.A(G204gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n906_), .A2(new_n915_), .A3(new_n321_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1353gat));
  OAI21_X1  g716(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n292_), .A2(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n906_), .B2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n923_), .ZN(new_n925_));
  AOI211_X1 g724(.A(new_n925_), .B(new_n920_), .C1(new_n902_), .C2(new_n905_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1354gat));
  INV_X1    g726(.A(G218gat), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n906_), .A2(new_n928_), .A3(new_n254_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n811_), .B1(new_n902_), .B2(new_n905_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n928_), .B2(new_n930_), .ZN(G1355gat));
endmodule


