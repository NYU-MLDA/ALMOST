//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT12), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G85gat), .B(G92gat), .Z(new_n211_));
  NOR2_X1   g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n211_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT8), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(KEYINPUT64), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n217_), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT10), .B(G99gat), .Z(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n211_), .A2(KEYINPUT9), .ZN(new_n230_));
  INV_X1    g029(.A(G85gat), .ZN(new_n231_));
  INV_X1    g030(.A(G92gat), .ZN(new_n232_));
  OR3_X1    g031(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT9), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n226_), .A2(new_n229_), .A3(new_n230_), .A4(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT65), .B1(new_n225_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236_));
  INV_X1    g035(.A(new_n234_), .ZN(new_n237_));
  AOI211_X1 g036(.A(new_n236_), .B(new_n237_), .C1(new_n221_), .C2(new_n224_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n210_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G230gat), .A2(G233gat), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n237_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n207_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n241_), .A2(new_n207_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n208_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n239_), .A2(new_n240_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n242_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(G230gat), .A3(G233gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(G120gat), .B(G148gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(G176gat), .B(G204gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n253_), .A2(KEYINPUT66), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n246_), .A2(new_n248_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT13), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT72), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G29gat), .B(G36gat), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n262_), .A2(KEYINPUT69), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(KEYINPUT69), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G43gat), .B(G50gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT70), .B(KEYINPUT15), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G232gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT35), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n270_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n241_), .A2(new_n280_), .B1(new_n277_), .B2(new_n276_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n273_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n273_), .B2(new_n281_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n261_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n273_), .A2(new_n281_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n278_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n273_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(KEYINPUT72), .A3(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G190gat), .B(G218gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT71), .ZN(new_n290_));
  XOR2_X1   g089(.A(G134gat), .B(G162gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT36), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n284_), .A2(new_n288_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT36), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n286_), .A2(new_n295_), .A3(new_n292_), .A4(new_n287_), .ZN(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n296_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n293_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT37), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G15gat), .B(G22gat), .ZN(new_n304_));
  INV_X1    g103(.A(G1gat), .ZN(new_n305_));
  INV_X1    g104(.A(G8gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT14), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G8gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n308_), .B(new_n309_), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n207_), .B(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G231gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT17), .ZN(new_n315_));
  XOR2_X1   g114(.A(G127gat), .B(G155gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT16), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G183gat), .B(G211gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  OR3_X1    g118(.A1(new_n314_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(KEYINPUT17), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n303_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n260_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT74), .ZN(new_n327_));
  INV_X1    g126(.A(new_n310_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n272_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n280_), .A2(new_n310_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G229gat), .A2(G233gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n270_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n334_), .B2(new_n331_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G141gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G169gat), .B(G197gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n337_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT86), .ZN(new_n343_));
  OR2_X1    g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT21), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n344_), .A2(KEYINPUT21), .A3(new_n345_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n349_), .A2(new_n350_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(KEYINPUT1), .B2(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n355_), .A2(KEYINPUT1), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(G141gat), .A2(G148gat), .ZN(new_n359_));
  INV_X1    g158(.A(G141gat), .ZN(new_n360_));
  INV_X1    g159(.A(G148gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n354_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n355_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(KEYINPUT83), .A3(new_n355_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT3), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n371_), .B1(G141gat), .B2(G148gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  AND3_X1   g172(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n373_), .A2(new_n376_), .A3(KEYINPUT82), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT82), .B1(new_n373_), .B2(new_n376_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n369_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT84), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(KEYINPUT84), .B(new_n369_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n363_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n343_), .B(new_n353_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n386_), .B(new_n353_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n387_));
  AND2_X1   g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388_));
  AOI22_X1  g187(.A1(KEYINPUT87), .A2(new_n385_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n385_), .A2(KEYINPUT87), .A3(new_n388_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT89), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n385_), .A2(KEYINPUT87), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n387_), .A2(new_n388_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n385_), .A2(KEYINPUT87), .A3(new_n388_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n392_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n393_), .A3(new_n398_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT88), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n397_), .A2(new_n404_), .A3(new_n393_), .A4(new_n398_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n394_), .A2(new_n401_), .A3(new_n403_), .A4(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G22gat), .B(G50gat), .Z(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n383_), .A2(new_n384_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n408_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n413_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n407_), .A3(new_n411_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT90), .B1(new_n399_), .B2(new_n392_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n402_), .A2(new_n417_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n399_), .A2(KEYINPUT90), .A3(new_n392_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n406_), .A2(new_n418_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT23), .ZN(new_n424_));
  INV_X1    g223(.A(G183gat), .ZN(new_n425_));
  INV_X1    g224(.A(G190gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT25), .B(G183gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT26), .B1(new_n426_), .B2(KEYINPUT76), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n426_), .A2(KEYINPUT26), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n438_), .B(new_n439_), .C1(new_n440_), .C2(KEYINPUT76), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n431_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(KEYINPUT22), .B(G169gat), .Z(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT78), .B1(new_n443_), .B2(G176gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT22), .B(G169gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT78), .ZN(new_n446_));
  INV_X1    g245(.A(G176gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n425_), .A2(new_n426_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n427_), .A2(new_n428_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n434_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n442_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT20), .B1(new_n453_), .B2(new_n353_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G226gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT19), .ZN(new_n456_));
  INV_X1    g255(.A(new_n353_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT92), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n443_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n445_), .A2(KEYINPUT92), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n447_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n451_), .A2(KEYINPUT93), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n451_), .A2(KEYINPUT93), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n434_), .A4(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n436_), .A2(new_n432_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n438_), .B(KEYINPUT91), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT26), .B(G190gat), .Z(new_n467_));
  OAI211_X1 g266(.A(new_n431_), .B(new_n465_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n457_), .B1(new_n464_), .B2(new_n468_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n454_), .A2(new_n456_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n456_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT20), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n453_), .B2(new_n353_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n464_), .A2(new_n468_), .A3(new_n457_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n471_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n456_), .B1(new_n454_), .B2(new_n469_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G8gat), .B(G36gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT18), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G64gat), .B(G92gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT32), .ZN(new_n484_));
  MUX2_X1   g283(.A(new_n476_), .B(new_n479_), .S(new_n484_), .Z(new_n485_));
  INV_X1    g284(.A(new_n363_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n373_), .A2(new_n376_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n373_), .A2(new_n376_), .A3(KEYINPUT82), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT84), .B1(new_n491_), .B2(new_n369_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n382_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n486_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G127gat), .B(G134gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G113gat), .B(G120gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n494_), .A2(KEYINPUT95), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT95), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(new_n383_), .B2(new_n497_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT96), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n383_), .A2(KEYINPUT96), .A3(new_n497_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n502_), .A2(KEYINPUT4), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G225gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT4), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n494_), .A2(new_n508_), .A3(new_n498_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT97), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT97), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n494_), .A2(new_n511_), .A3(new_n508_), .A4(new_n498_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n507_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n506_), .A2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n504_), .A2(new_n505_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(new_n507_), .A3(new_n502_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G29gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(G85gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT0), .B(G57gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  AND3_X1   g319(.A1(new_n514_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n520_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n485_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT98), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n483_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n442_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n452_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n472_), .B1(new_n529_), .B2(new_n457_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n464_), .A2(new_n468_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n353_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n471_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n353_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n534_));
  AND4_X1   g333(.A1(KEYINPUT20), .A2(new_n474_), .A3(new_n471_), .A4(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n526_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n477_), .A2(new_n483_), .A3(new_n478_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT94), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n477_), .A2(new_n478_), .A3(new_n539_), .A4(new_n483_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n507_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n515_), .A2(new_n542_), .A3(new_n502_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n520_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n542_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n506_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n541_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n521_), .A2(KEYINPUT33), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n514_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT33), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n549_), .A3(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(KEYINPUT98), .B(new_n485_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n423_), .A2(new_n525_), .A3(new_n553_), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G227gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT80), .ZN(new_n557_));
  XOR2_X1   g356(.A(G71gat), .B(G99gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n453_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G15gat), .B(G43gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT79), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT30), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n560_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT81), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n497_), .B(KEYINPUT31), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n564_), .A2(KEYINPUT81), .ZN(new_n568_));
  MUX2_X1   g367(.A(new_n567_), .B(new_n566_), .S(new_n568_), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT27), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n541_), .A2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(KEYINPUT27), .B(new_n537_), .C1(new_n476_), .C2(new_n483_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT99), .B1(new_n521_), .B2(new_n522_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n514_), .A2(new_n516_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n544_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n550_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n574_), .B1(new_n575_), .B2(new_n579_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n555_), .B(new_n570_), .C1(new_n423_), .C2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n575_), .A2(new_n579_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n574_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n423_), .A2(new_n582_), .A3(new_n583_), .A4(new_n569_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n342_), .B1(new_n581_), .B2(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n327_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n582_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n305_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT38), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n294_), .A2(new_n296_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n581_), .B2(new_n584_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n260_), .A2(new_n342_), .A3(new_n323_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n582_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n588_), .A2(new_n589_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n590_), .A2(new_n596_), .A3(new_n597_), .ZN(G1324gat));
  NAND3_X1  g397(.A1(new_n586_), .A2(new_n306_), .A3(new_n574_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G8gat), .B1(new_n595_), .B2(new_n583_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT100), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(KEYINPUT100), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n602_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n599_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n606_), .B(new_n608_), .ZN(G1325gat));
  OAI21_X1  g408(.A(G15gat), .B1(new_n595_), .B2(new_n570_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT41), .Z(new_n611_));
  INV_X1    g410(.A(G15gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n586_), .A2(new_n612_), .A3(new_n569_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(G1326gat));
  OAI21_X1  g413(.A(G22gat), .B1(new_n595_), .B2(new_n423_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT42), .ZN(new_n616_));
  INV_X1    g415(.A(G22gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n423_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n586_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(G1327gat));
  NAND2_X1  g419(.A1(new_n592_), .A2(new_n323_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n260_), .A2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n585_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(G29gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n624_), .A3(new_n587_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n260_), .A2(new_n342_), .A3(new_n324_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT43), .ZN(new_n627_));
  AND4_X1   g426(.A1(new_n423_), .A2(new_n525_), .A3(new_n553_), .A4(new_n554_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n570_), .B1(new_n580_), .B2(new_n423_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n584_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n298_), .A2(KEYINPUT102), .A3(new_n302_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT102), .B1(new_n298_), .B2(new_n302_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n627_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n303_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n627_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n581_), .B2(new_n584_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n626_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(KEYINPUT44), .B(new_n626_), .C1(new_n634_), .C2(new_n637_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n587_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(KEYINPUT103), .A3(G29gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT103), .B1(new_n643_), .B2(G29gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n625_), .B1(new_n644_), .B2(new_n645_), .ZN(G1328gat));
  NAND3_X1  g445(.A1(new_n640_), .A2(new_n574_), .A3(new_n641_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(new_n648_), .A3(G36gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n574_), .B(KEYINPUT105), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(G36gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n585_), .A2(new_n622_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT106), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n585_), .A2(new_n622_), .A3(new_n654_), .A4(new_n651_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n653_), .A2(new_n655_), .A3(KEYINPUT45), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT45), .B1(new_n653_), .B2(new_n655_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n649_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n648_), .B1(new_n647_), .B2(G36gat), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT107), .B(KEYINPUT46), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n647_), .A2(G36gat), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT104), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n649_), .A3(new_n658_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT46), .B1(new_n665_), .B2(KEYINPUT107), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n662_), .A2(new_n666_), .ZN(G1329gat));
  AOI21_X1  g466(.A(G43gat), .B1(new_n623_), .B2(new_n569_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT108), .Z(new_n669_));
  NAND3_X1  g468(.A1(new_n642_), .A2(G43gat), .A3(new_n569_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g471(.A(G50gat), .B1(new_n623_), .B2(new_n618_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n618_), .A2(G50gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n642_), .B2(new_n674_), .ZN(G1331gat));
  AOI21_X1  g474(.A(new_n341_), .B1(new_n581_), .B2(new_n584_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n325_), .A2(new_n259_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(G57gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n587_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n259_), .A2(new_n341_), .A3(new_n323_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n593_), .A2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(new_n587_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n684_), .B2(new_n680_), .ZN(G1332gat));
  INV_X1    g484(.A(G64gat), .ZN(new_n686_));
  INV_X1    g485(.A(new_n650_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n683_), .B2(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT48), .Z(new_n689_));
  NAND3_X1  g488(.A1(new_n679_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT109), .ZN(G1333gat));
  INV_X1    g491(.A(G71gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n683_), .B2(new_n569_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT49), .Z(new_n695_));
  NAND2_X1  g494(.A1(new_n569_), .A2(new_n693_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n678_), .B2(new_n696_), .ZN(G1334gat));
  INV_X1    g496(.A(G78gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n683_), .B2(new_n618_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT50), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n679_), .A2(new_n698_), .A3(new_n618_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1335gat));
  NOR2_X1   g501(.A1(new_n259_), .A2(new_n621_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n676_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n231_), .A3(new_n587_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n634_), .A2(new_n637_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n259_), .A2(new_n341_), .A3(new_n324_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT110), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT110), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(new_n587_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n706_), .B1(new_n713_), .B2(new_n231_), .ZN(G1336gat));
  OAI21_X1  g513(.A(new_n232_), .B1(new_n704_), .B2(new_n583_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT111), .Z(new_n716_));
  NAND2_X1  g515(.A1(new_n687_), .A2(G92gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT112), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n712_), .B2(new_n718_), .ZN(G1337gat));
  NAND4_X1  g518(.A1(new_n676_), .A2(new_n703_), .A3(new_n569_), .A4(new_n227_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT113), .Z(new_n721_));
  NAND2_X1  g520(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n569_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(G99gat), .ZN(new_n725_));
  NOR2_X1   g524(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT115), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n725_), .B(new_n728_), .ZN(G1338gat));
  NAND3_X1  g528(.A1(new_n705_), .A2(new_n228_), .A3(new_n618_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n707_), .A2(new_n618_), .A3(new_n708_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n228_), .B1(KEYINPUT116), .B2(KEYINPUT52), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n730_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g536(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n239_), .A2(KEYINPUT55), .A3(new_n245_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n240_), .A2(KEYINPUT117), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n246_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n253_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n740_), .B2(new_n742_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT118), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(KEYINPUT56), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n246_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n341_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n258_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n335_), .A2(new_n340_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n331_), .B1(new_n280_), .B2(new_n310_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n330_), .A2(new_n333_), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n329_), .A2(new_n758_), .B1(new_n759_), .B2(new_n331_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n760_), .B2(new_n340_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n756_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n591_), .B(new_n739_), .C1(new_n755_), .C2(new_n762_), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n751_), .A2(new_n754_), .B1(new_n756_), .B2(new_n761_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n738_), .B1(new_n764_), .B2(new_n592_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT120), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n752_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n748_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT56), .B1(new_n745_), .B2(new_n747_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(KEYINPUT58), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n635_), .B1(new_n771_), .B2(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n763_), .B(new_n765_), .C1(new_n773_), .C2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n326_), .A2(new_n342_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT54), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n326_), .A2(new_n779_), .A3(new_n342_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n776_), .A2(new_n323_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  NOR4_X1   g580(.A1(new_n618_), .A2(new_n582_), .A3(new_n574_), .A4(new_n570_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(G113gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(new_n341_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n781_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT59), .A3(new_n782_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT59), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n342_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n786_), .B1(new_n791_), .B2(new_n785_), .ZN(G1340gat));
  INV_X1    g591(.A(G120gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n259_), .B2(KEYINPUT60), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n784_), .B(new_n794_), .C1(KEYINPUT60), .C2(new_n793_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n259_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n793_), .ZN(G1341gat));
  INV_X1    g596(.A(KEYINPUT121), .ZN(new_n798_));
  INV_X1    g597(.A(G127gat), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n788_), .A2(new_n790_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n324_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n784_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n324_), .A2(new_n799_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n798_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n323_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n806_));
  OAI221_X1 g605(.A(KEYINPUT121), .B1(new_n802_), .B2(new_n803_), .C1(new_n806_), .C2(new_n799_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1342gat));
  INV_X1    g607(.A(G134gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n784_), .A2(new_n809_), .A3(new_n592_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n303_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n809_), .ZN(G1343gat));
  NAND4_X1  g611(.A1(new_n650_), .A2(new_n618_), .A3(new_n587_), .A4(new_n570_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT122), .Z(new_n814_));
  NAND2_X1  g613(.A1(new_n787_), .A2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n342_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(new_n360_), .ZN(G1344gat));
  NOR2_X1   g616(.A1(new_n815_), .A2(new_n259_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(new_n361_), .ZN(G1345gat));
  NOR2_X1   g618(.A1(new_n815_), .A2(new_n323_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT61), .B(G155gat), .Z(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1346gat));
  INV_X1    g621(.A(G162gat), .ZN(new_n823_));
  NOR4_X1   g622(.A1(new_n815_), .A2(new_n823_), .A3(new_n632_), .A4(new_n631_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n815_), .B2(new_n591_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n825_), .A2(KEYINPUT123), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(KEYINPUT123), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n824_), .B1(new_n826_), .B2(new_n827_), .ZN(G1347gat));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n829_));
  NOR4_X1   g628(.A1(new_n650_), .A2(new_n618_), .A3(new_n587_), .A4(new_n570_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n787_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n342_), .ZN(new_n832_));
  INV_X1    g631(.A(G169gat), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT124), .B(new_n829_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n833_), .B1(new_n836_), .B2(KEYINPUT62), .ZN(new_n837_));
  OAI221_X1 g636(.A(new_n837_), .B1(new_n836_), .B2(KEYINPUT62), .C1(new_n831_), .C2(new_n342_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n834_), .A2(new_n835_), .A3(new_n838_), .ZN(G1348gat));
  INV_X1    g638(.A(new_n831_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n260_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n447_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT125), .B(G176gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n841_), .B2(new_n844_), .ZN(G1349gat));
  NOR2_X1   g644(.A1(new_n831_), .A2(new_n323_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(G183gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n466_), .B2(new_n846_), .ZN(G1350gat));
  OAI21_X1  g647(.A(G190gat), .B1(new_n831_), .B2(new_n303_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n591_), .A2(new_n467_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n831_), .B2(new_n850_), .ZN(G1351gat));
  NOR4_X1   g650(.A1(new_n650_), .A2(new_n587_), .A3(new_n423_), .A4(new_n569_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n787_), .A2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n342_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT126), .B(G197gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1352gat));
  INV_X1    g655(.A(new_n853_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT127), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n259_), .B1(new_n858_), .B2(G204gat), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(G204gat), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n860_), .B(new_n861_), .Z(G1353gat));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n324_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n864_));
  AND2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n863_), .B2(new_n864_), .ZN(G1354gat));
  OR3_X1    g666(.A1(new_n853_), .A2(G218gat), .A3(new_n591_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G218gat), .B1(new_n853_), .B2(new_n303_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1355gat));
endmodule


