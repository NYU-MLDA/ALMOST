//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT73), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT73), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(new_n204_), .A3(new_n206_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT15), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT76), .ZN(new_n213_));
  INV_X1    g012(.A(G15gat), .ZN(new_n214_));
  INV_X1    g013(.A(G22gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G15gat), .A2(G22gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G1gat), .A2(G8gat), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n216_), .A2(new_n217_), .B1(KEYINPUT14), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n213_), .B(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n211_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n210_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT78), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n220_), .B(new_n210_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(G229gat), .A3(G233gat), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G113gat), .B(G141gat), .Z(new_n230_));
  XNOR2_X1  g029(.A(G169gat), .B(G197gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n229_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G64gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G57gat), .ZN(new_n236_));
  INV_X1    g035(.A(G57gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G64gat), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n236_), .A2(new_n238_), .A3(KEYINPUT11), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT68), .B(G71gat), .ZN(new_n241_));
  INV_X1    g040(.A(G78gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n241_), .A2(new_n242_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n240_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT68), .B(G71gat), .Z(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G78gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT11), .B1(new_n236_), .B2(new_n238_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n248_), .B(new_n243_), .C1(new_n249_), .C2(new_n239_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n252_), .A2(KEYINPUT9), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(KEYINPUT9), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n253_), .A2(G85gat), .A3(G92gat), .A4(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G85gat), .ZN(new_n256_));
  INV_X1    g055(.A(G92gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G85gat), .A2(G92gat), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n258_), .A2(new_n252_), .A3(KEYINPUT9), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT66), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(G99gat), .ZN(new_n264_));
  INV_X1    g063(.A(G106gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT6), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(G99gat), .A3(G106gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n255_), .A2(KEYINPUT66), .A3(new_n260_), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT10), .B(G99gat), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n265_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n263_), .A2(new_n269_), .A3(new_n270_), .A4(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT8), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G99gat), .A2(G106gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT7), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n266_), .A2(new_n268_), .A3(KEYINPUT67), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n276_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n258_), .A2(new_n259_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n274_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n274_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(new_n269_), .B2(new_n278_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n251_), .B(new_n273_), .C1(new_n282_), .C2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G230gat), .A2(G233gat), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT64), .Z(new_n289_));
  OAI21_X1  g088(.A(new_n273_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n251_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n287_), .B(new_n289_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n291_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n285_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n289_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G120gat), .B(G148gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT5), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G176gat), .B(G204gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n295_), .A2(new_n299_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n304_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT13), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT13), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(KEYINPUT71), .A3(new_n314_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n234_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(G127gat), .B(G155gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT16), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G183gat), .B(G211gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT17), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G231gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n220_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(new_n251_), .ZN(new_n329_));
  AOI211_X1 g128(.A(new_n326_), .B(new_n329_), .C1(new_n325_), .C2(new_n323_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n326_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n319_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G85gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT0), .B(G57gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT86), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT85), .B(KEYINPUT3), .ZN(new_n343_));
  OR2_X1    g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT3), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n347_), .A2(KEYINPUT85), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(KEYINPUT85), .ZN(new_n349_));
  OAI211_X1 g148(.A(KEYINPUT86), .B(new_n346_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT2), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(G141gat), .A3(G148gat), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n352_), .A2(new_n354_), .B1(new_n344_), .B2(KEYINPUT3), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n345_), .A2(new_n350_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n344_), .A2(new_n351_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n359_), .B1(KEYINPUT1), .B2(new_n357_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n357_), .A2(KEYINPUT1), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n365_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT87), .ZN(new_n371_));
  XOR2_X1   g170(.A(G127gat), .B(G134gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(G113gat), .B(G120gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n369_), .A2(new_n371_), .A3(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n341_), .B1(new_n375_), .B2(KEYINPUT4), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n367_), .A2(new_n374_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(KEYINPUT4), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT92), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n375_), .A2(new_n378_), .A3(KEYINPUT92), .A4(KEYINPUT4), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n376_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n375_), .A2(new_n378_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(new_n341_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n339_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n381_), .A2(new_n382_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n376_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n338_), .B1(new_n384_), .B2(new_n341_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT95), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT95), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n383_), .A2(new_n393_), .A3(new_n390_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n386_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT96), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n389_), .A2(KEYINPUT95), .A3(new_n391_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n393_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT96), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n386_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT27), .ZN(new_n403_));
  OR2_X1    g202(.A1(G197gat), .A2(G204gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G197gat), .A2(G204gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT21), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(KEYINPUT21), .A3(new_n405_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n409_), .A2(new_n410_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G169gat), .ZN(new_n416_));
  INV_X1    g215(.A(G183gat), .ZN(new_n417_));
  INV_X1    g216(.A(G190gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT23), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT23), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(G183gat), .A3(G190gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(KEYINPUT82), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT82), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n423_), .B(KEYINPUT23), .C1(new_n417_), .C2(new_n418_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT79), .B(G190gat), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n426_), .A2(new_n417_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n416_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT26), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n418_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT25), .B(G183gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT24), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(G169gat), .B2(G176gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436_));
  INV_X1    g235(.A(G169gat), .ZN(new_n437_));
  INV_X1    g236(.A(G176gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n433_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n440_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n434_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n419_), .A2(new_n421_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n446_), .B(new_n447_), .C1(new_n442_), .C2(new_n441_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n414_), .B(new_n428_), .C1(new_n444_), .C2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n416_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n419_), .A2(new_n421_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT26), .B(G190gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n432_), .A2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n446_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n425_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT90), .A4(new_n441_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n446_), .A2(new_n441_), .A3(new_n454_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n458_), .B1(new_n459_), .B2(new_n425_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n452_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n461_));
  OAI211_X1 g260(.A(KEYINPUT20), .B(new_n449_), .C1(new_n461_), .C2(new_n414_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT19), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n428_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n467_));
  AOI211_X1 g266(.A(new_n466_), .B(new_n464_), .C1(new_n467_), .C2(new_n413_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n461_), .A2(new_n414_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(G8gat), .B(G36gat), .Z(new_n472_));
  XNOR2_X1  g271(.A(G64gat), .B(G92gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n462_), .A2(new_n464_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n476_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n403_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n413_), .A2(new_n452_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n455_), .A2(new_n456_), .A3(new_n441_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n466_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n467_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(new_n414_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n486_), .A2(new_n464_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n462_), .A2(new_n464_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n476_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n478_), .A2(new_n479_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT27), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n481_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G15gat), .B(G43gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G71gat), .B(G99gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n467_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n467_), .A2(new_n496_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G227gat), .A2(G233gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n500_), .B(KEYINPUT83), .Z(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT30), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n497_), .A2(new_n502_), .A3(new_n498_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n374_), .B(KEYINPUT31), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n506_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n510_));
  MUX2_X1   g309(.A(new_n509_), .B(new_n508_), .S(new_n510_), .Z(new_n511_));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n413_), .B1(new_n370_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G228gat), .ZN(new_n515_));
  INV_X1    g314(.A(G233gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT87), .B1(new_n361_), .B2(new_n366_), .ZN(new_n519_));
  AOI211_X1 g318(.A(new_n368_), .B(new_n365_), .C1(new_n356_), .C2(new_n360_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n513_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n414_), .A2(new_n517_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n518_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G78gat), .B(G106gat), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n512_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n513_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G22gat), .B(G50gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT28), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n527_), .B(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT89), .B1(new_n526_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n531_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n369_), .A2(KEYINPUT29), .A3(new_n371_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n534_), .A2(new_n522_), .B1(new_n517_), .B2(new_n514_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n525_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT88), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n524_), .B(new_n536_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n526_), .A2(KEYINPUT89), .A3(new_n531_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n538_), .B1(new_n533_), .B2(new_n537_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n493_), .A2(new_n511_), .A3(new_n541_), .A4(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n402_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n541_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT33), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n477_), .A2(new_n480_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n375_), .A2(KEYINPUT4), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(new_n341_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n519_), .A2(new_n520_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n377_), .B1(new_n555_), .B2(new_n374_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT92), .B1(new_n556_), .B2(KEYINPUT4), .ZN(new_n557_));
  INV_X1    g356(.A(new_n382_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n554_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n338_), .B1(new_n556_), .B2(new_n341_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n551_), .A2(new_n552_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n390_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n564_), .B2(KEYINPUT33), .ZN(new_n565_));
  NOR4_X1   g364(.A1(new_n383_), .A2(KEYINPUT93), .A3(new_n550_), .A4(new_n390_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n562_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n479_), .A2(KEYINPUT32), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT94), .B1(new_n471_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n478_), .A2(new_n571_), .A3(new_n568_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n569_), .B1(new_n488_), .B2(new_n487_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n399_), .B2(new_n386_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n549_), .B1(new_n567_), .B2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n492_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n396_), .A2(new_n578_), .A3(new_n401_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n511_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n547_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT36), .Z(new_n586_));
  NAND2_X1  g385(.A1(new_n211_), .A2(new_n290_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT74), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n210_), .B(new_n273_), .C1(new_n282_), .C2(new_n284_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n595_), .A2(KEYINPUT75), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(KEYINPUT75), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n596_), .A2(new_n597_), .B1(new_n592_), .B2(new_n591_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n588_), .A2(new_n594_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n594_), .B1(new_n588_), .B2(new_n598_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n586_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n601_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n585_), .A2(KEYINPUT36), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n599_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n582_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n334_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n402_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G1gat), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT97), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n396_), .A2(new_n578_), .A3(new_n401_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n575_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n395_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n564_), .A2(KEYINPUT33), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT93), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n471_), .A2(new_n476_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n490_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n564_), .A2(new_n563_), .A3(KEYINPUT33), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n617_), .A2(new_n620_), .A3(new_n621_), .A4(new_n551_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n548_), .B1(new_n615_), .B2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n581_), .B1(new_n613_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n547_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT37), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n627_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n602_), .A2(new_n605_), .A3(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n333_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n626_), .A2(new_n633_), .A3(new_n319_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n634_), .A2(G1gat), .A3(new_n610_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT38), .Z(new_n636_));
  NAND2_X1  g435(.A1(new_n612_), .A2(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n334_), .A2(new_n492_), .A3(new_n608_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(G8gat), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n638_), .A3(G8gat), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n634_), .A2(G8gat), .A3(new_n493_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1325gat));
  OAI21_X1  g448(.A(G15gat), .B1(new_n609_), .B2(new_n581_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n511_), .A2(new_n214_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n652_), .B(new_n653_), .C1(new_n634_), .C2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT101), .ZN(G1326gat));
  OAI21_X1  g455(.A(G22gat), .B1(new_n609_), .B2(new_n549_), .ZN(new_n657_));
  XOR2_X1   g456(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n548_), .A2(new_n215_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT103), .Z(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n634_), .B2(new_n661_), .ZN(G1327gat));
  OAI21_X1  g461(.A(KEYINPUT43), .B1(new_n582_), .B2(new_n631_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n629_), .A2(new_n630_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n511_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n664_), .B(new_n665_), .C1(new_n666_), .C2(new_n547_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n317_), .A2(new_n318_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n332_), .A3(new_n233_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT44), .B1(new_n668_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n673_), .B(new_n670_), .C1(new_n663_), .C2(new_n667_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n402_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n676_), .A2(KEYINPUT104), .A3(G29gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT104), .B1(new_n676_), .B2(G29gat), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n333_), .A2(new_n606_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n626_), .A2(new_n319_), .A3(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n610_), .A2(G29gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT105), .ZN(new_n682_));
  OAI22_X1  g481(.A1(new_n677_), .A2(new_n678_), .B1(new_n680_), .B2(new_n682_), .ZN(G1328gat));
  INV_X1    g482(.A(new_n680_), .ZN(new_n684_));
  INV_X1    g483(.A(G36gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n492_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT45), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n672_), .A2(new_n674_), .A3(new_n493_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(new_n685_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1329gat));
  INV_X1    g490(.A(G43gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n692_), .B1(new_n680_), .B2(new_n581_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT107), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n511_), .A2(G43gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT106), .B1(new_n675_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698_));
  NOR4_X1   g497(.A1(new_n672_), .A2(new_n674_), .A3(new_n698_), .A4(new_n695_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT47), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n702_), .B(new_n694_), .C1(new_n697_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1330gat));
  INV_X1    g503(.A(G50gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n684_), .A2(new_n705_), .A3(new_n548_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n675_), .A2(new_n548_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(G50gat), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT108), .B(new_n705_), .C1(new_n675_), .C2(new_n548_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(G1331gat));
  NOR2_X1   g510(.A1(new_n632_), .A2(new_n669_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT109), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n582_), .A2(new_n233_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n237_), .B1(new_n715_), .B2(new_n610_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n669_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n332_), .A2(new_n233_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n608_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G57gat), .B1(new_n610_), .B2(KEYINPUT110), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n720_), .B(new_n721_), .C1(KEYINPUT110), .C2(G57gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n716_), .A2(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT111), .Z(G1332gat));
  OAI21_X1  g523(.A(G64gat), .B1(new_n719_), .B2(new_n493_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT48), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n492_), .A2(new_n235_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n715_), .B2(new_n727_), .ZN(G1333gat));
  OAI21_X1  g527(.A(G71gat), .B1(new_n719_), .B2(new_n581_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT49), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n581_), .A2(G71gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n715_), .B2(new_n731_), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n720_), .A2(new_n548_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(G78gat), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n733_), .B2(G78gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n548_), .A2(new_n242_), .ZN(new_n738_));
  OAI22_X1  g537(.A1(new_n736_), .A2(new_n737_), .B1(new_n715_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT112), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT112), .ZN(new_n741_));
  OAI221_X1 g540(.A(new_n741_), .B1(new_n715_), .B2(new_n738_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1335gat));
  NOR3_X1   g542(.A1(new_n669_), .A2(new_n606_), .A3(new_n333_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n714_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n256_), .B1(new_n745_), .B2(new_n610_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT113), .Z(new_n747_));
  NOR3_X1   g546(.A1(new_n669_), .A2(new_n333_), .A3(new_n233_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n665_), .B1(new_n626_), .B2(new_n664_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n667_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT114), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n668_), .A2(new_n753_), .A3(new_n748_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n610_), .A2(new_n256_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n747_), .B1(new_n755_), .B2(new_n756_), .ZN(G1336gat));
  AOI21_X1  g556(.A(new_n493_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n492_), .A2(new_n257_), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n758_), .A2(new_n257_), .B1(new_n745_), .B2(new_n759_), .ZN(G1337gat));
  OR2_X1    g559(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n761_));
  NAND2_X1  g560(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n264_), .B1(new_n755_), .B2(new_n511_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n511_), .A2(new_n271_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n745_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n761_), .B(new_n762_), .C1(new_n763_), .C2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n754_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n753_), .B1(new_n668_), .B2(new_n748_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n511_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G99gat), .ZN(new_n770_));
  INV_X1    g569(.A(new_n765_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n770_), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n766_), .A2(new_n772_), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n668_), .A2(new_n548_), .A3(new_n748_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G106gat), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n549_), .A2(G106gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n714_), .A2(new_n744_), .A3(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT116), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n777_), .A2(new_n778_), .A3(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g582(.A(new_n225_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n222_), .A2(new_n223_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n232_), .B1(new_n227_), .B2(new_n225_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n229_), .A2(new_n232_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n311_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n233_), .A2(new_n305_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n295_), .A2(KEYINPUT118), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT55), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n295_), .A2(KEYINPUT118), .A3(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n287_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n298_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n790_), .A2(KEYINPUT55), .B1(new_n794_), .B2(new_n298_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT119), .B1(new_n799_), .B2(new_n793_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n303_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n796_), .A2(new_n797_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n799_), .A2(KEYINPUT119), .A3(new_n793_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n303_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n789_), .B1(new_n803_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n788_), .B1(new_n808_), .B2(KEYINPUT120), .ZN(new_n809_));
  INV_X1    g608(.A(new_n789_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n806_), .B2(new_n303_), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n802_), .B(new_n304_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT120), .B(new_n810_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n606_), .B1(new_n809_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n813_), .A3(new_n788_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n607_), .A2(new_n816_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n787_), .A2(new_n305_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n631_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n821_), .A2(new_n822_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n333_), .B1(new_n817_), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n315_), .A2(KEYINPUT117), .A3(new_n718_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n631_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT117), .B1(new_n315_), .B2(new_n718_), .ZN(new_n832_));
  OR3_X1    g631(.A1(new_n831_), .A2(KEYINPUT54), .A3(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT54), .B1(new_n831_), .B2(new_n832_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n829_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n549_), .A2(new_n511_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n402_), .A3(new_n493_), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(KEYINPUT121), .Z(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n837_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(G113gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n233_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n837_), .B2(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n821_), .A2(new_n822_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n826_), .A2(new_n827_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT57), .B1(new_n821_), .B2(new_n606_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n332_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n835_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(KEYINPUT59), .A3(new_n841_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n234_), .B1(new_n847_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n845_), .B1(new_n855_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n669_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n843_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n857_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n669_), .B1(new_n847_), .B2(new_n854_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n857_), .ZN(G1341gat));
  INV_X1    g660(.A(G127gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n843_), .A2(new_n862_), .A3(new_n333_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n332_), .B1(new_n847_), .B2(new_n854_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1342gat));
  OAI211_X1 g664(.A(new_n607_), .B(new_n841_), .C1(new_n829_), .C2(new_n836_), .ZN(new_n866_));
  INV_X1    g665(.A(G134gat), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n866_), .A2(KEYINPUT122), .A3(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n847_), .A2(new_n854_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n631_), .A2(new_n867_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n870_), .A2(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1343gat));
  NAND3_X1  g673(.A1(new_n402_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n852_), .B2(new_n835_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n233_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n717_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n333_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  INV_X1    g682(.A(G162gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n876_), .A2(new_n884_), .A3(new_n607_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n837_), .A2(new_n631_), .A3(new_n875_), .ZN(new_n886_));
  OAI211_X1 g685(.A(KEYINPUT123), .B(new_n885_), .C1(new_n886_), .C2(new_n884_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n884_), .B1(new_n876_), .B2(new_n664_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n607_), .A2(new_n884_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n837_), .A2(new_n875_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n888_), .B1(new_n889_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n887_), .A2(new_n892_), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n402_), .A2(new_n493_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n839_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n853_), .A2(new_n233_), .A3(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n897_), .A2(new_n898_), .A3(G169gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n897_), .B2(G169gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n853_), .A2(new_n896_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT22), .B(G169gat), .Z(new_n902_));
  NOR2_X1   g701(.A1(new_n234_), .A2(new_n902_), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT124), .Z(new_n904_));
  OAI22_X1  g703(.A1(new_n899_), .A2(new_n900_), .B1(new_n901_), .B2(new_n904_), .ZN(G1348gat));
  NOR2_X1   g704(.A1(new_n837_), .A2(new_n895_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n438_), .A2(KEYINPUT125), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n438_), .A2(KEYINPUT125), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n906_), .A2(new_n717_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n901_), .A2(new_n669_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n908_), .ZN(G1349gat));
  OAI211_X1 g710(.A(new_n333_), .B(new_n896_), .C1(new_n829_), .C2(new_n836_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n417_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n432_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n853_), .A2(new_n914_), .A3(new_n333_), .A4(new_n896_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n913_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n913_), .B2(new_n915_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1350gat));
  NAND3_X1  g718(.A1(new_n906_), .A2(new_n453_), .A3(new_n607_), .ZN(new_n920_));
  OAI21_X1  g719(.A(G190gat), .B1(new_n901_), .B2(new_n631_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1351gat));
  NAND3_X1  g721(.A1(new_n894_), .A2(new_n548_), .A3(new_n581_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n837_), .A2(new_n923_), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n924_), .A2(G197gat), .A3(new_n233_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G197gat), .B1(new_n924_), .B2(new_n233_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1352gat));
  INV_X1    g726(.A(new_n924_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G204gat), .B1(new_n928_), .B2(new_n669_), .ZN(new_n929_));
  INV_X1    g728(.A(G204gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n924_), .A2(new_n930_), .A3(new_n717_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1353gat));
  AOI21_X1  g731(.A(new_n332_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n934_));
  OR3_X1    g733(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n924_), .A2(new_n933_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n924_), .A2(new_n933_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(new_n935_), .ZN(G1354gat));
  OAI21_X1  g737(.A(G218gat), .B1(new_n928_), .B2(new_n631_), .ZN(new_n939_));
  INV_X1    g738(.A(G218gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n924_), .A2(new_n940_), .A3(new_n607_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1355gat));
endmodule


