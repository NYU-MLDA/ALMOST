// Benchmark "../Benchmarks/c6288" written by ABC on Fri Feb  4 08:49:25 2022

module c6288  ( 
    G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat,
    G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat  );
  input  G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat;
  output G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat;
  wire new_G546gat_, new_G549gat_, new_G552gat_, new_G555gat_, new_G558gat_,
    new_G561gat_, new_G564gat_, new_G567gat_, new_G570gat_, new_G573gat_,
    new_G576gat_, new_G579gat_, new_G582gat_, new_G585gat_, new_G588gat_,
    new_G591gat_, new_G594gat_, new_G597gat_, new_G600gat_, new_G603gat_,
    new_G606gat_, new_G609gat_, new_G612gat_, new_G615gat_, new_G618gat_,
    new_G621gat_, new_G624gat_, new_G627gat_, new_G630gat_, new_G633gat_,
    new_G636gat_, new_G639gat_, new_G642gat_, new_G645gat_, new_G648gat_,
    new_G651gat_, new_G654gat_, new_G657gat_, new_G660gat_, new_G663gat_,
    new_G666gat_, new_G669gat_, new_G672gat_, new_G675gat_, new_G678gat_,
    new_G681gat_, new_G684gat_, new_G687gat_, new_G690gat_, new_G693gat_,
    new_G696gat_, new_G699gat_, new_G702gat_, new_G705gat_, new_G708gat_,
    new_G711gat_, new_G714gat_, new_G717gat_, new_G720gat_, new_G723gat_,
    new_G726gat_, new_G729gat_, new_G732gat_, new_G735gat_, new_G738gat_,
    new_G741gat_, new_G744gat_, new_G747gat_, new_G750gat_, new_G753gat_,
    new_G756gat_, new_G759gat_, new_G762gat_, new_G765gat_, new_G768gat_,
    new_G771gat_, new_G774gat_, new_G777gat_, new_G780gat_, new_G783gat_,
    new_G786gat_, new_G789gat_, new_G792gat_, new_G795gat_, new_G798gat_,
    new_G801gat_, new_G804gat_, new_G807gat_, new_G810gat_, new_G813gat_,
    new_G816gat_, new_G819gat_, new_G822gat_, new_G825gat_, new_G828gat_,
    new_G831gat_, new_G834gat_, new_G837gat_, new_G840gat_, new_G843gat_,
    new_G846gat_, new_G849gat_, new_G852gat_, new_G855gat_, new_G858gat_,
    new_G861gat_, new_G864gat_, new_G867gat_, new_G870gat_, new_G873gat_,
    new_G876gat_, new_G879gat_, new_G882gat_, new_G885gat_, new_G888gat_,
    new_G891gat_, new_G894gat_, new_G897gat_, new_G900gat_, new_G903gat_,
    new_G906gat_, new_G909gat_, new_G912gat_, new_G915gat_, new_G918gat_,
    new_G921gat_, new_G924gat_, new_G927gat_, new_G930gat_, new_G933gat_,
    new_G936gat_, new_G939gat_, new_G942gat_, new_G945gat_, new_G948gat_,
    new_G951gat_, new_G954gat_, new_G957gat_, new_G960gat_, new_G963gat_,
    new_G966gat_, new_G969gat_, new_G972gat_, new_G975gat_, new_G978gat_,
    new_G981gat_, new_G984gat_, new_G987gat_, new_G990gat_, new_G993gat_,
    new_G996gat_, new_G999gat_, new_G1002gat_, new_G1005gat_,
    new_G1008gat_, new_G1011gat_, new_G1014gat_, new_G1017gat_,
    new_G1020gat_, new_G1023gat_, new_G1026gat_, new_G1029gat_,
    new_G1032gat_, new_G1035gat_, new_G1038gat_, new_G1041gat_,
    new_G1044gat_, new_G1047gat_, new_G1050gat_, new_G1053gat_,
    new_G1056gat_, new_G1059gat_, new_G1062gat_, new_G1065gat_,
    new_G1068gat_, new_G1071gat_, new_G1074gat_, new_G1077gat_,
    new_G1080gat_, new_G1083gat_, new_G1086gat_, new_G1089gat_,
    new_G1092gat_, new_G1095gat_, new_G1098gat_, new_G1101gat_,
    new_G1104gat_, new_G1107gat_, new_G1110gat_, new_G1113gat_,
    new_G1116gat_, new_G1119gat_, new_G1122gat_, new_G1125gat_,
    new_G1128gat_, new_G1131gat_, new_G1134gat_, new_G1137gat_,
    new_G1140gat_, new_G1143gat_, new_G1146gat_, new_G1149gat_,
    new_G1152gat_, new_G1155gat_, new_G1158gat_, new_G1161gat_,
    new_G1164gat_, new_G1167gat_, new_G1170gat_, new_G1173gat_,
    new_G1176gat_, new_G1179gat_, new_G1182gat_, new_G1185gat_,
    new_G1188gat_, new_G1191gat_, new_G1194gat_, new_G1197gat_,
    new_G1200gat_, new_G1203gat_, new_G1206gat_, new_G1209gat_,
    new_G1212gat_, new_G1215gat_, new_G1218gat_, new_G1221gat_,
    new_G1224gat_, new_G1227gat_, new_G1230gat_, new_G1233gat_,
    new_G1236gat_, new_G1239gat_, new_G1242gat_, new_G1245gat_,
    new_G1248gat_, new_G1251gat_, new_G1254gat_, new_G1257gat_,
    new_G1260gat_, new_G1263gat_, new_G1266gat_, new_G1269gat_,
    new_G1272gat_, new_G1275gat_, new_G1278gat_, new_G1281gat_,
    new_G1284gat_, new_G1287gat_, new_G1290gat_, new_G1293gat_,
    new_G1296gat_, new_G1299gat_, new_G1302gat_, new_G1305gat_,
    new_G1308gat_, new_G1311gat_, new_G1315gat_, new_G1319gat_,
    new_G1323gat_, new_G1327gat_, new_G1331gat_, new_G1335gat_,
    new_G1339gat_, new_G1343gat_, new_G1347gat_, new_G1351gat_,
    new_G1355gat_, new_G1359gat_, new_G1363gat_, new_G1367gat_,
    new_G1371gat_, new_G1372gat_, new_G1373gat_, new_G1374gat_,
    new_G1375gat_, new_G1376gat_, new_G1377gat_, new_G1378gat_,
    new_G1379gat_, new_G1380gat_, new_G1381gat_, new_G1382gat_,
    new_G1383gat_, new_G1384gat_, new_G1385gat_, new_G1386gat_,
    new_G1387gat_, new_G1388gat_, new_G1389gat_, new_G1390gat_,
    new_G1391gat_, new_G1392gat_, new_G1393gat_, new_G1394gat_,
    new_G1395gat_, new_G1396gat_, new_G1397gat_, new_G1398gat_,
    new_G1399gat_, new_G1400gat_, new_G1401gat_, new_G1404gat_,
    new_G1407gat_, new_G1410gat_, new_G1413gat_, new_G1416gat_,
    new_G1419gat_, new_G1422gat_, new_G1425gat_, new_G1428gat_,
    new_G1431gat_, new_G1434gat_, new_G1437gat_, new_G1440gat_,
    new_G1443gat_, new_G1446gat_, new_G1450gat_, new_G1454gat_,
    new_G1458gat_, new_G1462gat_, new_G1466gat_, new_G1470gat_,
    new_G1474gat_, new_G1478gat_, new_G1482gat_, new_G1486gat_,
    new_G1490gat_, new_G1494gat_, new_G1498gat_, new_G1502gat_,
    new_G1506gat_, new_G1507gat_, new_G1508gat_, new_G1511gat_,
    new_G1512gat_, new_G1513gat_, new_G1516gat_, new_G1517gat_,
    new_G1518gat_, new_G1521gat_, new_G1522gat_, new_G1523gat_,
    new_G1526gat_, new_G1527gat_, new_G1528gat_, new_G1531gat_,
    new_G1532gat_, new_G1533gat_, new_G1536gat_, new_G1537gat_,
    new_G1538gat_, new_G1541gat_, new_G1542gat_, new_G1543gat_,
    new_G1546gat_, new_G1547gat_, new_G1548gat_, new_G1551gat_,
    new_G1552gat_, new_G1553gat_, new_G1556gat_, new_G1557gat_,
    new_G1558gat_, new_G1561gat_, new_G1562gat_, new_G1563gat_,
    new_G1566gat_, new_G1567gat_, new_G1568gat_, new_G1571gat_,
    new_G1572gat_, new_G1573gat_, new_G1576gat_, new_G1577gat_,
    new_G1578gat_, new_G1582gat_, new_G1585gat_, new_G1588gat_,
    new_G1591gat_, new_G1594gat_, new_G1597gat_, new_G1600gat_,
    new_G1603gat_, new_G1606gat_, new_G1609gat_, new_G1612gat_,
    new_G1615gat_, new_G1618gat_, new_G1621gat_, new_G1624gat_,
    new_G1628gat_, new_G1632gat_, new_G1636gat_, new_G1640gat_,
    new_G1644gat_, new_G1648gat_, new_G1652gat_, new_G1656gat_,
    new_G1660gat_, new_G1664gat_, new_G1668gat_, new_G1672gat_,
    new_G1676gat_, new_G1680gat_, new_G1684gat_, new_G1685gat_,
    new_G1686gat_, new_G1687gat_, new_G1688gat_, new_G1689gat_,
    new_G1690gat_, new_G1691gat_, new_G1692gat_, new_G1693gat_,
    new_G1694gat_, new_G1695gat_, new_G1696gat_, new_G1697gat_,
    new_G1698gat_, new_G1699gat_, new_G1700gat_, new_G1701gat_,
    new_G1702gat_, new_G1703gat_, new_G1704gat_, new_G1705gat_,
    new_G1706gat_, new_G1707gat_, new_G1708gat_, new_G1709gat_,
    new_G1710gat_, new_G1711gat_, new_G1712gat_, new_G1713gat_,
    new_G1714gat_, new_G1717gat_, new_G1720gat_, new_G1723gat_,
    new_G1726gat_, new_G1729gat_, new_G1732gat_, new_G1735gat_,
    new_G1738gat_, new_G1741gat_, new_G1744gat_, new_G1747gat_,
    new_G1750gat_, new_G1753gat_, new_G1756gat_, new_G1759gat_,
    new_G1763gat_, new_G1767gat_, new_G1771gat_, new_G1775gat_,
    new_G1779gat_, new_G1783gat_, new_G1787gat_, new_G1791gat_,
    new_G1795gat_, new_G1799gat_, new_G1803gat_, new_G1807gat_,
    new_G1811gat_, new_G1815gat_, new_G1819gat_, new_G1820gat_,
    new_G1821gat_, new_G1824gat_, new_G1825gat_, new_G1826gat_,
    new_G1829gat_, new_G1830gat_, new_G1831gat_, new_G1834gat_,
    new_G1835gat_, new_G1836gat_, new_G1839gat_, new_G1840gat_,
    new_G1841gat_, new_G1844gat_, new_G1845gat_, new_G1846gat_,
    new_G1849gat_, new_G1850gat_, new_G1851gat_, new_G1854gat_,
    new_G1855gat_, new_G1856gat_, new_G1859gat_, new_G1860gat_,
    new_G1861gat_, new_G1864gat_, new_G1865gat_, new_G1866gat_,
    new_G1869gat_, new_G1870gat_, new_G1871gat_, new_G1874gat_,
    new_G1875gat_, new_G1876gat_, new_G1879gat_, new_G1880gat_,
    new_G1881gat_, new_G1884gat_, new_G1885gat_, new_G1886gat_,
    new_G1889gat_, new_G1890gat_, new_G1891gat_, new_G1894gat_,
    new_G1897gat_, new_G1902gat_, new_G1905gat_, new_G1908gat_,
    new_G1911gat_, new_G1914gat_, new_G1917gat_, new_G1920gat_,
    new_G1923gat_, new_G1926gat_, new_G1929gat_, new_G1932gat_,
    new_G1935gat_, new_G1938gat_, new_G1941gat_, new_G1945gat_,
    new_G1946gat_, new_G1947gat_, new_G1951gat_, new_G1955gat_,
    new_G1959gat_, new_G1963gat_, new_G1967gat_, new_G1971gat_,
    new_G1975gat_, new_G1979gat_, new_G1983gat_, new_G1987gat_,
    new_G1991gat_, new_G1995gat_, new_G1999gat_, new_G2000gat_,
    new_G2001gat_, new_G2004gat_, new_G2005gat_, new_G2006gat_,
    new_G2007gat_, new_G2008gat_, new_G2009gat_, new_G2010gat_,
    new_G2011gat_, new_G2012gat_, new_G2013gat_, new_G2014gat_,
    new_G2015gat_, new_G2016gat_, new_G2017gat_, new_G2018gat_,
    new_G2019gat_, new_G2020gat_, new_G2021gat_, new_G2022gat_,
    new_G2023gat_, new_G2024gat_, new_G2025gat_, new_G2026gat_,
    new_G2027gat_, new_G2028gat_, new_G2029gat_, new_G2030gat_,
    new_G2033gat_, new_G2037gat_, new_G2040gat_, new_G2043gat_,
    new_G2046gat_, new_G2049gat_, new_G2052gat_, new_G2055gat_,
    new_G2058gat_, new_G2061gat_, new_G2064gat_, new_G2067gat_,
    new_G2070gat_, new_G2073gat_, new_G2076gat_, new_G2080gat_,
    new_G2081gat_, new_G2082gat_, new_G2085gat_, new_G2089gat_,
    new_G2093gat_, new_G2097gat_, new_G2101gat_, new_G2105gat_,
    new_G2109gat_, new_G2113gat_, new_G2117gat_, new_G2121gat_,
    new_G2125gat_, new_G2129gat_, new_G2133gat_, new_G2137gat_,
    new_G2138gat_, new_G2139gat_, new_G2142gat_, new_G2145gat_,
    new_G2149gat_, new_G2150gat_, new_G2151gat_, new_G2154gat_,
    new_G2155gat_, new_G2156gat_, new_G2159gat_, new_G2160gat_,
    new_G2161gat_, new_G2164gat_, new_G2165gat_, new_G2166gat_,
    new_G2169gat_, new_G2170gat_, new_G2171gat_, new_G2174gat_,
    new_G2175gat_, new_G2176gat_, new_G2179gat_, new_G2180gat_,
    new_G2181gat_, new_G2184gat_, new_G2185gat_, new_G2186gat_,
    new_G2189gat_, new_G2190gat_, new_G2191gat_, new_G2194gat_,
    new_G2195gat_, new_G2196gat_, new_G2199gat_, new_G2200gat_,
    new_G2201gat_, new_G2204gat_, new_G2205gat_, new_G2206gat_,
    new_G2209gat_, new_G2210gat_, new_G2211gat_, new_G2214gat_,
    new_G2217gat_, new_G2221gat_, new_G2222gat_, new_G2224gat_,
    new_G2227gat_, new_G2230gat_, new_G2233gat_, new_G2236gat_,
    new_G2239gat_, new_G2242gat_, new_G2245gat_, new_G2248gat_,
    new_G2251gat_, new_G2254gat_, new_G2257gat_, new_G2260gat_,
    new_G2264gat_, new_G2265gat_, new_G2266gat_, new_G2269gat_,
    new_G2273gat_, new_G2277gat_, new_G2281gat_, new_G2285gat_,
    new_G2289gat_, new_G2293gat_, new_G2297gat_, new_G2301gat_,
    new_G2305gat_, new_G2309gat_, new_G2313gat_, new_G2317gat_,
    new_G2318gat_, new_G2319gat_, new_G2322gat_, new_G2326gat_,
    new_G2327gat_, new_G2328gat_, new_G2329gat_, new_G2330gat_,
    new_G2331gat_, new_G2332gat_, new_G2333gat_, new_G2334gat_,
    new_G2335gat_, new_G2336gat_, new_G2337gat_, new_G2338gat_,
    new_G2339gat_, new_G2340gat_, new_G2341gat_, new_G2342gat_,
    new_G2343gat_, new_G2344gat_, new_G2345gat_, new_G2346gat_,
    new_G2347gat_, new_G2348gat_, new_G2349gat_, new_G2350gat_,
    new_G2353gat_, new_G2357gat_, new_G2358gat_, new_G2359gat_,
    new_G2362gat_, new_G2365gat_, new_G2368gat_, new_G2371gat_,
    new_G2374gat_, new_G2377gat_, new_G2380gat_, new_G2383gat_,
    new_G2386gat_, new_G2389gat_, new_G2392gat_, new_G2395gat_,
    new_G2398gat_, new_G2402gat_, new_G2403gat_, new_G2404gat_,
    new_G2407gat_, new_G2410gat_, new_G2414gat_, new_G2418gat_,
    new_G2422gat_, new_G2426gat_, new_G2430gat_, new_G2434gat_,
    new_G2438gat_, new_G2442gat_, new_G2446gat_, new_G2450gat_,
    new_G2454gat_, new_G2458gat_, new_G2462gat_, new_G2463gat_,
    new_G2464gat_, new_G2467gat_, new_G2470gat_, new_G2474gat_,
    new_G2475gat_, new_G2476gat_, new_G2477gat_, new_G2478gat_,
    new_G2481gat_, new_G2482gat_, new_G2483gat_, new_G2486gat_,
    new_G2487gat_, new_G2488gat_, new_G2491gat_, new_G2492gat_,
    new_G2493gat_, new_G2496gat_, new_G2497gat_, new_G2498gat_,
    new_G2501gat_, new_G2502gat_, new_G2503gat_, new_G2506gat_,
    new_G2507gat_, new_G2508gat_, new_G2511gat_, new_G2512gat_,
    new_G2513gat_, new_G2516gat_, new_G2517gat_, new_G2518gat_,
    new_G2521gat_, new_G2522gat_, new_G2523gat_, new_G2526gat_,
    new_G2527gat_, new_G2528gat_, new_G2531gat_, new_G2532gat_,
    new_G2533gat_, new_G2536gat_, new_G2539gat_, new_G2543gat_,
    new_G2544gat_, new_G2545gat_, new_G2549gat_, new_G2552gat_,
    new_G2555gat_, new_G2558gat_, new_G2561gat_, new_G2564gat_,
    new_G2567gat_, new_G2570gat_, new_G2573gat_, new_G2576gat_,
    new_G2579gat_, new_G2582gat_, new_G2586gat_, new_G2587gat_,
    new_G2588gat_, new_G2591gat_, new_G2595gat_, new_G2599gat_,
    new_G2603gat_, new_G2607gat_, new_G2611gat_, new_G2615gat_,
    new_G2619gat_, new_G2623gat_, new_G2627gat_, new_G2631gat_,
    new_G2635gat_, new_G2639gat_, new_G2640gat_, new_G2641gat_,
    new_G2644gat_, new_G2648gat_, new_G2649gat_, new_G2650gat_,
    new_G2653gat_, new_G2654gat_, new_G2655gat_, new_G2656gat_,
    new_G2657gat_, new_G2658gat_, new_G2659gat_, new_G2660gat_,
    new_G2661gat_, new_G2662gat_, new_G2663gat_, new_G2664gat_,
    new_G2665gat_, new_G2666gat_, new_G2667gat_, new_G2668gat_,
    new_G2669gat_, new_G2670gat_, new_G2671gat_, new_G2672gat_,
    new_G2673gat_, new_G2674gat_, new_G2675gat_, new_G2678gat_,
    new_G2682gat_, new_G2683gat_, new_G2684gat_, new_G2687gat_,
    new_G2690gat_, new_G2694gat_, new_G2697gat_, new_G2700gat_,
    new_G2703gat_, new_G2706gat_, new_G2709gat_, new_G2712gat_,
    new_G2715gat_, new_G2718gat_, new_G2721gat_, new_G2724gat_,
    new_G2727gat_, new_G2731gat_, new_G2732gat_, new_G2733gat_,
    new_G2736gat_, new_G2739gat_, new_G2743gat_, new_G2744gat_,
    new_G2745gat_, new_G2749gat_, new_G2753gat_, new_G2757gat_,
    new_G2761gat_, new_G2765gat_, new_G2769gat_, new_G2773gat_,
    new_G2777gat_, new_G2781gat_, new_G2785gat_, new_G2789gat_,
    new_G2790gat_, new_G2791gat_, new_G2794gat_, new_G2797gat_,
    new_G2801gat_, new_G2802gat_, new_G2803gat_, new_G2806gat_,
    new_G2807gat_, new_G2808gat_, new_G2811gat_, new_G2812gat_,
    new_G2813gat_, new_G2816gat_, new_G2817gat_, new_G2818gat_,
    new_G2821gat_, new_G2822gat_, new_G2823gat_, new_G2826gat_,
    new_G2827gat_, new_G2828gat_, new_G2831gat_, new_G2832gat_,
    new_G2833gat_, new_G2836gat_, new_G2837gat_, new_G2838gat_,
    new_G2841gat_, new_G2842gat_, new_G2843gat_, new_G2846gat_,
    new_G2847gat_, new_G2848gat_, new_G2851gat_, new_G2852gat_,
    new_G2853gat_, new_G2856gat_, new_G2857gat_, new_G2858gat_,
    new_G2861gat_, new_G2864gat_, new_G2868gat_, new_G2869gat_,
    new_G2870gat_, new_G2873gat_, new_G2878gat_, new_G2881gat_,
    new_G2884gat_, new_G2887gat_, new_G2890gat_, new_G2893gat_,
    new_G2896gat_, new_G2899gat_, new_G2902gat_, new_G2905gat_,
    new_G2908gat_, new_G2912gat_, new_G2913gat_, new_G2914gat_,
    new_G2917gat_, new_G2921gat_, new_G2922gat_, new_G2923gat_,
    new_G2926gat_, new_G2930gat_, new_G2934gat_, new_G2938gat_,
    new_G2942gat_, new_G2946gat_, new_G2950gat_, new_G2954gat_,
    new_G2958gat_, new_G2962gat_, new_G2966gat_, new_G2967gat_,
    new_G2968gat_, new_G2971gat_, new_G2975gat_, new_G2976gat_,
    new_G2977gat_, new_G2980gat_, new_G2983gat_, new_G2987gat_,
    new_G2988gat_, new_G2989gat_, new_G2990gat_, new_G2991gat_,
    new_G2992gat_, new_G2993gat_, new_G2994gat_, new_G2995gat_,
    new_G2996gat_, new_G2997gat_, new_G2998gat_, new_G2999gat_,
    new_G3000gat_, new_G3001gat_, new_G3002gat_, new_G3003gat_,
    new_G3004gat_, new_G3005gat_, new_G3006gat_, new_G3007gat_,
    new_G3010gat_, new_G3014gat_, new_G3015gat_, new_G3016gat_,
    new_G3019gat_, new_G3022gat_, new_G3026gat_, new_G3027gat_,
    new_G3028gat_, new_G3031gat_, new_G3034gat_, new_G3037gat_,
    new_G3040gat_, new_G3043gat_, new_G3046gat_, new_G3049gat_,
    new_G3052gat_, new_G3055gat_, new_G3058gat_, new_G3062gat_,
    new_G3063gat_, new_G3064gat_, new_G3067gat_, new_G3070gat_,
    new_G3074gat_, new_G3075gat_, new_G3076gat_, new_G3079gat_,
    new_G3083gat_, new_G3087gat_, new_G3091gat_, new_G3095gat_,
    new_G3099gat_, new_G3103gat_, new_G3107gat_, new_G3111gat_,
    new_G3115gat_, new_G3119gat_, new_G3120gat_, new_G3121gat_,
    new_G3124gat_, new_G3127gat_, new_G3131gat_, new_G3132gat_,
    new_G3133gat_, new_G3136gat_, new_G3140gat_, new_G3141gat_,
    new_G3142gat_, new_G3145gat_, new_G3146gat_, new_G3147gat_,
    new_G3150gat_, new_G3151gat_, new_G3152gat_, new_G3155gat_,
    new_G3156gat_, new_G3157gat_, new_G3160gat_, new_G3161gat_,
    new_G3162gat_, new_G3165gat_, new_G3166gat_, new_G3167gat_,
    new_G3170gat_, new_G3171gat_, new_G3172gat_, new_G3175gat_,
    new_G3176gat_, new_G3177gat_, new_G3180gat_, new_G3181gat_,
    new_G3182gat_, new_G3185gat_, new_G3186gat_, new_G3187gat_,
    new_G3190gat_, new_G3193gat_, new_G3197gat_, new_G3198gat_,
    new_G3199gat_, new_G3202gat_, new_G3206gat_, new_G3207gat_,
    new_G3208gat_, new_G3212gat_, new_G3215gat_, new_G3218gat_,
    new_G3221gat_, new_G3224gat_, new_G3227gat_, new_G3230gat_,
    new_G3233gat_, new_G3236gat_, new_G3239gat_, new_G3243gat_,
    new_G3244gat_, new_G3245gat_, new_G3248gat_, new_G3252gat_,
    new_G3253gat_, new_G3254gat_, new_G3257gat_, new_G3260gat_,
    new_G3264gat_, new_G3268gat_, new_G3272gat_, new_G3276gat_,
    new_G3280gat_, new_G3284gat_, new_G3288gat_, new_G3292gat_,
    new_G3296gat_, new_G3300gat_, new_G3301gat_, new_G3302gat_,
    new_G3305gat_, new_G3309gat_, new_G3310gat_, new_G3311gat_,
    new_G3314gat_, new_G3317gat_, new_G3321gat_, new_G3322gat_,
    new_G3323gat_, new_G3324gat_, new_G3325gat_, new_G3326gat_,
    new_G3327gat_, new_G3328gat_, new_G3329gat_, new_G3330gat_,
    new_G3331gat_, new_G3332gat_, new_G3333gat_, new_G3334gat_,
    new_G3335gat_, new_G3336gat_, new_G3337gat_, new_G3338gat_,
    new_G3339gat_, new_G3340gat_, new_G3341gat_, new_G3344gat_,
    new_G3348gat_, new_G3349gat_, new_G3350gat_, new_G3353gat_,
    new_G3356gat_, new_G3360gat_, new_G3361gat_, new_G3362gat_,
    new_G3365gat_, new_G3368gat_, new_G3371gat_, new_G3374gat_,
    new_G3377gat_, new_G3380gat_, new_G3383gat_, new_G3386gat_,
    new_G3389gat_, new_G3392gat_, new_G3396gat_, new_G3397gat_,
    new_G3398gat_, new_G3401gat_, new_G3404gat_, new_G3408gat_,
    new_G3409gat_, new_G3410gat_, new_G3413gat_, new_G3417gat_,
    new_G3421gat_, new_G3425gat_, new_G3429gat_, new_G3433gat_,
    new_G3437gat_, new_G3441gat_, new_G3445gat_, new_G3449gat_,
    new_G3453gat_, new_G3454gat_, new_G3455gat_, new_G3458gat_,
    new_G3461gat_, new_G3465gat_, new_G3466gat_, new_G3467gat_,
    new_G3470gat_, new_G3474gat_, new_G3475gat_, new_G3476gat_,
    new_G3479gat_, new_G3480gat_, new_G3481gat_, new_G3484gat_,
    new_G3485gat_, new_G3486gat_, new_G3489gat_, new_G3490gat_,
    new_G3491gat_, new_G3494gat_, new_G3495gat_, new_G3496gat_,
    new_G3499gat_, new_G3500gat_, new_G3501gat_, new_G3504gat_,
    new_G3505gat_, new_G3506gat_, new_G3509gat_, new_G3510gat_,
    new_G3511gat_, new_G3514gat_, new_G3515gat_, new_G3516gat_,
    new_G3519gat_, new_G3520gat_, new_G3521gat_, new_G3524gat_,
    new_G3527gat_, new_G3531gat_, new_G3532gat_, new_G3533gat_,
    new_G3536gat_, new_G3540gat_, new_G3541gat_, new_G3542gat_,
    new_G3545gat_, new_G3548gat_, new_G3553gat_, new_G3556gat_,
    new_G3559gat_, new_G3562gat_, new_G3565gat_, new_G3568gat_,
    new_G3571gat_, new_G3574gat_, new_G3577gat_, new_G3581gat_,
    new_G3582gat_, new_G3583gat_, new_G3586gat_, new_G3590gat_,
    new_G3591gat_, new_G3592gat_, new_G3595gat_, new_G3598gat_,
    new_G3602gat_, new_G3603gat_, new_G3604gat_, new_G3608gat_,
    new_G3612gat_, new_G3616gat_, new_G3620gat_, new_G3624gat_,
    new_G3628gat_, new_G3632gat_, new_G3636gat_, new_G3637gat_,
    new_G3638gat_, new_G3641gat_, new_G3645gat_, new_G3646gat_,
    new_G3647gat_, new_G3650gat_, new_G3653gat_, new_G3657gat_,
    new_G3658gat_, new_G3659gat_, new_G3662gat_, new_G3663gat_,
    new_G3664gat_, new_G3665gat_, new_G3666gat_, new_G3667gat_,
    new_G3668gat_, new_G3669gat_, new_G3670gat_, new_G3671gat_,
    new_G3672gat_, new_G3673gat_, new_G3674gat_, new_G3675gat_,
    new_G3676gat_, new_G3677gat_, new_G3678gat_, new_G3681gat_,
    new_G3685gat_, new_G3686gat_, new_G3687gat_, new_G3690gat_,
    new_G3693gat_, new_G3697gat_, new_G3698gat_, new_G3699gat_,
    new_G3702gat_, new_G3706gat_, new_G3709gat_, new_G3712gat_,
    new_G3715gat_, new_G3718gat_, new_G3721gat_, new_G3724gat_,
    new_G3727gat_, new_G3730gat_, new_G3734gat_, new_G3735gat_,
    new_G3736gat_, new_G3739gat_, new_G3742gat_, new_G3746gat_,
    new_G3747gat_, new_G3748gat_, new_G3751gat_, new_G3755gat_,
    new_G3756gat_, new_G3757gat_, new_G3760gat_, new_G3764gat_,
    new_G3768gat_, new_G3772gat_, new_G3776gat_, new_G3780gat_,
    new_G3784gat_, new_G3788gat_, new_G3792gat_, new_G3793gat_,
    new_G3794gat_, new_G3797gat_, new_G3800gat_, new_G3804gat_,
    new_G3805gat_, new_G3806gat_, new_G3809gat_, new_G3813gat_,
    new_G3814gat_, new_G3815gat_, new_G3818gat_, new_G3821gat_,
    new_G3825gat_, new_G3826gat_, new_G3827gat_, new_G3830gat_,
    new_G3831gat_, new_G3832gat_, new_G3835gat_, new_G3836gat_,
    new_G3837gat_, new_G3840gat_, new_G3841gat_, new_G3842gat_,
    new_G3845gat_, new_G3846gat_, new_G3847gat_, new_G3850gat_,
    new_G3851gat_, new_G3852gat_, new_G3855gat_, new_G3856gat_,
    new_G3857gat_, new_G3860gat_, new_G3861gat_, new_G3862gat_,
    new_G3865gat_, new_G3868gat_, new_G3872gat_, new_G3873gat_,
    new_G3874gat_, new_G3877gat_, new_G3881gat_, new_G3882gat_,
    new_G3883gat_, new_G3886gat_, new_G3889gat_, new_G3893gat_,
    new_G3894gat_, new_G3896gat_, new_G3899gat_, new_G3902gat_,
    new_G3905gat_, new_G3908gat_, new_G3911gat_, new_G3914gat_,
    new_G3917gat_, new_G3921gat_, new_G3922gat_, new_G3923gat_,
    new_G3926gat_, new_G3930gat_, new_G3931gat_, new_G3932gat_,
    new_G3935gat_, new_G3938gat_, new_G3942gat_, new_G3943gat_,
    new_G3944gat_, new_G3947gat_, new_G3951gat_, new_G3955gat_,
    new_G3959gat_, new_G3963gat_, new_G3967gat_, new_G3971gat_,
    new_G3975gat_, new_G3976gat_, new_G3977gat_, new_G3980gat_,
    new_G3984gat_, new_G3985gat_, new_G3986gat_, new_G3989gat_,
    new_G3992gat_, new_G3996gat_, new_G3997gat_, new_G3998gat_,
    new_G4001gat_, new_G4005gat_, new_G4006gat_, new_G4007gat_,
    new_G4008gat_, new_G4009gat_, new_G4010gat_, new_G4011gat_,
    new_G4012gat_, new_G4013gat_, new_G4014gat_, new_G4015gat_,
    new_G4016gat_, new_G4017gat_, new_G4018gat_, new_G4019gat_,
    new_G4022gat_, new_G4026gat_, new_G4027gat_, new_G4028gat_,
    new_G4031gat_, new_G4034gat_, new_G4038gat_, new_G4039gat_,
    new_G4040gat_, new_G4043gat_, new_G4047gat_, new_G4048gat_,
    new_G4049gat_, new_G4052gat_, new_G4055gat_, new_G4058gat_,
    new_G4061gat_, new_G4064gat_, new_G4067gat_, new_G4070gat_,
    new_G4073gat_, new_G4077gat_, new_G4078gat_, new_G4079gat_,
    new_G4082gat_, new_G4085gat_, new_G4089gat_, new_G4090gat_,
    new_G4091gat_, new_G4094gat_, new_G4098gat_, new_G4099gat_,
    new_G4100gat_, new_G4103gat_, new_G4106gat_, new_G4110gat_,
    new_G4114gat_, new_G4118gat_, new_G4122gat_, new_G4126gat_,
    new_G4130gat_, new_G4134gat_, new_G4138gat_, new_G4139gat_,
    new_G4140gat_, new_G4143gat_, new_G4146gat_, new_G4150gat_,
    new_G4151gat_, new_G4152gat_, new_G4155gat_, new_G4159gat_,
    new_G4160gat_, new_G4161gat_, new_G4164gat_, new_G4167gat_,
    new_G4171gat_, new_G4172gat_, new_G4173gat_, new_G4174gat_,
    new_G4175gat_, new_G4178gat_, new_G4179gat_, new_G4180gat_,
    new_G4183gat_, new_G4184gat_, new_G4185gat_, new_G4188gat_,
    new_G4189gat_, new_G4190gat_, new_G4193gat_, new_G4194gat_,
    new_G4195gat_, new_G4198gat_, new_G4199gat_, new_G4200gat_,
    new_G4203gat_, new_G4204gat_, new_G4205gat_, new_G4208gat_,
    new_G4211gat_, new_G4215gat_, new_G4216gat_, new_G4217gat_,
    new_G4220gat_, new_G4224gat_, new_G4225gat_, new_G4226gat_,
    new_G4229gat_, new_G4232gat_, new_G4236gat_, new_G4237gat_,
    new_G4238gat_, new_G4242gat_, new_G4245gat_, new_G4248gat_,
    new_G4251gat_, new_G4254gat_, new_G4257gat_, new_G4260gat_,
    new_G4264gat_, new_G4265gat_, new_G4266gat_, new_G4269gat_,
    new_G4273gat_, new_G4274gat_, new_G4275gat_, new_G4278gat_,
    new_G4281gat_, new_G4285gat_, new_G4286gat_, new_G4287gat_,
    new_G4290gat_, new_G4294gat_, new_G4298gat_, new_G4302gat_,
    new_G4306gat_, new_G4310gat_, new_G4314gat_, new_G4318gat_,
    new_G4319gat_, new_G4320gat_, new_G4323gat_, new_G4327gat_,
    new_G4328gat_, new_G4329gat_, new_G4332gat_, new_G4335gat_,
    new_G4339gat_, new_G4340gat_, new_G4341gat_, new_G4344gat_,
    new_G4348gat_, new_G4349gat_, new_G4350gat_, new_G4353gat_,
    new_G4354gat_, new_G4355gat_, new_G4356gat_, new_G4357gat_,
    new_G4358gat_, new_G4359gat_, new_G4360gat_, new_G4361gat_,
    new_G4362gat_, new_G4363gat_, new_G4364gat_, new_G4365gat_,
    new_G4368gat_, new_G4372gat_, new_G4373gat_, new_G4374gat_,
    new_G4377gat_, new_G4380gat_, new_G4384gat_, new_G4385gat_,
    new_G4386gat_, new_G4389gat_, new_G4393gat_, new_G4394gat_,
    new_G4395gat_, new_G4398gat_, new_G4401gat_, new_G4405gat_,
    new_G4408gat_, new_G4411gat_, new_G4414gat_, new_G4417gat_,
    new_G4420gat_, new_G4423gat_, new_G4427gat_, new_G4428gat_,
    new_G4429gat_, new_G4432gat_, new_G4435gat_, new_G4439gat_,
    new_G4440gat_, new_G4441gat_, new_G4444gat_, new_G4448gat_,
    new_G4449gat_, new_G4450gat_, new_G4453gat_, new_G4456gat_,
    new_G4460gat_, new_G4461gat_, new_G4462gat_, new_G4466gat_,
    new_G4470gat_, new_G4474gat_, new_G4478gat_, new_G4482gat_,
    new_G4486gat_, new_G4487gat_, new_G4488gat_, new_G4491gat_,
    new_G4494gat_, new_G4498gat_, new_G4499gat_, new_G4500gat_,
    new_G4503gat_, new_G4507gat_, new_G4508gat_, new_G4509gat_,
    new_G4512gat_, new_G4515gat_, new_G4519gat_, new_G4520gat_,
    new_G4521gat_, new_G4524gat_, new_G4525gat_, new_G4526gat_,
    new_G4529gat_, new_G4530gat_, new_G4531gat_, new_G4534gat_,
    new_G4535gat_, new_G4536gat_, new_G4539gat_, new_G4540gat_,
    new_G4541gat_, new_G4544gat_, new_G4545gat_, new_G4546gat_,
    new_G4549gat_, new_G4550gat_, new_G4551gat_, new_G4554gat_,
    new_G4557gat_, new_G4561gat_, new_G4562gat_, new_G4563gat_,
    new_G4566gat_, new_G4570gat_, new_G4571gat_, new_G4572gat_,
    new_G4575gat_, new_G4578gat_, new_G4582gat_, new_G4583gat_,
    new_G4584gat_, new_G4587gat_, new_G4592gat_, new_G4595gat_,
    new_G4598gat_, new_G4601gat_, new_G4604gat_, new_G4607gat_,
    new_G4611gat_, new_G4612gat_, new_G4613gat_, new_G4616gat_,
    new_G4620gat_, new_G4621gat_, new_G4622gat_, new_G4625gat_,
    new_G4628gat_, new_G4632gat_, new_G4633gat_, new_G4634gat_,
    new_G4637gat_, new_G4641gat_, new_G4642gat_, new_G4643gat_,
    new_G4646gat_, new_G4650gat_, new_G4654gat_, new_G4658gat_,
    new_G4662gat_, new_G4666gat_, new_G4667gat_, new_G4668gat_,
    new_G4671gat_, new_G4675gat_, new_G4676gat_, new_G4677gat_,
    new_G4680gat_, new_G4683gat_, new_G4687gat_, new_G4688gat_,
    new_G4689gat_, new_G4692gat_, new_G4696gat_, new_G4697gat_,
    new_G4698gat_, new_G4701gat_, new_G4704gat_, new_G4708gat_,
    new_G4709gat_, new_G4710gat_, new_G4711gat_, new_G4712gat_,
    new_G4713gat_, new_G4714gat_, new_G4715gat_, new_G4716gat_,
    new_G4717gat_, new_G4718gat_, new_G4721gat_, new_G4725gat_,
    new_G4726gat_, new_G4727gat_, new_G4730gat_, new_G4733gat_,
    new_G4737gat_, new_G4738gat_, new_G4739gat_, new_G4742gat_,
    new_G4746gat_, new_G4747gat_, new_G4748gat_, new_G4751gat_,
    new_G4754gat_, new_G4758gat_, new_G4759gat_, new_G4760gat_,
    new_G4763gat_, new_G4766gat_, new_G4769gat_, new_G4772gat_,
    new_G4775gat_, new_G4779gat_, new_G4780gat_, new_G4781gat_,
    new_G4784gat_, new_G4787gat_, new_G4791gat_, new_G4792gat_,
    new_G4793gat_, new_G4796gat_, new_G4800gat_, new_G4801gat_,
    new_G4802gat_, new_G4805gat_, new_G4808gat_, new_G4812gat_,
    new_G4813gat_, new_G4814gat_, new_G4817gat_, new_G4821gat_,
    new_G4825gat_, new_G4829gat_, new_G4833gat_, new_G4837gat_,
    new_G4838gat_, new_G4839gat_, new_G4842gat_, new_G4845gat_,
    new_G4849gat_, new_G4850gat_, new_G4851gat_, new_G4854gat_,
    new_G4858gat_, new_G4859gat_, new_G4860gat_, new_G4863gat_,
    new_G4866gat_, new_G4870gat_, new_G4871gat_, new_G4872gat_,
    new_G4875gat_, new_G4879gat_, new_G4880gat_, new_G4881gat_,
    new_G4884gat_, new_G4885gat_, new_G4886gat_, new_G4889gat_,
    new_G4890gat_, new_G4891gat_, new_G4894gat_, new_G4895gat_,
    new_G4896gat_, new_G4899gat_, new_G4900gat_, new_G4901gat_,
    new_G4904gat_, new_G4907gat_, new_G4911gat_, new_G4912gat_,
    new_G4913gat_, new_G4916gat_, new_G4920gat_, new_G4921gat_,
    new_G4922gat_, new_G4925gat_, new_G4928gat_, new_G4932gat_,
    new_G4933gat_, new_G4934gat_, new_G4937gat_, new_G4941gat_,
    new_G4942gat_, new_G4943gat_, new_G4947gat_, new_G4950gat_,
    new_G4953gat_, new_G4956gat_, new_G4959gat_, new_G4963gat_,
    new_G4964gat_, new_G4965gat_, new_G4968gat_, new_G4972gat_,
    new_G4973gat_, new_G4974gat_, new_G4977gat_, new_G4980gat_,
    new_G4984gat_, new_G4985gat_, new_G4986gat_, new_G4989gat_,
    new_G4993gat_, new_G4994gat_, new_G4995gat_, new_G4998gat_,
    new_G5001gat_, new_G5005gat_, new_G5009gat_, new_G5013gat_,
    new_G5017gat_, new_G5021gat_, new_G5022gat_, new_G5023gat_,
    new_G5026gat_, new_G5030gat_, new_G5031gat_, new_G5032gat_,
    new_G5035gat_, new_G5038gat_, new_G5042gat_, new_G5043gat_,
    new_G5044gat_, new_G5047gat_, new_G5051gat_, new_G5052gat_,
    new_G5053gat_, new_G5056gat_, new_G5059gat_, new_G5063gat_,
    new_G5064gat_, new_G5065gat_, new_G5066gat_, new_G5067gat_,
    new_G5068gat_, new_G5069gat_, new_G5070gat_, new_G5071gat_,
    new_G5072gat_, new_G5073gat_, new_G5076gat_, new_G5080gat_,
    new_G5081gat_, new_G5082gat_, new_G5085gat_, new_G5088gat_,
    new_G5092gat_, new_G5093gat_, new_G5094gat_, new_G5097gat_,
    new_G5101gat_, new_G5102gat_, new_G5103gat_, new_G5106gat_,
    new_G5109gat_, new_G5113gat_, new_G5114gat_, new_G5115gat_,
    new_G5118gat_, new_G5121gat_, new_G5124gat_, new_G5127gat_,
    new_G5130gat_, new_G5134gat_, new_G5135gat_, new_G5136gat_,
    new_G5139gat_, new_G5142gat_, new_G5146gat_, new_G5147gat_,
    new_G5148gat_, new_G5151gat_, new_G5155gat_, new_G5156gat_,
    new_G5157gat_, new_G5160gat_, new_G5163gat_, new_G5167gat_,
    new_G5168gat_, new_G5169gat_, new_G5172gat_, new_G5176gat_,
    new_G5180gat_, new_G5184gat_, new_G5188gat_, new_G5192gat_,
    new_G5193gat_, new_G5194gat_, new_G5197gat_, new_G5200gat_,
    new_G5204gat_, new_G5205gat_, new_G5206gat_, new_G5209gat_,
    new_G5213gat_, new_G5214gat_, new_G5215gat_, new_G5218gat_,
    new_G5221gat_, new_G5225gat_, new_G5226gat_, new_G5227gat_,
    new_G5230gat_, new_G5234gat_, new_G5235gat_, new_G5236gat_,
    new_G5239gat_, new_G5240gat_, new_G5241gat_, new_G5244gat_,
    new_G5245gat_, new_G5246gat_, new_G5249gat_, new_G5250gat_,
    new_G5251gat_, new_G5254gat_, new_G5255gat_, new_G5256gat_,
    new_G5259gat_, new_G5262gat_, new_G5266gat_, new_G5267gat_,
    new_G5268gat_, new_G5271gat_, new_G5275gat_, new_G5276gat_,
    new_G5277gat_, new_G5280gat_, new_G5283gat_, new_G5287gat_,
    new_G5288gat_, new_G5289gat_, new_G5292gat_, new_G5296gat_,
    new_G5297gat_, new_G5298gat_, new_G5301gat_, new_G5304gat_,
    new_G5309gat_, new_G5312gat_, new_G5315gat_, new_G5318gat_,
    new_G5322gat_, new_G5323gat_, new_G5324gat_, new_G5327gat_,
    new_G5331gat_, new_G5332gat_, new_G5333gat_, new_G5336gat_,
    new_G5339gat_, new_G5343gat_, new_G5344gat_, new_G5345gat_,
    new_G5348gat_, new_G5352gat_, new_G5353gat_, new_G5354gat_,
    new_G5357gat_, new_G5360gat_, new_G5364gat_, new_G5365gat_,
    new_G5366gat_, new_G5370gat_, new_G5374gat_, new_G5378gat_,
    new_G5379gat_, new_G5380gat_, new_G5383gat_, new_G5387gat_,
    new_G5388gat_, new_G5389gat_, new_G5392gat_, new_G5395gat_,
    new_G5399gat_, new_G5400gat_, new_G5401gat_, new_G5404gat_,
    new_G5408gat_, new_G5409gat_, new_G5410gat_, new_G5413gat_,
    new_G5416gat_, new_G5420gat_, new_G5421gat_, new_G5422gat_,
    new_G5425gat_, new_G5426gat_, new_G5427gat_, new_G5428gat_,
    new_G5429gat_, new_G5430gat_, new_G5431gat_, new_G5434gat_,
    new_G5438gat_, new_G5439gat_, new_G5440gat_, new_G5443gat_,
    new_G5446gat_, new_G5450gat_, new_G5451gat_, new_G5452gat_,
    new_G5455gat_, new_G5459gat_, new_G5460gat_, new_G5461gat_,
    new_G5464gat_, new_G5467gat_, new_G5471gat_, new_G5472gat_,
    new_G5473gat_, new_G5476gat_, new_G5480gat_, new_G5483gat_,
    new_G5486gat_, new_G5489gat_, new_G5493gat_, new_G5494gat_,
    new_G5495gat_, new_G5498gat_, new_G5501gat_, new_G5505gat_,
    new_G5506gat_, new_G5507gat_, new_G5510gat_, new_G5514gat_,
    new_G5515gat_, new_G5516gat_, new_G5519gat_, new_G5522gat_,
    new_G5526gat_, new_G5527gat_, new_G5528gat_, new_G5531gat_,
    new_G5535gat_, new_G5536gat_, new_G5537gat_, new_G5540gat_,
    new_G5544gat_, new_G5548gat_, new_G5552gat_, new_G5553gat_,
    new_G5554gat_, new_G5557gat_, new_G5560gat_, new_G5564gat_,
    new_G5565gat_, new_G5566gat_, new_G5569gat_, new_G5573gat_,
    new_G5574gat_, new_G5575gat_, new_G5578gat_, new_G5581gat_,
    new_G5585gat_, new_G5586gat_, new_G5587gat_, new_G5590gat_,
    new_G5594gat_, new_G5595gat_, new_G5596gat_, new_G5599gat_,
    new_G5602gat_, new_G5606gat_, new_G5607gat_, new_G5608gat_,
    new_G5611gat_, new_G5612gat_, new_G5613gat_, new_G5616gat_,
    new_G5617gat_, new_G5618gat_, new_G5621gat_, new_G5624gat_,
    new_G5628gat_, new_G5629gat_, new_G5630gat_, new_G5633gat_,
    new_G5637gat_, new_G5638gat_, new_G5639gat_, new_G5642gat_,
    new_G5645gat_, new_G5649gat_, new_G5650gat_, new_G5651gat_,
    new_G5654gat_, new_G5658gat_, new_G5659gat_, new_G5660gat_,
    new_G5663gat_, new_G5666gat_, new_G5670gat_, new_G5671gat_,
    new_G5673gat_, new_G5676gat_, new_G5679gat_, new_G5683gat_,
    new_G5684gat_, new_G5685gat_, new_G5688gat_, new_G5692gat_,
    new_G5693gat_, new_G5694gat_, new_G5697gat_, new_G5700gat_,
    new_G5704gat_, new_G5705gat_, new_G5706gat_, new_G5709gat_,
    new_G5713gat_, new_G5714gat_, new_G5715gat_, new_G5718gat_,
    new_G5721gat_, new_G5725gat_, new_G5726gat_, new_G5727gat_,
    new_G5730gat_, new_G5734gat_, new_G5738gat_, new_G5739gat_,
    new_G5740gat_, new_G5743gat_, new_G5747gat_, new_G5748gat_,
    new_G5749gat_, new_G5752gat_, new_G5755gat_, new_G5759gat_,
    new_G5760gat_, new_G5761gat_, new_G5764gat_, new_G5768gat_,
    new_G5769gat_, new_G5770gat_, new_G5773gat_, new_G5776gat_,
    new_G5780gat_, new_G5781gat_, new_G5782gat_, new_G5785gat_,
    new_G5786gat_, new_G5787gat_, new_G5788gat_, new_G5789gat_,
    new_G5792gat_, new_G5796gat_, new_G5797gat_, new_G5798gat_,
    new_G5801gat_, new_G5804gat_, new_G5808gat_, new_G5809gat_,
    new_G5810gat_, new_G5813gat_, new_G5817gat_, new_G5818gat_,
    new_G5819gat_, new_G5822gat_, new_G5825gat_, new_G5829gat_,
    new_G5830gat_, new_G5831gat_, new_G5834gat_, new_G5837gat_,
    new_G5840gat_, new_G5844gat_, new_G5845gat_, new_G5846gat_,
    new_G5849gat_, new_G5852gat_, new_G5856gat_, new_G5857gat_,
    new_G5858gat_, new_G5861gat_, new_G5865gat_, new_G5866gat_,
    new_G5867gat_, new_G5870gat_, new_G5873gat_, new_G5877gat_,
    new_G5878gat_, new_G5879gat_, new_G5882gat_, new_G5886gat_,
    new_G5890gat_, new_G5891gat_, new_G5892gat_, new_G5895gat_,
    new_G5898gat_, new_G5902gat_, new_G5903gat_, new_G5904gat_,
    new_G5907gat_, new_G5911gat_, new_G5912gat_, new_G5913gat_,
    new_G5916gat_, new_G5919gat_, new_G5923gat_, new_G5924gat_,
    new_G5925gat_, new_G5928gat_, new_G5929gat_, new_G5930gat_,
    new_G5933gat_, new_G5934gat_, new_G5935gat_, new_G5938gat_,
    new_G5941gat_, new_G5945gat_, new_G5946gat_, new_G5947gat_,
    new_G5950gat_, new_G5954gat_, new_G5955gat_, new_G5956gat_,
    new_G5959gat_, new_G5962gat_, new_G5966gat_, new_G5967gat_,
    new_G5968gat_, new_G5972gat_, new_G5975gat_, new_G5979gat_,
    new_G5980gat_, new_G5981gat_, new_G5984gat_, new_G5988gat_,
    new_G5989gat_, new_G5990gat_, new_G5993gat_, new_G5996gat_,
    new_G6000gat_, new_G6001gat_, new_G6002gat_, new_G6005gat_,
    new_G6009gat_, new_G6010gat_, new_G6011gat_, new_G6014gat_,
    new_G6018gat_, new_G6019gat_, new_G6020gat_, new_G6023gat_,
    new_G6026gat_, new_G6030gat_, new_G6031gat_, new_G6032gat_,
    new_G6035gat_, new_G6036gat_, new_G6037gat_, new_G6040gat_,
    new_G6044gat_, new_G6045gat_, new_G6046gat_, new_G6049gat_,
    new_G6052gat_, new_G6056gat_, new_G6057gat_, new_G6058gat_,
    new_G6061gat_, new_G6064gat_, new_G6068gat_, new_G6069gat_,
    new_G6070gat_, new_G6073gat_, new_G6076gat_, new_G6080gat_,
    new_G6081gat_, new_G6082gat_, new_G6085gat_, new_G6089gat_,
    new_G6090gat_, new_G6091gat_, new_G6094gat_, new_G6097gat_,
    new_G6101gat_, new_G6102gat_, new_G6103gat_, new_G6106gat_,
    new_G6107gat_, new_G6108gat_, new_G6111gat_, new_G6114gat_,
    new_G6118gat_, new_G6119gat_, new_G6120gat_, new_G6124gat_,
    new_G6128gat_, new_G6129gat_, new_G6130gat_, new_G6133gat_,
    new_G6134gat_, new_G6135gat_, new_G6138gat_, new_G6141gat_,
    new_G6145gat_, new_G6146gat_, new_G6147gat_, new_G6151gat_,
    new_G6155gat_, new_G6156gat_, new_G6157gat_, new_G6161gat_,
    new_G6165gat_, new_G6166gat_, new_G6167gat_, new_G6171gat_,
    new_G6175gat_, new_G6176gat_, new_G6177gat_, new_G6181gat_,
    new_G6185gat_, new_G6186gat_, new_G6187gat_, new_G6191gat_,
    new_G6195gat_, new_G6196gat_, new_G6197gat_, new_G6201gat_,
    new_G6205gat_, new_G6206gat_, new_G6207gat_, new_G6211gat_,
    new_G6215gat_, new_G6216gat_, new_G6217gat_, new_G6221gat_,
    new_G6225gat_, new_G6226gat_, new_G6227gat_, new_G6231gat_,
    new_G6235gat_, new_G6236gat_, new_G6237gat_, new_G6241gat_,
    new_G6245gat_, new_G6246gat_, new_G6247gat_, new_G6251gat_,
    new_G6255gat_, new_G6256gat_, new_G6257gat_, new_G6261gat_,
    new_G6265gat_, new_G6266gat_, new_G6267gat_, new_G6271gat_,
    new_G6275gat_, new_G6276gat_, new_G6277gat_, new_G6281gat_,
    new_G6285gat_, new_G6286gat_;
  assign G545gat = G1gat & G273gat;
  assign new_G546gat_ = G1gat & G290gat;
  assign new_G549gat_ = G1gat & G307gat;
  assign new_G552gat_ = G1gat & G324gat;
  assign new_G555gat_ = G1gat & G341gat;
  assign new_G558gat_ = G1gat & G358gat;
  assign new_G561gat_ = G1gat & G375gat;
  assign new_G564gat_ = G1gat & G392gat;
  assign new_G567gat_ = G1gat & G409gat;
  assign new_G570gat_ = G1gat & G426gat;
  assign new_G573gat_ = G1gat & G443gat;
  assign new_G576gat_ = G1gat & G460gat;
  assign new_G579gat_ = G1gat & G477gat;
  assign new_G582gat_ = G1gat & G494gat;
  assign new_G585gat_ = G1gat & G511gat;
  assign new_G588gat_ = G1gat & G528gat;
  assign new_G591gat_ = G18gat & G273gat;
  assign new_G594gat_ = G18gat & G290gat;
  assign new_G597gat_ = G18gat & G307gat;
  assign new_G600gat_ = G18gat & G324gat;
  assign new_G603gat_ = G18gat & G341gat;
  assign new_G606gat_ = G18gat & G358gat;
  assign new_G609gat_ = G18gat & G375gat;
  assign new_G612gat_ = G18gat & G392gat;
  assign new_G615gat_ = G18gat & G409gat;
  assign new_G618gat_ = G18gat & G426gat;
  assign new_G621gat_ = G18gat & G443gat;
  assign new_G624gat_ = G18gat & G460gat;
  assign new_G627gat_ = G18gat & G477gat;
  assign new_G630gat_ = G18gat & G494gat;
  assign new_G633gat_ = G18gat & G511gat;
  assign new_G636gat_ = G18gat & G528gat;
  assign new_G639gat_ = G35gat & G273gat;
  assign new_G642gat_ = G35gat & G290gat;
  assign new_G645gat_ = G35gat & G307gat;
  assign new_G648gat_ = G35gat & G324gat;
  assign new_G651gat_ = G35gat & G341gat;
  assign new_G654gat_ = G35gat & G358gat;
  assign new_G657gat_ = G35gat & G375gat;
  assign new_G660gat_ = G35gat & G392gat;
  assign new_G663gat_ = G35gat & G409gat;
  assign new_G666gat_ = G35gat & G426gat;
  assign new_G669gat_ = G35gat & G443gat;
  assign new_G672gat_ = G35gat & G460gat;
  assign new_G675gat_ = G35gat & G477gat;
  assign new_G678gat_ = G35gat & G494gat;
  assign new_G681gat_ = G35gat & G511gat;
  assign new_G684gat_ = G35gat & G528gat;
  assign new_G687gat_ = G52gat & G273gat;
  assign new_G690gat_ = G52gat & G290gat;
  assign new_G693gat_ = G52gat & G307gat;
  assign new_G696gat_ = G52gat & G324gat;
  assign new_G699gat_ = G52gat & G341gat;
  assign new_G702gat_ = G52gat & G358gat;
  assign new_G705gat_ = G52gat & G375gat;
  assign new_G708gat_ = G52gat & G392gat;
  assign new_G711gat_ = G52gat & G409gat;
  assign new_G714gat_ = G52gat & G426gat;
  assign new_G717gat_ = G52gat & G443gat;
  assign new_G720gat_ = G52gat & G460gat;
  assign new_G723gat_ = G52gat & G477gat;
  assign new_G726gat_ = G52gat & G494gat;
  assign new_G729gat_ = G52gat & G511gat;
  assign new_G732gat_ = G52gat & G528gat;
  assign new_G735gat_ = G69gat & G273gat;
  assign new_G738gat_ = G69gat & G290gat;
  assign new_G741gat_ = G69gat & G307gat;
  assign new_G744gat_ = G69gat & G324gat;
  assign new_G747gat_ = G69gat & G341gat;
  assign new_G750gat_ = G69gat & G358gat;
  assign new_G753gat_ = G69gat & G375gat;
  assign new_G756gat_ = G69gat & G392gat;
  assign new_G759gat_ = G69gat & G409gat;
  assign new_G762gat_ = G69gat & G426gat;
  assign new_G765gat_ = G69gat & G443gat;
  assign new_G768gat_ = G69gat & G460gat;
  assign new_G771gat_ = G69gat & G477gat;
  assign new_G774gat_ = G69gat & G494gat;
  assign new_G777gat_ = G69gat & G511gat;
  assign new_G780gat_ = G69gat & G528gat;
  assign new_G783gat_ = G86gat & G273gat;
  assign new_G786gat_ = G86gat & G290gat;
  assign new_G789gat_ = G86gat & G307gat;
  assign new_G792gat_ = G86gat & G324gat;
  assign new_G795gat_ = G86gat & G341gat;
  assign new_G798gat_ = G86gat & G358gat;
  assign new_G801gat_ = G86gat & G375gat;
  assign new_G804gat_ = G86gat & G392gat;
  assign new_G807gat_ = G86gat & G409gat;
  assign new_G810gat_ = G86gat & G426gat;
  assign new_G813gat_ = G86gat & G443gat;
  assign new_G816gat_ = G86gat & G460gat;
  assign new_G819gat_ = G86gat & G477gat;
  assign new_G822gat_ = G86gat & G494gat;
  assign new_G825gat_ = G86gat & G511gat;
  assign new_G828gat_ = G86gat & G528gat;
  assign new_G831gat_ = G103gat & G273gat;
  assign new_G834gat_ = G103gat & G290gat;
  assign new_G837gat_ = G103gat & G307gat;
  assign new_G840gat_ = G103gat & G324gat;
  assign new_G843gat_ = G103gat & G341gat;
  assign new_G846gat_ = G103gat & G358gat;
  assign new_G849gat_ = G103gat & G375gat;
  assign new_G852gat_ = G103gat & G392gat;
  assign new_G855gat_ = G103gat & G409gat;
  assign new_G858gat_ = G103gat & G426gat;
  assign new_G861gat_ = G103gat & G443gat;
  assign new_G864gat_ = G103gat & G460gat;
  assign new_G867gat_ = G103gat & G477gat;
  assign new_G870gat_ = G103gat & G494gat;
  assign new_G873gat_ = G103gat & G511gat;
  assign new_G876gat_ = G103gat & G528gat;
  assign new_G879gat_ = G120gat & G273gat;
  assign new_G882gat_ = G120gat & G290gat;
  assign new_G885gat_ = G120gat & G307gat;
  assign new_G888gat_ = G120gat & G324gat;
  assign new_G891gat_ = G120gat & G341gat;
  assign new_G894gat_ = G120gat & G358gat;
  assign new_G897gat_ = G120gat & G375gat;
  assign new_G900gat_ = G120gat & G392gat;
  assign new_G903gat_ = G120gat & G409gat;
  assign new_G906gat_ = G120gat & G426gat;
  assign new_G909gat_ = G120gat & G443gat;
  assign new_G912gat_ = G120gat & G460gat;
  assign new_G915gat_ = G120gat & G477gat;
  assign new_G918gat_ = G120gat & G494gat;
  assign new_G921gat_ = G120gat & G511gat;
  assign new_G924gat_ = G120gat & G528gat;
  assign new_G927gat_ = G137gat & G273gat;
  assign new_G930gat_ = G137gat & G290gat;
  assign new_G933gat_ = G137gat & G307gat;
  assign new_G936gat_ = G137gat & G324gat;
  assign new_G939gat_ = G137gat & G341gat;
  assign new_G942gat_ = G137gat & G358gat;
  assign new_G945gat_ = G137gat & G375gat;
  assign new_G948gat_ = G137gat & G392gat;
  assign new_G951gat_ = G137gat & G409gat;
  assign new_G954gat_ = G137gat & G426gat;
  assign new_G957gat_ = G137gat & G443gat;
  assign new_G960gat_ = G137gat & G460gat;
  assign new_G963gat_ = G137gat & G477gat;
  assign new_G966gat_ = G137gat & G494gat;
  assign new_G969gat_ = G137gat & G511gat;
  assign new_G972gat_ = G137gat & G528gat;
  assign new_G975gat_ = G154gat & G273gat;
  assign new_G978gat_ = G154gat & G290gat;
  assign new_G981gat_ = G154gat & G307gat;
  assign new_G984gat_ = G154gat & G324gat;
  assign new_G987gat_ = G154gat & G341gat;
  assign new_G990gat_ = G154gat & G358gat;
  assign new_G993gat_ = G154gat & G375gat;
  assign new_G996gat_ = G154gat & G392gat;
  assign new_G999gat_ = G154gat & G409gat;
  assign new_G1002gat_ = G154gat & G426gat;
  assign new_G1005gat_ = G154gat & G443gat;
  assign new_G1008gat_ = G154gat & G460gat;
  assign new_G1011gat_ = G154gat & G477gat;
  assign new_G1014gat_ = G154gat & G494gat;
  assign new_G1017gat_ = G154gat & G511gat;
  assign new_G1020gat_ = G154gat & G528gat;
  assign new_G1023gat_ = G171gat & G273gat;
  assign new_G1026gat_ = G171gat & G290gat;
  assign new_G1029gat_ = G171gat & G307gat;
  assign new_G1032gat_ = G171gat & G324gat;
  assign new_G1035gat_ = G171gat & G341gat;
  assign new_G1038gat_ = G171gat & G358gat;
  assign new_G1041gat_ = G171gat & G375gat;
  assign new_G1044gat_ = G171gat & G392gat;
  assign new_G1047gat_ = G171gat & G409gat;
  assign new_G1050gat_ = G171gat & G426gat;
  assign new_G1053gat_ = G171gat & G443gat;
  assign new_G1056gat_ = G171gat & G460gat;
  assign new_G1059gat_ = G171gat & G477gat;
  assign new_G1062gat_ = G171gat & G494gat;
  assign new_G1065gat_ = G171gat & G511gat;
  assign new_G1068gat_ = G171gat & G528gat;
  assign new_G1071gat_ = G188gat & G273gat;
  assign new_G1074gat_ = G188gat & G290gat;
  assign new_G1077gat_ = G188gat & G307gat;
  assign new_G1080gat_ = G188gat & G324gat;
  assign new_G1083gat_ = G188gat & G341gat;
  assign new_G1086gat_ = G188gat & G358gat;
  assign new_G1089gat_ = G188gat & G375gat;
  assign new_G1092gat_ = G188gat & G392gat;
  assign new_G1095gat_ = G188gat & G409gat;
  assign new_G1098gat_ = G188gat & G426gat;
  assign new_G1101gat_ = G188gat & G443gat;
  assign new_G1104gat_ = G188gat & G460gat;
  assign new_G1107gat_ = G188gat & G477gat;
  assign new_G1110gat_ = G188gat & G494gat;
  assign new_G1113gat_ = G188gat & G511gat;
  assign new_G1116gat_ = G188gat & G528gat;
  assign new_G1119gat_ = G205gat & G273gat;
  assign new_G1122gat_ = G205gat & G290gat;
  assign new_G1125gat_ = G205gat & G307gat;
  assign new_G1128gat_ = G205gat & G324gat;
  assign new_G1131gat_ = G205gat & G341gat;
  assign new_G1134gat_ = G205gat & G358gat;
  assign new_G1137gat_ = G205gat & G375gat;
  assign new_G1140gat_ = G205gat & G392gat;
  assign new_G1143gat_ = G205gat & G409gat;
  assign new_G1146gat_ = G205gat & G426gat;
  assign new_G1149gat_ = G205gat & G443gat;
  assign new_G1152gat_ = G205gat & G460gat;
  assign new_G1155gat_ = G205gat & G477gat;
  assign new_G1158gat_ = G205gat & G494gat;
  assign new_G1161gat_ = G205gat & G511gat;
  assign new_G1164gat_ = G205gat & G528gat;
  assign new_G1167gat_ = G222gat & G273gat;
  assign new_G1170gat_ = G222gat & G290gat;
  assign new_G1173gat_ = G222gat & G307gat;
  assign new_G1176gat_ = G222gat & G324gat;
  assign new_G1179gat_ = G222gat & G341gat;
  assign new_G1182gat_ = G222gat & G358gat;
  assign new_G1185gat_ = G222gat & G375gat;
  assign new_G1188gat_ = G222gat & G392gat;
  assign new_G1191gat_ = G222gat & G409gat;
  assign new_G1194gat_ = G222gat & G426gat;
  assign new_G1197gat_ = G222gat & G443gat;
  assign new_G1200gat_ = G222gat & G460gat;
  assign new_G1203gat_ = G222gat & G477gat;
  assign new_G1206gat_ = G222gat & G494gat;
  assign new_G1209gat_ = G222gat & G511gat;
  assign new_G1212gat_ = G222gat & G528gat;
  assign new_G1215gat_ = G239gat & G273gat;
  assign new_G1218gat_ = G239gat & G290gat;
  assign new_G1221gat_ = G239gat & G307gat;
  assign new_G1224gat_ = G239gat & G324gat;
  assign new_G1227gat_ = G239gat & G341gat;
  assign new_G1230gat_ = G239gat & G358gat;
  assign new_G1233gat_ = G239gat & G375gat;
  assign new_G1236gat_ = G239gat & G392gat;
  assign new_G1239gat_ = G239gat & G409gat;
  assign new_G1242gat_ = G239gat & G426gat;
  assign new_G1245gat_ = G239gat & G443gat;
  assign new_G1248gat_ = G239gat & G460gat;
  assign new_G1251gat_ = G239gat & G477gat;
  assign new_G1254gat_ = G239gat & G494gat;
  assign new_G1257gat_ = G239gat & G511gat;
  assign new_G1260gat_ = G239gat & G528gat;
  assign new_G1263gat_ = G256gat & G273gat;
  assign new_G1266gat_ = G256gat & G290gat;
  assign new_G1269gat_ = G256gat & G307gat;
  assign new_G1272gat_ = G256gat & G324gat;
  assign new_G1275gat_ = G256gat & G341gat;
  assign new_G1278gat_ = G256gat & G358gat;
  assign new_G1281gat_ = G256gat & G375gat;
  assign new_G1284gat_ = G256gat & G392gat;
  assign new_G1287gat_ = G256gat & G409gat;
  assign new_G1290gat_ = G256gat & G426gat;
  assign new_G1293gat_ = G256gat & G443gat;
  assign new_G1296gat_ = G256gat & G460gat;
  assign new_G1299gat_ = G256gat & G477gat;
  assign new_G1302gat_ = G256gat & G494gat;
  assign new_G1305gat_ = G256gat & G511gat;
  assign new_G1308gat_ = G256gat & G528gat;
  assign new_G1311gat_ = ~new_G591gat_;
  assign new_G1315gat_ = ~new_G639gat_;
  assign new_G1319gat_ = ~new_G687gat_;
  assign new_G1323gat_ = ~new_G735gat_;
  assign new_G1327gat_ = ~new_G783gat_;
  assign new_G1331gat_ = ~new_G831gat_;
  assign new_G1335gat_ = ~new_G879gat_;
  assign new_G1339gat_ = ~new_G927gat_;
  assign new_G1343gat_ = ~new_G975gat_;
  assign new_G1347gat_ = ~new_G1023gat_;
  assign new_G1351gat_ = ~new_G1071gat_;
  assign new_G1355gat_ = ~new_G1119gat_;
  assign new_G1359gat_ = ~new_G1167gat_;
  assign new_G1363gat_ = ~new_G1215gat_;
  assign new_G1367gat_ = ~new_G1263gat_;
  assign new_G1371gat_ = ~new_G591gat_ & ~new_G1311gat_;
  assign new_G1372gat_ = ~new_G1311gat_;
  assign new_G1373gat_ = ~new_G639gat_ & ~new_G1315gat_;
  assign new_G1374gat_ = ~new_G1315gat_;
  assign new_G1375gat_ = ~new_G687gat_ & ~new_G1319gat_;
  assign new_G1376gat_ = ~new_G1319gat_;
  assign new_G1377gat_ = ~new_G735gat_ & ~new_G1323gat_;
  assign new_G1378gat_ = ~new_G1323gat_;
  assign new_G1379gat_ = ~new_G783gat_ & ~new_G1327gat_;
  assign new_G1380gat_ = ~new_G1327gat_;
  assign new_G1381gat_ = ~new_G831gat_ & ~new_G1331gat_;
  assign new_G1382gat_ = ~new_G1331gat_;
  assign new_G1383gat_ = ~new_G879gat_ & ~new_G1335gat_;
  assign new_G1384gat_ = ~new_G1335gat_;
  assign new_G1385gat_ = ~new_G927gat_ & ~new_G1339gat_;
  assign new_G1386gat_ = ~new_G1339gat_;
  assign new_G1387gat_ = ~new_G975gat_ & ~new_G1343gat_;
  assign new_G1388gat_ = ~new_G1343gat_;
  assign new_G1389gat_ = ~new_G1023gat_ & ~new_G1347gat_;
  assign new_G1390gat_ = ~new_G1347gat_;
  assign new_G1391gat_ = ~new_G1071gat_ & ~new_G1351gat_;
  assign new_G1392gat_ = ~new_G1351gat_;
  assign new_G1393gat_ = ~new_G1119gat_ & ~new_G1355gat_;
  assign new_G1394gat_ = ~new_G1355gat_;
  assign new_G1395gat_ = ~new_G1167gat_ & ~new_G1359gat_;
  assign new_G1396gat_ = ~new_G1359gat_;
  assign new_G1397gat_ = ~new_G1215gat_ & ~new_G1363gat_;
  assign new_G1398gat_ = ~new_G1363gat_;
  assign new_G1399gat_ = ~new_G1263gat_ & ~new_G1367gat_;
  assign new_G1400gat_ = ~new_G1367gat_;
  assign new_G1401gat_ = ~new_G1371gat_ & ~new_G1372gat_;
  assign new_G1404gat_ = ~new_G1373gat_ & ~new_G1374gat_;
  assign new_G1407gat_ = ~new_G1375gat_ & ~new_G1376gat_;
  assign new_G1410gat_ = ~new_G1377gat_ & ~new_G1378gat_;
  assign new_G1413gat_ = ~new_G1379gat_ & ~new_G1380gat_;
  assign new_G1416gat_ = ~new_G1381gat_ & ~new_G1382gat_;
  assign new_G1419gat_ = ~new_G1383gat_ & ~new_G1384gat_;
  assign new_G1422gat_ = ~new_G1385gat_ & ~new_G1386gat_;
  assign new_G1425gat_ = ~new_G1387gat_ & ~new_G1388gat_;
  assign new_G1428gat_ = ~new_G1389gat_ & ~new_G1390gat_;
  assign new_G1431gat_ = ~new_G1391gat_ & ~new_G1392gat_;
  assign new_G1434gat_ = ~new_G1393gat_ & ~new_G1394gat_;
  assign new_G1437gat_ = ~new_G1395gat_ & ~new_G1396gat_;
  assign new_G1440gat_ = ~new_G1397gat_ & ~new_G1398gat_;
  assign new_G1443gat_ = ~new_G1399gat_ & ~new_G1400gat_;
  assign new_G1446gat_ = ~new_G1401gat_ & ~new_G546gat_;
  assign new_G1450gat_ = ~new_G1404gat_ & ~new_G594gat_;
  assign new_G1454gat_ = ~new_G1407gat_ & ~new_G642gat_;
  assign new_G1458gat_ = ~new_G1410gat_ & ~new_G690gat_;
  assign new_G1462gat_ = ~new_G1413gat_ & ~new_G738gat_;
  assign new_G1466gat_ = ~new_G1416gat_ & ~new_G786gat_;
  assign new_G1470gat_ = ~new_G1419gat_ & ~new_G834gat_;
  assign new_G1474gat_ = ~new_G1422gat_ & ~new_G882gat_;
  assign new_G1478gat_ = ~new_G1425gat_ & ~new_G930gat_;
  assign new_G1482gat_ = ~new_G1428gat_ & ~new_G978gat_;
  assign new_G1486gat_ = ~new_G1431gat_ & ~new_G1026gat_;
  assign new_G1490gat_ = ~new_G1434gat_ & ~new_G1074gat_;
  assign new_G1494gat_ = ~new_G1437gat_ & ~new_G1122gat_;
  assign new_G1498gat_ = ~new_G1440gat_ & ~new_G1170gat_;
  assign new_G1502gat_ = ~new_G1443gat_ & ~new_G1218gat_;
  assign new_G1506gat_ = ~new_G1401gat_ & ~new_G1446gat_;
  assign new_G1507gat_ = ~new_G1446gat_ & ~new_G546gat_;
  assign new_G1508gat_ = ~new_G1311gat_ & ~new_G1446gat_;
  assign new_G1511gat_ = ~new_G1404gat_ & ~new_G1450gat_;
  assign new_G1512gat_ = ~new_G1450gat_ & ~new_G594gat_;
  assign new_G1513gat_ = ~new_G1315gat_ & ~new_G1450gat_;
  assign new_G1516gat_ = ~new_G1407gat_ & ~new_G1454gat_;
  assign new_G1517gat_ = ~new_G1454gat_ & ~new_G642gat_;
  assign new_G1518gat_ = ~new_G1319gat_ & ~new_G1454gat_;
  assign new_G1521gat_ = ~new_G1410gat_ & ~new_G1458gat_;
  assign new_G1522gat_ = ~new_G1458gat_ & ~new_G690gat_;
  assign new_G1523gat_ = ~new_G1323gat_ & ~new_G1458gat_;
  assign new_G1526gat_ = ~new_G1413gat_ & ~new_G1462gat_;
  assign new_G1527gat_ = ~new_G1462gat_ & ~new_G738gat_;
  assign new_G1528gat_ = ~new_G1327gat_ & ~new_G1462gat_;
  assign new_G1531gat_ = ~new_G1416gat_ & ~new_G1466gat_;
  assign new_G1532gat_ = ~new_G1466gat_ & ~new_G786gat_;
  assign new_G1533gat_ = ~new_G1331gat_ & ~new_G1466gat_;
  assign new_G1536gat_ = ~new_G1419gat_ & ~new_G1470gat_;
  assign new_G1537gat_ = ~new_G1470gat_ & ~new_G834gat_;
  assign new_G1538gat_ = ~new_G1335gat_ & ~new_G1470gat_;
  assign new_G1541gat_ = ~new_G1422gat_ & ~new_G1474gat_;
  assign new_G1542gat_ = ~new_G1474gat_ & ~new_G882gat_;
  assign new_G1543gat_ = ~new_G1339gat_ & ~new_G1474gat_;
  assign new_G1546gat_ = ~new_G1425gat_ & ~new_G1478gat_;
  assign new_G1547gat_ = ~new_G1478gat_ & ~new_G930gat_;
  assign new_G1548gat_ = ~new_G1343gat_ & ~new_G1478gat_;
  assign new_G1551gat_ = ~new_G1428gat_ & ~new_G1482gat_;
  assign new_G1552gat_ = ~new_G1482gat_ & ~new_G978gat_;
  assign new_G1553gat_ = ~new_G1347gat_ & ~new_G1482gat_;
  assign new_G1556gat_ = ~new_G1431gat_ & ~new_G1486gat_;
  assign new_G1557gat_ = ~new_G1486gat_ & ~new_G1026gat_;
  assign new_G1558gat_ = ~new_G1351gat_ & ~new_G1486gat_;
  assign new_G1561gat_ = ~new_G1434gat_ & ~new_G1490gat_;
  assign new_G1562gat_ = ~new_G1490gat_ & ~new_G1074gat_;
  assign new_G1563gat_ = ~new_G1355gat_ & ~new_G1490gat_;
  assign new_G1566gat_ = ~new_G1437gat_ & ~new_G1494gat_;
  assign new_G1567gat_ = ~new_G1494gat_ & ~new_G1122gat_;
  assign new_G1568gat_ = ~new_G1359gat_ & ~new_G1494gat_;
  assign new_G1571gat_ = ~new_G1440gat_ & ~new_G1498gat_;
  assign new_G1572gat_ = ~new_G1498gat_ & ~new_G1170gat_;
  assign new_G1573gat_ = ~new_G1363gat_ & ~new_G1498gat_;
  assign new_G1576gat_ = ~new_G1443gat_ & ~new_G1502gat_;
  assign new_G1577gat_ = ~new_G1502gat_ & ~new_G1218gat_;
  assign new_G1578gat_ = ~new_G1367gat_ & ~new_G1502gat_;
  assign G1581gat = ~new_G1506gat_ & ~new_G1507gat_;
  assign new_G1582gat_ = ~new_G1511gat_ & ~new_G1512gat_;
  assign new_G1585gat_ = ~new_G1516gat_ & ~new_G1517gat_;
  assign new_G1588gat_ = ~new_G1521gat_ & ~new_G1522gat_;
  assign new_G1591gat_ = ~new_G1526gat_ & ~new_G1527gat_;
  assign new_G1594gat_ = ~new_G1531gat_ & ~new_G1532gat_;
  assign new_G1597gat_ = ~new_G1536gat_ & ~new_G1537gat_;
  assign new_G1600gat_ = ~new_G1541gat_ & ~new_G1542gat_;
  assign new_G1603gat_ = ~new_G1546gat_ & ~new_G1547gat_;
  assign new_G1606gat_ = ~new_G1551gat_ & ~new_G1552gat_;
  assign new_G1609gat_ = ~new_G1556gat_ & ~new_G1557gat_;
  assign new_G1612gat_ = ~new_G1561gat_ & ~new_G1562gat_;
  assign new_G1615gat_ = ~new_G1566gat_ & ~new_G1567gat_;
  assign new_G1618gat_ = ~new_G1571gat_ & ~new_G1572gat_;
  assign new_G1621gat_ = ~new_G1576gat_ & ~new_G1577gat_;
  assign new_G1624gat_ = ~new_G1266gat_ & ~new_G1578gat_;
  assign new_G1628gat_ = ~new_G1582gat_ & ~new_G1508gat_;
  assign new_G1632gat_ = ~new_G1585gat_ & ~new_G1513gat_;
  assign new_G1636gat_ = ~new_G1588gat_ & ~new_G1518gat_;
  assign new_G1640gat_ = ~new_G1591gat_ & ~new_G1523gat_;
  assign new_G1644gat_ = ~new_G1594gat_ & ~new_G1528gat_;
  assign new_G1648gat_ = ~new_G1597gat_ & ~new_G1533gat_;
  assign new_G1652gat_ = ~new_G1600gat_ & ~new_G1538gat_;
  assign new_G1656gat_ = ~new_G1603gat_ & ~new_G1543gat_;
  assign new_G1660gat_ = ~new_G1606gat_ & ~new_G1548gat_;
  assign new_G1664gat_ = ~new_G1609gat_ & ~new_G1553gat_;
  assign new_G1668gat_ = ~new_G1612gat_ & ~new_G1558gat_;
  assign new_G1672gat_ = ~new_G1615gat_ & ~new_G1563gat_;
  assign new_G1676gat_ = ~new_G1618gat_ & ~new_G1568gat_;
  assign new_G1680gat_ = ~new_G1621gat_ & ~new_G1573gat_;
  assign new_G1684gat_ = ~new_G1266gat_ & ~new_G1624gat_;
  assign new_G1685gat_ = ~new_G1624gat_ & ~new_G1578gat_;
  assign new_G1686gat_ = ~new_G1582gat_ & ~new_G1628gat_;
  assign new_G1687gat_ = ~new_G1628gat_ & ~new_G1508gat_;
  assign new_G1688gat_ = ~new_G1585gat_ & ~new_G1632gat_;
  assign new_G1689gat_ = ~new_G1632gat_ & ~new_G1513gat_;
  assign new_G1690gat_ = ~new_G1588gat_ & ~new_G1636gat_;
  assign new_G1691gat_ = ~new_G1636gat_ & ~new_G1518gat_;
  assign new_G1692gat_ = ~new_G1591gat_ & ~new_G1640gat_;
  assign new_G1693gat_ = ~new_G1640gat_ & ~new_G1523gat_;
  assign new_G1694gat_ = ~new_G1594gat_ & ~new_G1644gat_;
  assign new_G1695gat_ = ~new_G1644gat_ & ~new_G1528gat_;
  assign new_G1696gat_ = ~new_G1597gat_ & ~new_G1648gat_;
  assign new_G1697gat_ = ~new_G1648gat_ & ~new_G1533gat_;
  assign new_G1698gat_ = ~new_G1600gat_ & ~new_G1652gat_;
  assign new_G1699gat_ = ~new_G1652gat_ & ~new_G1538gat_;
  assign new_G1700gat_ = ~new_G1603gat_ & ~new_G1656gat_;
  assign new_G1701gat_ = ~new_G1656gat_ & ~new_G1543gat_;
  assign new_G1702gat_ = ~new_G1606gat_ & ~new_G1660gat_;
  assign new_G1703gat_ = ~new_G1660gat_ & ~new_G1548gat_;
  assign new_G1704gat_ = ~new_G1609gat_ & ~new_G1664gat_;
  assign new_G1705gat_ = ~new_G1664gat_ & ~new_G1553gat_;
  assign new_G1706gat_ = ~new_G1612gat_ & ~new_G1668gat_;
  assign new_G1707gat_ = ~new_G1668gat_ & ~new_G1558gat_;
  assign new_G1708gat_ = ~new_G1615gat_ & ~new_G1672gat_;
  assign new_G1709gat_ = ~new_G1672gat_ & ~new_G1563gat_;
  assign new_G1710gat_ = ~new_G1618gat_ & ~new_G1676gat_;
  assign new_G1711gat_ = ~new_G1676gat_ & ~new_G1568gat_;
  assign new_G1712gat_ = ~new_G1621gat_ & ~new_G1680gat_;
  assign new_G1713gat_ = ~new_G1680gat_ & ~new_G1573gat_;
  assign new_G1714gat_ = ~new_G1684gat_ & ~new_G1685gat_;
  assign new_G1717gat_ = ~new_G1686gat_ & ~new_G1687gat_;
  assign new_G1720gat_ = ~new_G1688gat_ & ~new_G1689gat_;
  assign new_G1723gat_ = ~new_G1690gat_ & ~new_G1691gat_;
  assign new_G1726gat_ = ~new_G1692gat_ & ~new_G1693gat_;
  assign new_G1729gat_ = ~new_G1694gat_ & ~new_G1695gat_;
  assign new_G1732gat_ = ~new_G1696gat_ & ~new_G1697gat_;
  assign new_G1735gat_ = ~new_G1698gat_ & ~new_G1699gat_;
  assign new_G1738gat_ = ~new_G1700gat_ & ~new_G1701gat_;
  assign new_G1741gat_ = ~new_G1702gat_ & ~new_G1703gat_;
  assign new_G1744gat_ = ~new_G1704gat_ & ~new_G1705gat_;
  assign new_G1747gat_ = ~new_G1706gat_ & ~new_G1707gat_;
  assign new_G1750gat_ = ~new_G1708gat_ & ~new_G1709gat_;
  assign new_G1753gat_ = ~new_G1710gat_ & ~new_G1711gat_;
  assign new_G1756gat_ = ~new_G1712gat_ & ~new_G1713gat_;
  assign new_G1759gat_ = ~new_G1714gat_ & ~new_G1221gat_;
  assign new_G1763gat_ = ~new_G1717gat_ & ~new_G549gat_;
  assign new_G1767gat_ = ~new_G1720gat_ & ~new_G597gat_;
  assign new_G1771gat_ = ~new_G1723gat_ & ~new_G645gat_;
  assign new_G1775gat_ = ~new_G1726gat_ & ~new_G693gat_;
  assign new_G1779gat_ = ~new_G1729gat_ & ~new_G741gat_;
  assign new_G1783gat_ = ~new_G1732gat_ & ~new_G789gat_;
  assign new_G1787gat_ = ~new_G1735gat_ & ~new_G837gat_;
  assign new_G1791gat_ = ~new_G1738gat_ & ~new_G885gat_;
  assign new_G1795gat_ = ~new_G1741gat_ & ~new_G933gat_;
  assign new_G1799gat_ = ~new_G1744gat_ & ~new_G981gat_;
  assign new_G1803gat_ = ~new_G1747gat_ & ~new_G1029gat_;
  assign new_G1807gat_ = ~new_G1750gat_ & ~new_G1077gat_;
  assign new_G1811gat_ = ~new_G1753gat_ & ~new_G1125gat_;
  assign new_G1815gat_ = ~new_G1756gat_ & ~new_G1173gat_;
  assign new_G1819gat_ = ~new_G1714gat_ & ~new_G1759gat_;
  assign new_G1820gat_ = ~new_G1759gat_ & ~new_G1221gat_;
  assign new_G1821gat_ = ~new_G1624gat_ & ~new_G1759gat_;
  assign new_G1824gat_ = ~new_G1717gat_ & ~new_G1763gat_;
  assign new_G1825gat_ = ~new_G1763gat_ & ~new_G549gat_;
  assign new_G1826gat_ = ~new_G1628gat_ & ~new_G1763gat_;
  assign new_G1829gat_ = ~new_G1720gat_ & ~new_G1767gat_;
  assign new_G1830gat_ = ~new_G1767gat_ & ~new_G597gat_;
  assign new_G1831gat_ = ~new_G1632gat_ & ~new_G1767gat_;
  assign new_G1834gat_ = ~new_G1723gat_ & ~new_G1771gat_;
  assign new_G1835gat_ = ~new_G1771gat_ & ~new_G645gat_;
  assign new_G1836gat_ = ~new_G1636gat_ & ~new_G1771gat_;
  assign new_G1839gat_ = ~new_G1726gat_ & ~new_G1775gat_;
  assign new_G1840gat_ = ~new_G1775gat_ & ~new_G693gat_;
  assign new_G1841gat_ = ~new_G1640gat_ & ~new_G1775gat_;
  assign new_G1844gat_ = ~new_G1729gat_ & ~new_G1779gat_;
  assign new_G1845gat_ = ~new_G1779gat_ & ~new_G741gat_;
  assign new_G1846gat_ = ~new_G1644gat_ & ~new_G1779gat_;
  assign new_G1849gat_ = ~new_G1732gat_ & ~new_G1783gat_;
  assign new_G1850gat_ = ~new_G1783gat_ & ~new_G789gat_;
  assign new_G1851gat_ = ~new_G1648gat_ & ~new_G1783gat_;
  assign new_G1854gat_ = ~new_G1735gat_ & ~new_G1787gat_;
  assign new_G1855gat_ = ~new_G1787gat_ & ~new_G837gat_;
  assign new_G1856gat_ = ~new_G1652gat_ & ~new_G1787gat_;
  assign new_G1859gat_ = ~new_G1738gat_ & ~new_G1791gat_;
  assign new_G1860gat_ = ~new_G1791gat_ & ~new_G885gat_;
  assign new_G1861gat_ = ~new_G1656gat_ & ~new_G1791gat_;
  assign new_G1864gat_ = ~new_G1741gat_ & ~new_G1795gat_;
  assign new_G1865gat_ = ~new_G1795gat_ & ~new_G933gat_;
  assign new_G1866gat_ = ~new_G1660gat_ & ~new_G1795gat_;
  assign new_G1869gat_ = ~new_G1744gat_ & ~new_G1799gat_;
  assign new_G1870gat_ = ~new_G1799gat_ & ~new_G981gat_;
  assign new_G1871gat_ = ~new_G1664gat_ & ~new_G1799gat_;
  assign new_G1874gat_ = ~new_G1747gat_ & ~new_G1803gat_;
  assign new_G1875gat_ = ~new_G1803gat_ & ~new_G1029gat_;
  assign new_G1876gat_ = ~new_G1668gat_ & ~new_G1803gat_;
  assign new_G1879gat_ = ~new_G1750gat_ & ~new_G1807gat_;
  assign new_G1880gat_ = ~new_G1807gat_ & ~new_G1077gat_;
  assign new_G1881gat_ = ~new_G1672gat_ & ~new_G1807gat_;
  assign new_G1884gat_ = ~new_G1753gat_ & ~new_G1811gat_;
  assign new_G1885gat_ = ~new_G1811gat_ & ~new_G1125gat_;
  assign new_G1886gat_ = ~new_G1676gat_ & ~new_G1811gat_;
  assign new_G1889gat_ = ~new_G1756gat_ & ~new_G1815gat_;
  assign new_G1890gat_ = ~new_G1815gat_ & ~new_G1173gat_;
  assign new_G1891gat_ = ~new_G1680gat_ & ~new_G1815gat_;
  assign new_G1894gat_ = ~new_G1819gat_ & ~new_G1820gat_;
  assign new_G1897gat_ = ~new_G1269gat_ & ~new_G1821gat_;
  assign G1901gat = ~new_G1824gat_ & ~new_G1825gat_;
  assign new_G1902gat_ = ~new_G1829gat_ & ~new_G1830gat_;
  assign new_G1905gat_ = ~new_G1834gat_ & ~new_G1835gat_;
  assign new_G1908gat_ = ~new_G1839gat_ & ~new_G1840gat_;
  assign new_G1911gat_ = ~new_G1844gat_ & ~new_G1845gat_;
  assign new_G1914gat_ = ~new_G1849gat_ & ~new_G1850gat_;
  assign new_G1917gat_ = ~new_G1854gat_ & ~new_G1855gat_;
  assign new_G1920gat_ = ~new_G1859gat_ & ~new_G1860gat_;
  assign new_G1923gat_ = ~new_G1864gat_ & ~new_G1865gat_;
  assign new_G1926gat_ = ~new_G1869gat_ & ~new_G1870gat_;
  assign new_G1929gat_ = ~new_G1874gat_ & ~new_G1875gat_;
  assign new_G1932gat_ = ~new_G1879gat_ & ~new_G1880gat_;
  assign new_G1935gat_ = ~new_G1884gat_ & ~new_G1885gat_;
  assign new_G1938gat_ = ~new_G1889gat_ & ~new_G1890gat_;
  assign new_G1941gat_ = ~new_G1894gat_ & ~new_G1891gat_;
  assign new_G1945gat_ = ~new_G1269gat_ & ~new_G1897gat_;
  assign new_G1946gat_ = ~new_G1897gat_ & ~new_G1821gat_;
  assign new_G1947gat_ = ~new_G1902gat_ & ~new_G1826gat_;
  assign new_G1951gat_ = ~new_G1905gat_ & ~new_G1831gat_;
  assign new_G1955gat_ = ~new_G1908gat_ & ~new_G1836gat_;
  assign new_G1959gat_ = ~new_G1911gat_ & ~new_G1841gat_;
  assign new_G1963gat_ = ~new_G1914gat_ & ~new_G1846gat_;
  assign new_G1967gat_ = ~new_G1917gat_ & ~new_G1851gat_;
  assign new_G1971gat_ = ~new_G1920gat_ & ~new_G1856gat_;
  assign new_G1975gat_ = ~new_G1923gat_ & ~new_G1861gat_;
  assign new_G1979gat_ = ~new_G1926gat_ & ~new_G1866gat_;
  assign new_G1983gat_ = ~new_G1929gat_ & ~new_G1871gat_;
  assign new_G1987gat_ = ~new_G1932gat_ & ~new_G1876gat_;
  assign new_G1991gat_ = ~new_G1935gat_ & ~new_G1881gat_;
  assign new_G1995gat_ = ~new_G1938gat_ & ~new_G1886gat_;
  assign new_G1999gat_ = ~new_G1894gat_ & ~new_G1941gat_;
  assign new_G2000gat_ = ~new_G1941gat_ & ~new_G1891gat_;
  assign new_G2001gat_ = ~new_G1945gat_ & ~new_G1946gat_;
  assign new_G2004gat_ = ~new_G1902gat_ & ~new_G1947gat_;
  assign new_G2005gat_ = ~new_G1947gat_ & ~new_G1826gat_;
  assign new_G2006gat_ = ~new_G1905gat_ & ~new_G1951gat_;
  assign new_G2007gat_ = ~new_G1951gat_ & ~new_G1831gat_;
  assign new_G2008gat_ = ~new_G1908gat_ & ~new_G1955gat_;
  assign new_G2009gat_ = ~new_G1955gat_ & ~new_G1836gat_;
  assign new_G2010gat_ = ~new_G1911gat_ & ~new_G1959gat_;
  assign new_G2011gat_ = ~new_G1959gat_ & ~new_G1841gat_;
  assign new_G2012gat_ = ~new_G1914gat_ & ~new_G1963gat_;
  assign new_G2013gat_ = ~new_G1963gat_ & ~new_G1846gat_;
  assign new_G2014gat_ = ~new_G1917gat_ & ~new_G1967gat_;
  assign new_G2015gat_ = ~new_G1967gat_ & ~new_G1851gat_;
  assign new_G2016gat_ = ~new_G1920gat_ & ~new_G1971gat_;
  assign new_G2017gat_ = ~new_G1971gat_ & ~new_G1856gat_;
  assign new_G2018gat_ = ~new_G1923gat_ & ~new_G1975gat_;
  assign new_G2019gat_ = ~new_G1975gat_ & ~new_G1861gat_;
  assign new_G2020gat_ = ~new_G1926gat_ & ~new_G1979gat_;
  assign new_G2021gat_ = ~new_G1979gat_ & ~new_G1866gat_;
  assign new_G2022gat_ = ~new_G1929gat_ & ~new_G1983gat_;
  assign new_G2023gat_ = ~new_G1983gat_ & ~new_G1871gat_;
  assign new_G2024gat_ = ~new_G1932gat_ & ~new_G1987gat_;
  assign new_G2025gat_ = ~new_G1987gat_ & ~new_G1876gat_;
  assign new_G2026gat_ = ~new_G1935gat_ & ~new_G1991gat_;
  assign new_G2027gat_ = ~new_G1991gat_ & ~new_G1881gat_;
  assign new_G2028gat_ = ~new_G1938gat_ & ~new_G1995gat_;
  assign new_G2029gat_ = ~new_G1995gat_ & ~new_G1886gat_;
  assign new_G2030gat_ = ~new_G1999gat_ & ~new_G2000gat_;
  assign new_G2033gat_ = ~new_G2001gat_ & ~new_G1224gat_;
  assign new_G2037gat_ = ~new_G2004gat_ & ~new_G2005gat_;
  assign new_G2040gat_ = ~new_G2006gat_ & ~new_G2007gat_;
  assign new_G2043gat_ = ~new_G2008gat_ & ~new_G2009gat_;
  assign new_G2046gat_ = ~new_G2010gat_ & ~new_G2011gat_;
  assign new_G2049gat_ = ~new_G2012gat_ & ~new_G2013gat_;
  assign new_G2052gat_ = ~new_G2014gat_ & ~new_G2015gat_;
  assign new_G2055gat_ = ~new_G2016gat_ & ~new_G2017gat_;
  assign new_G2058gat_ = ~new_G2018gat_ & ~new_G2019gat_;
  assign new_G2061gat_ = ~new_G2020gat_ & ~new_G2021gat_;
  assign new_G2064gat_ = ~new_G2022gat_ & ~new_G2023gat_;
  assign new_G2067gat_ = ~new_G2024gat_ & ~new_G2025gat_;
  assign new_G2070gat_ = ~new_G2026gat_ & ~new_G2027gat_;
  assign new_G2073gat_ = ~new_G2028gat_ & ~new_G2029gat_;
  assign new_G2076gat_ = ~new_G2030gat_ & ~new_G1176gat_;
  assign new_G2080gat_ = ~new_G2001gat_ & ~new_G2033gat_;
  assign new_G2081gat_ = ~new_G2033gat_ & ~new_G1224gat_;
  assign new_G2082gat_ = ~new_G1897gat_ & ~new_G2033gat_;
  assign new_G2085gat_ = ~new_G2037gat_ & ~new_G552gat_;
  assign new_G2089gat_ = ~new_G2040gat_ & ~new_G600gat_;
  assign new_G2093gat_ = ~new_G2043gat_ & ~new_G648gat_;
  assign new_G2097gat_ = ~new_G2046gat_ & ~new_G696gat_;
  assign new_G2101gat_ = ~new_G2049gat_ & ~new_G744gat_;
  assign new_G2105gat_ = ~new_G2052gat_ & ~new_G792gat_;
  assign new_G2109gat_ = ~new_G2055gat_ & ~new_G840gat_;
  assign new_G2113gat_ = ~new_G2058gat_ & ~new_G888gat_;
  assign new_G2117gat_ = ~new_G2061gat_ & ~new_G936gat_;
  assign new_G2121gat_ = ~new_G2064gat_ & ~new_G984gat_;
  assign new_G2125gat_ = ~new_G2067gat_ & ~new_G1032gat_;
  assign new_G2129gat_ = ~new_G2070gat_ & ~new_G1080gat_;
  assign new_G2133gat_ = ~new_G2073gat_ & ~new_G1128gat_;
  assign new_G2137gat_ = ~new_G2030gat_ & ~new_G2076gat_;
  assign new_G2138gat_ = ~new_G2076gat_ & ~new_G1176gat_;
  assign new_G2139gat_ = ~new_G1941gat_ & ~new_G2076gat_;
  assign new_G2142gat_ = ~new_G2080gat_ & ~new_G2081gat_;
  assign new_G2145gat_ = ~new_G1272gat_ & ~new_G2082gat_;
  assign new_G2149gat_ = ~new_G2037gat_ & ~new_G2085gat_;
  assign new_G2150gat_ = ~new_G2085gat_ & ~new_G552gat_;
  assign new_G2151gat_ = ~new_G1947gat_ & ~new_G2085gat_;
  assign new_G2154gat_ = ~new_G2040gat_ & ~new_G2089gat_;
  assign new_G2155gat_ = ~new_G2089gat_ & ~new_G600gat_;
  assign new_G2156gat_ = ~new_G1951gat_ & ~new_G2089gat_;
  assign new_G2159gat_ = ~new_G2043gat_ & ~new_G2093gat_;
  assign new_G2160gat_ = ~new_G2093gat_ & ~new_G648gat_;
  assign new_G2161gat_ = ~new_G1955gat_ & ~new_G2093gat_;
  assign new_G2164gat_ = ~new_G2046gat_ & ~new_G2097gat_;
  assign new_G2165gat_ = ~new_G2097gat_ & ~new_G696gat_;
  assign new_G2166gat_ = ~new_G1959gat_ & ~new_G2097gat_;
  assign new_G2169gat_ = ~new_G2049gat_ & ~new_G2101gat_;
  assign new_G2170gat_ = ~new_G2101gat_ & ~new_G744gat_;
  assign new_G2171gat_ = ~new_G1963gat_ & ~new_G2101gat_;
  assign new_G2174gat_ = ~new_G2052gat_ & ~new_G2105gat_;
  assign new_G2175gat_ = ~new_G2105gat_ & ~new_G792gat_;
  assign new_G2176gat_ = ~new_G1967gat_ & ~new_G2105gat_;
  assign new_G2179gat_ = ~new_G2055gat_ & ~new_G2109gat_;
  assign new_G2180gat_ = ~new_G2109gat_ & ~new_G840gat_;
  assign new_G2181gat_ = ~new_G1971gat_ & ~new_G2109gat_;
  assign new_G2184gat_ = ~new_G2058gat_ & ~new_G2113gat_;
  assign new_G2185gat_ = ~new_G2113gat_ & ~new_G888gat_;
  assign new_G2186gat_ = ~new_G1975gat_ & ~new_G2113gat_;
  assign new_G2189gat_ = ~new_G2061gat_ & ~new_G2117gat_;
  assign new_G2190gat_ = ~new_G2117gat_ & ~new_G936gat_;
  assign new_G2191gat_ = ~new_G1979gat_ & ~new_G2117gat_;
  assign new_G2194gat_ = ~new_G2064gat_ & ~new_G2121gat_;
  assign new_G2195gat_ = ~new_G2121gat_ & ~new_G984gat_;
  assign new_G2196gat_ = ~new_G1983gat_ & ~new_G2121gat_;
  assign new_G2199gat_ = ~new_G2067gat_ & ~new_G2125gat_;
  assign new_G2200gat_ = ~new_G2125gat_ & ~new_G1032gat_;
  assign new_G2201gat_ = ~new_G1987gat_ & ~new_G2125gat_;
  assign new_G2204gat_ = ~new_G2070gat_ & ~new_G2129gat_;
  assign new_G2205gat_ = ~new_G2129gat_ & ~new_G1080gat_;
  assign new_G2206gat_ = ~new_G1991gat_ & ~new_G2129gat_;
  assign new_G2209gat_ = ~new_G2073gat_ & ~new_G2133gat_;
  assign new_G2210gat_ = ~new_G2133gat_ & ~new_G1128gat_;
  assign new_G2211gat_ = ~new_G1995gat_ & ~new_G2133gat_;
  assign new_G2214gat_ = ~new_G2137gat_ & ~new_G2138gat_;
  assign new_G2217gat_ = ~new_G2142gat_ & ~new_G2139gat_;
  assign new_G2221gat_ = ~new_G1272gat_ & ~new_G2145gat_;
  assign new_G2222gat_ = ~new_G2145gat_ & ~new_G2082gat_;
  assign G2223gat = ~new_G2149gat_ & ~new_G2150gat_;
  assign new_G2224gat_ = ~new_G2154gat_ & ~new_G2155gat_;
  assign new_G2227gat_ = ~new_G2159gat_ & ~new_G2160gat_;
  assign new_G2230gat_ = ~new_G2164gat_ & ~new_G2165gat_;
  assign new_G2233gat_ = ~new_G2169gat_ & ~new_G2170gat_;
  assign new_G2236gat_ = ~new_G2174gat_ & ~new_G2175gat_;
  assign new_G2239gat_ = ~new_G2179gat_ & ~new_G2180gat_;
  assign new_G2242gat_ = ~new_G2184gat_ & ~new_G2185gat_;
  assign new_G2245gat_ = ~new_G2189gat_ & ~new_G2190gat_;
  assign new_G2248gat_ = ~new_G2194gat_ & ~new_G2195gat_;
  assign new_G2251gat_ = ~new_G2199gat_ & ~new_G2200gat_;
  assign new_G2254gat_ = ~new_G2204gat_ & ~new_G2205gat_;
  assign new_G2257gat_ = ~new_G2209gat_ & ~new_G2210gat_;
  assign new_G2260gat_ = ~new_G2214gat_ & ~new_G2211gat_;
  assign new_G2264gat_ = ~new_G2142gat_ & ~new_G2217gat_;
  assign new_G2265gat_ = ~new_G2217gat_ & ~new_G2139gat_;
  assign new_G2266gat_ = ~new_G2221gat_ & ~new_G2222gat_;
  assign new_G2269gat_ = ~new_G2224gat_ & ~new_G2151gat_;
  assign new_G2273gat_ = ~new_G2227gat_ & ~new_G2156gat_;
  assign new_G2277gat_ = ~new_G2230gat_ & ~new_G2161gat_;
  assign new_G2281gat_ = ~new_G2233gat_ & ~new_G2166gat_;
  assign new_G2285gat_ = ~new_G2236gat_ & ~new_G2171gat_;
  assign new_G2289gat_ = ~new_G2239gat_ & ~new_G2176gat_;
  assign new_G2293gat_ = ~new_G2242gat_ & ~new_G2181gat_;
  assign new_G2297gat_ = ~new_G2245gat_ & ~new_G2186gat_;
  assign new_G2301gat_ = ~new_G2248gat_ & ~new_G2191gat_;
  assign new_G2305gat_ = ~new_G2251gat_ & ~new_G2196gat_;
  assign new_G2309gat_ = ~new_G2254gat_ & ~new_G2201gat_;
  assign new_G2313gat_ = ~new_G2257gat_ & ~new_G2206gat_;
  assign new_G2317gat_ = ~new_G2214gat_ & ~new_G2260gat_;
  assign new_G2318gat_ = ~new_G2260gat_ & ~new_G2211gat_;
  assign new_G2319gat_ = ~new_G2264gat_ & ~new_G2265gat_;
  assign new_G2322gat_ = ~new_G2266gat_ & ~new_G1227gat_;
  assign new_G2326gat_ = ~new_G2224gat_ & ~new_G2269gat_;
  assign new_G2327gat_ = ~new_G2269gat_ & ~new_G2151gat_;
  assign new_G2328gat_ = ~new_G2227gat_ & ~new_G2273gat_;
  assign new_G2329gat_ = ~new_G2273gat_ & ~new_G2156gat_;
  assign new_G2330gat_ = ~new_G2230gat_ & ~new_G2277gat_;
  assign new_G2331gat_ = ~new_G2277gat_ & ~new_G2161gat_;
  assign new_G2332gat_ = ~new_G2233gat_ & ~new_G2281gat_;
  assign new_G2333gat_ = ~new_G2281gat_ & ~new_G2166gat_;
  assign new_G2334gat_ = ~new_G2236gat_ & ~new_G2285gat_;
  assign new_G2335gat_ = ~new_G2285gat_ & ~new_G2171gat_;
  assign new_G2336gat_ = ~new_G2239gat_ & ~new_G2289gat_;
  assign new_G2337gat_ = ~new_G2289gat_ & ~new_G2176gat_;
  assign new_G2338gat_ = ~new_G2242gat_ & ~new_G2293gat_;
  assign new_G2339gat_ = ~new_G2293gat_ & ~new_G2181gat_;
  assign new_G2340gat_ = ~new_G2245gat_ & ~new_G2297gat_;
  assign new_G2341gat_ = ~new_G2297gat_ & ~new_G2186gat_;
  assign new_G2342gat_ = ~new_G2248gat_ & ~new_G2301gat_;
  assign new_G2343gat_ = ~new_G2301gat_ & ~new_G2191gat_;
  assign new_G2344gat_ = ~new_G2251gat_ & ~new_G2305gat_;
  assign new_G2345gat_ = ~new_G2305gat_ & ~new_G2196gat_;
  assign new_G2346gat_ = ~new_G2254gat_ & ~new_G2309gat_;
  assign new_G2347gat_ = ~new_G2309gat_ & ~new_G2201gat_;
  assign new_G2348gat_ = ~new_G2257gat_ & ~new_G2313gat_;
  assign new_G2349gat_ = ~new_G2313gat_ & ~new_G2206gat_;
  assign new_G2350gat_ = ~new_G2317gat_ & ~new_G2318gat_;
  assign new_G2353gat_ = ~new_G2319gat_ & ~new_G1179gat_;
  assign new_G2357gat_ = ~new_G2266gat_ & ~new_G2322gat_;
  assign new_G2358gat_ = ~new_G2322gat_ & ~new_G1227gat_;
  assign new_G2359gat_ = ~new_G2145gat_ & ~new_G2322gat_;
  assign new_G2362gat_ = ~new_G2326gat_ & ~new_G2327gat_;
  assign new_G2365gat_ = ~new_G2328gat_ & ~new_G2329gat_;
  assign new_G2368gat_ = ~new_G2330gat_ & ~new_G2331gat_;
  assign new_G2371gat_ = ~new_G2332gat_ & ~new_G2333gat_;
  assign new_G2374gat_ = ~new_G2334gat_ & ~new_G2335gat_;
  assign new_G2377gat_ = ~new_G2336gat_ & ~new_G2337gat_;
  assign new_G2380gat_ = ~new_G2338gat_ & ~new_G2339gat_;
  assign new_G2383gat_ = ~new_G2340gat_ & ~new_G2341gat_;
  assign new_G2386gat_ = ~new_G2342gat_ & ~new_G2343gat_;
  assign new_G2389gat_ = ~new_G2344gat_ & ~new_G2345gat_;
  assign new_G2392gat_ = ~new_G2346gat_ & ~new_G2347gat_;
  assign new_G2395gat_ = ~new_G2348gat_ & ~new_G2349gat_;
  assign new_G2398gat_ = ~new_G2350gat_ & ~new_G1131gat_;
  assign new_G2402gat_ = ~new_G2319gat_ & ~new_G2353gat_;
  assign new_G2403gat_ = ~new_G2353gat_ & ~new_G1179gat_;
  assign new_G2404gat_ = ~new_G2217gat_ & ~new_G2353gat_;
  assign new_G2407gat_ = ~new_G2357gat_ & ~new_G2358gat_;
  assign new_G2410gat_ = ~new_G1275gat_ & ~new_G2359gat_;
  assign new_G2414gat_ = ~new_G2362gat_ & ~new_G555gat_;
  assign new_G2418gat_ = ~new_G2365gat_ & ~new_G603gat_;
  assign new_G2422gat_ = ~new_G2368gat_ & ~new_G651gat_;
  assign new_G2426gat_ = ~new_G2371gat_ & ~new_G699gat_;
  assign new_G2430gat_ = ~new_G2374gat_ & ~new_G747gat_;
  assign new_G2434gat_ = ~new_G2377gat_ & ~new_G795gat_;
  assign new_G2438gat_ = ~new_G2380gat_ & ~new_G843gat_;
  assign new_G2442gat_ = ~new_G2383gat_ & ~new_G891gat_;
  assign new_G2446gat_ = ~new_G2386gat_ & ~new_G939gat_;
  assign new_G2450gat_ = ~new_G2389gat_ & ~new_G987gat_;
  assign new_G2454gat_ = ~new_G2392gat_ & ~new_G1035gat_;
  assign new_G2458gat_ = ~new_G2395gat_ & ~new_G1083gat_;
  assign new_G2462gat_ = ~new_G2350gat_ & ~new_G2398gat_;
  assign new_G2463gat_ = ~new_G2398gat_ & ~new_G1131gat_;
  assign new_G2464gat_ = ~new_G2260gat_ & ~new_G2398gat_;
  assign new_G2467gat_ = ~new_G2402gat_ & ~new_G2403gat_;
  assign new_G2470gat_ = ~new_G2407gat_ & ~new_G2404gat_;
  assign new_G2474gat_ = ~new_G1275gat_ & ~new_G2410gat_;
  assign new_G2475gat_ = ~new_G2410gat_ & ~new_G2359gat_;
  assign new_G2476gat_ = ~new_G2362gat_ & ~new_G2414gat_;
  assign new_G2477gat_ = ~new_G2414gat_ & ~new_G555gat_;
  assign new_G2478gat_ = ~new_G2269gat_ & ~new_G2414gat_;
  assign new_G2481gat_ = ~new_G2365gat_ & ~new_G2418gat_;
  assign new_G2482gat_ = ~new_G2418gat_ & ~new_G603gat_;
  assign new_G2483gat_ = ~new_G2273gat_ & ~new_G2418gat_;
  assign new_G2486gat_ = ~new_G2368gat_ & ~new_G2422gat_;
  assign new_G2487gat_ = ~new_G2422gat_ & ~new_G651gat_;
  assign new_G2488gat_ = ~new_G2277gat_ & ~new_G2422gat_;
  assign new_G2491gat_ = ~new_G2371gat_ & ~new_G2426gat_;
  assign new_G2492gat_ = ~new_G2426gat_ & ~new_G699gat_;
  assign new_G2493gat_ = ~new_G2281gat_ & ~new_G2426gat_;
  assign new_G2496gat_ = ~new_G2374gat_ & ~new_G2430gat_;
  assign new_G2497gat_ = ~new_G2430gat_ & ~new_G747gat_;
  assign new_G2498gat_ = ~new_G2285gat_ & ~new_G2430gat_;
  assign new_G2501gat_ = ~new_G2377gat_ & ~new_G2434gat_;
  assign new_G2502gat_ = ~new_G2434gat_ & ~new_G795gat_;
  assign new_G2503gat_ = ~new_G2289gat_ & ~new_G2434gat_;
  assign new_G2506gat_ = ~new_G2380gat_ & ~new_G2438gat_;
  assign new_G2507gat_ = ~new_G2438gat_ & ~new_G843gat_;
  assign new_G2508gat_ = ~new_G2293gat_ & ~new_G2438gat_;
  assign new_G2511gat_ = ~new_G2383gat_ & ~new_G2442gat_;
  assign new_G2512gat_ = ~new_G2442gat_ & ~new_G891gat_;
  assign new_G2513gat_ = ~new_G2297gat_ & ~new_G2442gat_;
  assign new_G2516gat_ = ~new_G2386gat_ & ~new_G2446gat_;
  assign new_G2517gat_ = ~new_G2446gat_ & ~new_G939gat_;
  assign new_G2518gat_ = ~new_G2301gat_ & ~new_G2446gat_;
  assign new_G2521gat_ = ~new_G2389gat_ & ~new_G2450gat_;
  assign new_G2522gat_ = ~new_G2450gat_ & ~new_G987gat_;
  assign new_G2523gat_ = ~new_G2305gat_ & ~new_G2450gat_;
  assign new_G2526gat_ = ~new_G2392gat_ & ~new_G2454gat_;
  assign new_G2527gat_ = ~new_G2454gat_ & ~new_G1035gat_;
  assign new_G2528gat_ = ~new_G2309gat_ & ~new_G2454gat_;
  assign new_G2531gat_ = ~new_G2395gat_ & ~new_G2458gat_;
  assign new_G2532gat_ = ~new_G2458gat_ & ~new_G1083gat_;
  assign new_G2533gat_ = ~new_G2313gat_ & ~new_G2458gat_;
  assign new_G2536gat_ = ~new_G2462gat_ & ~new_G2463gat_;
  assign new_G2539gat_ = ~new_G2467gat_ & ~new_G2464gat_;
  assign new_G2543gat_ = ~new_G2407gat_ & ~new_G2470gat_;
  assign new_G2544gat_ = ~new_G2470gat_ & ~new_G2404gat_;
  assign new_G2545gat_ = ~new_G2474gat_ & ~new_G2475gat_;
  assign G2548gat = ~new_G2476gat_ & ~new_G2477gat_;
  assign new_G2549gat_ = ~new_G2481gat_ & ~new_G2482gat_;
  assign new_G2552gat_ = ~new_G2486gat_ & ~new_G2487gat_;
  assign new_G2555gat_ = ~new_G2491gat_ & ~new_G2492gat_;
  assign new_G2558gat_ = ~new_G2496gat_ & ~new_G2497gat_;
  assign new_G2561gat_ = ~new_G2501gat_ & ~new_G2502gat_;
  assign new_G2564gat_ = ~new_G2506gat_ & ~new_G2507gat_;
  assign new_G2567gat_ = ~new_G2511gat_ & ~new_G2512gat_;
  assign new_G2570gat_ = ~new_G2516gat_ & ~new_G2517gat_;
  assign new_G2573gat_ = ~new_G2521gat_ & ~new_G2522gat_;
  assign new_G2576gat_ = ~new_G2526gat_ & ~new_G2527gat_;
  assign new_G2579gat_ = ~new_G2531gat_ & ~new_G2532gat_;
  assign new_G2582gat_ = ~new_G2536gat_ & ~new_G2533gat_;
  assign new_G2586gat_ = ~new_G2467gat_ & ~new_G2539gat_;
  assign new_G2587gat_ = ~new_G2539gat_ & ~new_G2464gat_;
  assign new_G2588gat_ = ~new_G2543gat_ & ~new_G2544gat_;
  assign new_G2591gat_ = ~new_G2545gat_ & ~new_G1230gat_;
  assign new_G2595gat_ = ~new_G2549gat_ & ~new_G2478gat_;
  assign new_G2599gat_ = ~new_G2552gat_ & ~new_G2483gat_;
  assign new_G2603gat_ = ~new_G2555gat_ & ~new_G2488gat_;
  assign new_G2607gat_ = ~new_G2558gat_ & ~new_G2493gat_;
  assign new_G2611gat_ = ~new_G2561gat_ & ~new_G2498gat_;
  assign new_G2615gat_ = ~new_G2564gat_ & ~new_G2503gat_;
  assign new_G2619gat_ = ~new_G2567gat_ & ~new_G2508gat_;
  assign new_G2623gat_ = ~new_G2570gat_ & ~new_G2513gat_;
  assign new_G2627gat_ = ~new_G2573gat_ & ~new_G2518gat_;
  assign new_G2631gat_ = ~new_G2576gat_ & ~new_G2523gat_;
  assign new_G2635gat_ = ~new_G2579gat_ & ~new_G2528gat_;
  assign new_G2639gat_ = ~new_G2536gat_ & ~new_G2582gat_;
  assign new_G2640gat_ = ~new_G2582gat_ & ~new_G2533gat_;
  assign new_G2641gat_ = ~new_G2586gat_ & ~new_G2587gat_;
  assign new_G2644gat_ = ~new_G2588gat_ & ~new_G1182gat_;
  assign new_G2648gat_ = ~new_G2545gat_ & ~new_G2591gat_;
  assign new_G2649gat_ = ~new_G2591gat_ & ~new_G1230gat_;
  assign new_G2650gat_ = ~new_G2410gat_ & ~new_G2591gat_;
  assign new_G2653gat_ = ~new_G2549gat_ & ~new_G2595gat_;
  assign new_G2654gat_ = ~new_G2595gat_ & ~new_G2478gat_;
  assign new_G2655gat_ = ~new_G2552gat_ & ~new_G2599gat_;
  assign new_G2656gat_ = ~new_G2599gat_ & ~new_G2483gat_;
  assign new_G2657gat_ = ~new_G2555gat_ & ~new_G2603gat_;
  assign new_G2658gat_ = ~new_G2603gat_ & ~new_G2488gat_;
  assign new_G2659gat_ = ~new_G2558gat_ & ~new_G2607gat_;
  assign new_G2660gat_ = ~new_G2607gat_ & ~new_G2493gat_;
  assign new_G2661gat_ = ~new_G2561gat_ & ~new_G2611gat_;
  assign new_G2662gat_ = ~new_G2611gat_ & ~new_G2498gat_;
  assign new_G2663gat_ = ~new_G2564gat_ & ~new_G2615gat_;
  assign new_G2664gat_ = ~new_G2615gat_ & ~new_G2503gat_;
  assign new_G2665gat_ = ~new_G2567gat_ & ~new_G2619gat_;
  assign new_G2666gat_ = ~new_G2619gat_ & ~new_G2508gat_;
  assign new_G2667gat_ = ~new_G2570gat_ & ~new_G2623gat_;
  assign new_G2668gat_ = ~new_G2623gat_ & ~new_G2513gat_;
  assign new_G2669gat_ = ~new_G2573gat_ & ~new_G2627gat_;
  assign new_G2670gat_ = ~new_G2627gat_ & ~new_G2518gat_;
  assign new_G2671gat_ = ~new_G2576gat_ & ~new_G2631gat_;
  assign new_G2672gat_ = ~new_G2631gat_ & ~new_G2523gat_;
  assign new_G2673gat_ = ~new_G2579gat_ & ~new_G2635gat_;
  assign new_G2674gat_ = ~new_G2635gat_ & ~new_G2528gat_;
  assign new_G2675gat_ = ~new_G2639gat_ & ~new_G2640gat_;
  assign new_G2678gat_ = ~new_G2641gat_ & ~new_G1134gat_;
  assign new_G2682gat_ = ~new_G2588gat_ & ~new_G2644gat_;
  assign new_G2683gat_ = ~new_G2644gat_ & ~new_G1182gat_;
  assign new_G2684gat_ = ~new_G2470gat_ & ~new_G2644gat_;
  assign new_G2687gat_ = ~new_G2648gat_ & ~new_G2649gat_;
  assign new_G2690gat_ = ~new_G1278gat_ & ~new_G2650gat_;
  assign new_G2694gat_ = ~new_G2653gat_ & ~new_G2654gat_;
  assign new_G2697gat_ = ~new_G2655gat_ & ~new_G2656gat_;
  assign new_G2700gat_ = ~new_G2657gat_ & ~new_G2658gat_;
  assign new_G2703gat_ = ~new_G2659gat_ & ~new_G2660gat_;
  assign new_G2706gat_ = ~new_G2661gat_ & ~new_G2662gat_;
  assign new_G2709gat_ = ~new_G2663gat_ & ~new_G2664gat_;
  assign new_G2712gat_ = ~new_G2665gat_ & ~new_G2666gat_;
  assign new_G2715gat_ = ~new_G2667gat_ & ~new_G2668gat_;
  assign new_G2718gat_ = ~new_G2669gat_ & ~new_G2670gat_;
  assign new_G2721gat_ = ~new_G2671gat_ & ~new_G2672gat_;
  assign new_G2724gat_ = ~new_G2673gat_ & ~new_G2674gat_;
  assign new_G2727gat_ = ~new_G2675gat_ & ~new_G1086gat_;
  assign new_G2731gat_ = ~new_G2641gat_ & ~new_G2678gat_;
  assign new_G2732gat_ = ~new_G2678gat_ & ~new_G1134gat_;
  assign new_G2733gat_ = ~new_G2539gat_ & ~new_G2678gat_;
  assign new_G2736gat_ = ~new_G2682gat_ & ~new_G2683gat_;
  assign new_G2739gat_ = ~new_G2687gat_ & ~new_G2684gat_;
  assign new_G2743gat_ = ~new_G1278gat_ & ~new_G2690gat_;
  assign new_G2744gat_ = ~new_G2690gat_ & ~new_G2650gat_;
  assign new_G2745gat_ = ~new_G2694gat_ & ~new_G558gat_;
  assign new_G2749gat_ = ~new_G2697gat_ & ~new_G606gat_;
  assign new_G2753gat_ = ~new_G2700gat_ & ~new_G654gat_;
  assign new_G2757gat_ = ~new_G2703gat_ & ~new_G702gat_;
  assign new_G2761gat_ = ~new_G2706gat_ & ~new_G750gat_;
  assign new_G2765gat_ = ~new_G2709gat_ & ~new_G798gat_;
  assign new_G2769gat_ = ~new_G2712gat_ & ~new_G846gat_;
  assign new_G2773gat_ = ~new_G2715gat_ & ~new_G894gat_;
  assign new_G2777gat_ = ~new_G2718gat_ & ~new_G942gat_;
  assign new_G2781gat_ = ~new_G2721gat_ & ~new_G990gat_;
  assign new_G2785gat_ = ~new_G2724gat_ & ~new_G1038gat_;
  assign new_G2789gat_ = ~new_G2675gat_ & ~new_G2727gat_;
  assign new_G2790gat_ = ~new_G2727gat_ & ~new_G1086gat_;
  assign new_G2791gat_ = ~new_G2582gat_ & ~new_G2727gat_;
  assign new_G2794gat_ = ~new_G2731gat_ & ~new_G2732gat_;
  assign new_G2797gat_ = ~new_G2736gat_ & ~new_G2733gat_;
  assign new_G2801gat_ = ~new_G2687gat_ & ~new_G2739gat_;
  assign new_G2802gat_ = ~new_G2739gat_ & ~new_G2684gat_;
  assign new_G2803gat_ = ~new_G2743gat_ & ~new_G2744gat_;
  assign new_G2806gat_ = ~new_G2694gat_ & ~new_G2745gat_;
  assign new_G2807gat_ = ~new_G2745gat_ & ~new_G558gat_;
  assign new_G2808gat_ = ~new_G2595gat_ & ~new_G2745gat_;
  assign new_G2811gat_ = ~new_G2697gat_ & ~new_G2749gat_;
  assign new_G2812gat_ = ~new_G2749gat_ & ~new_G606gat_;
  assign new_G2813gat_ = ~new_G2599gat_ & ~new_G2749gat_;
  assign new_G2816gat_ = ~new_G2700gat_ & ~new_G2753gat_;
  assign new_G2817gat_ = ~new_G2753gat_ & ~new_G654gat_;
  assign new_G2818gat_ = ~new_G2603gat_ & ~new_G2753gat_;
  assign new_G2821gat_ = ~new_G2703gat_ & ~new_G2757gat_;
  assign new_G2822gat_ = ~new_G2757gat_ & ~new_G702gat_;
  assign new_G2823gat_ = ~new_G2607gat_ & ~new_G2757gat_;
  assign new_G2826gat_ = ~new_G2706gat_ & ~new_G2761gat_;
  assign new_G2827gat_ = ~new_G2761gat_ & ~new_G750gat_;
  assign new_G2828gat_ = ~new_G2611gat_ & ~new_G2761gat_;
  assign new_G2831gat_ = ~new_G2709gat_ & ~new_G2765gat_;
  assign new_G2832gat_ = ~new_G2765gat_ & ~new_G798gat_;
  assign new_G2833gat_ = ~new_G2615gat_ & ~new_G2765gat_;
  assign new_G2836gat_ = ~new_G2712gat_ & ~new_G2769gat_;
  assign new_G2837gat_ = ~new_G2769gat_ & ~new_G846gat_;
  assign new_G2838gat_ = ~new_G2619gat_ & ~new_G2769gat_;
  assign new_G2841gat_ = ~new_G2715gat_ & ~new_G2773gat_;
  assign new_G2842gat_ = ~new_G2773gat_ & ~new_G894gat_;
  assign new_G2843gat_ = ~new_G2623gat_ & ~new_G2773gat_;
  assign new_G2846gat_ = ~new_G2718gat_ & ~new_G2777gat_;
  assign new_G2847gat_ = ~new_G2777gat_ & ~new_G942gat_;
  assign new_G2848gat_ = ~new_G2627gat_ & ~new_G2777gat_;
  assign new_G2851gat_ = ~new_G2721gat_ & ~new_G2781gat_;
  assign new_G2852gat_ = ~new_G2781gat_ & ~new_G990gat_;
  assign new_G2853gat_ = ~new_G2631gat_ & ~new_G2781gat_;
  assign new_G2856gat_ = ~new_G2724gat_ & ~new_G2785gat_;
  assign new_G2857gat_ = ~new_G2785gat_ & ~new_G1038gat_;
  assign new_G2858gat_ = ~new_G2635gat_ & ~new_G2785gat_;
  assign new_G2861gat_ = ~new_G2789gat_ & ~new_G2790gat_;
  assign new_G2864gat_ = ~new_G2794gat_ & ~new_G2791gat_;
  assign new_G2868gat_ = ~new_G2736gat_ & ~new_G2797gat_;
  assign new_G2869gat_ = ~new_G2797gat_ & ~new_G2733gat_;
  assign new_G2870gat_ = ~new_G2801gat_ & ~new_G2802gat_;
  assign new_G2873gat_ = ~new_G2803gat_ & ~new_G1233gat_;
  assign G2877gat = ~new_G2806gat_ & ~new_G2807gat_;
  assign new_G2878gat_ = ~new_G2811gat_ & ~new_G2812gat_;
  assign new_G2881gat_ = ~new_G2816gat_ & ~new_G2817gat_;
  assign new_G2884gat_ = ~new_G2821gat_ & ~new_G2822gat_;
  assign new_G2887gat_ = ~new_G2826gat_ & ~new_G2827gat_;
  assign new_G2890gat_ = ~new_G2831gat_ & ~new_G2832gat_;
  assign new_G2893gat_ = ~new_G2836gat_ & ~new_G2837gat_;
  assign new_G2896gat_ = ~new_G2841gat_ & ~new_G2842gat_;
  assign new_G2899gat_ = ~new_G2846gat_ & ~new_G2847gat_;
  assign new_G2902gat_ = ~new_G2851gat_ & ~new_G2852gat_;
  assign new_G2905gat_ = ~new_G2856gat_ & ~new_G2857gat_;
  assign new_G2908gat_ = ~new_G2861gat_ & ~new_G2858gat_;
  assign new_G2912gat_ = ~new_G2794gat_ & ~new_G2864gat_;
  assign new_G2913gat_ = ~new_G2864gat_ & ~new_G2791gat_;
  assign new_G2914gat_ = ~new_G2868gat_ & ~new_G2869gat_;
  assign new_G2917gat_ = ~new_G2870gat_ & ~new_G1185gat_;
  assign new_G2921gat_ = ~new_G2803gat_ & ~new_G2873gat_;
  assign new_G2922gat_ = ~new_G2873gat_ & ~new_G1233gat_;
  assign new_G2923gat_ = ~new_G2690gat_ & ~new_G2873gat_;
  assign new_G2926gat_ = ~new_G2878gat_ & ~new_G2808gat_;
  assign new_G2930gat_ = ~new_G2881gat_ & ~new_G2813gat_;
  assign new_G2934gat_ = ~new_G2884gat_ & ~new_G2818gat_;
  assign new_G2938gat_ = ~new_G2887gat_ & ~new_G2823gat_;
  assign new_G2942gat_ = ~new_G2890gat_ & ~new_G2828gat_;
  assign new_G2946gat_ = ~new_G2893gat_ & ~new_G2833gat_;
  assign new_G2950gat_ = ~new_G2896gat_ & ~new_G2838gat_;
  assign new_G2954gat_ = ~new_G2899gat_ & ~new_G2843gat_;
  assign new_G2958gat_ = ~new_G2902gat_ & ~new_G2848gat_;
  assign new_G2962gat_ = ~new_G2905gat_ & ~new_G2853gat_;
  assign new_G2966gat_ = ~new_G2861gat_ & ~new_G2908gat_;
  assign new_G2967gat_ = ~new_G2908gat_ & ~new_G2858gat_;
  assign new_G2968gat_ = ~new_G2912gat_ & ~new_G2913gat_;
  assign new_G2971gat_ = ~new_G2914gat_ & ~new_G1137gat_;
  assign new_G2975gat_ = ~new_G2870gat_ & ~new_G2917gat_;
  assign new_G2976gat_ = ~new_G2917gat_ & ~new_G1185gat_;
  assign new_G2977gat_ = ~new_G2739gat_ & ~new_G2917gat_;
  assign new_G2980gat_ = ~new_G2921gat_ & ~new_G2922gat_;
  assign new_G2983gat_ = ~new_G1281gat_ & ~new_G2923gat_;
  assign new_G2987gat_ = ~new_G2878gat_ & ~new_G2926gat_;
  assign new_G2988gat_ = ~new_G2926gat_ & ~new_G2808gat_;
  assign new_G2989gat_ = ~new_G2881gat_ & ~new_G2930gat_;
  assign new_G2990gat_ = ~new_G2930gat_ & ~new_G2813gat_;
  assign new_G2991gat_ = ~new_G2884gat_ & ~new_G2934gat_;
  assign new_G2992gat_ = ~new_G2934gat_ & ~new_G2818gat_;
  assign new_G2993gat_ = ~new_G2887gat_ & ~new_G2938gat_;
  assign new_G2994gat_ = ~new_G2938gat_ & ~new_G2823gat_;
  assign new_G2995gat_ = ~new_G2890gat_ & ~new_G2942gat_;
  assign new_G2996gat_ = ~new_G2942gat_ & ~new_G2828gat_;
  assign new_G2997gat_ = ~new_G2893gat_ & ~new_G2946gat_;
  assign new_G2998gat_ = ~new_G2946gat_ & ~new_G2833gat_;
  assign new_G2999gat_ = ~new_G2896gat_ & ~new_G2950gat_;
  assign new_G3000gat_ = ~new_G2950gat_ & ~new_G2838gat_;
  assign new_G3001gat_ = ~new_G2899gat_ & ~new_G2954gat_;
  assign new_G3002gat_ = ~new_G2954gat_ & ~new_G2843gat_;
  assign new_G3003gat_ = ~new_G2902gat_ & ~new_G2958gat_;
  assign new_G3004gat_ = ~new_G2958gat_ & ~new_G2848gat_;
  assign new_G3005gat_ = ~new_G2905gat_ & ~new_G2962gat_;
  assign new_G3006gat_ = ~new_G2962gat_ & ~new_G2853gat_;
  assign new_G3007gat_ = ~new_G2966gat_ & ~new_G2967gat_;
  assign new_G3010gat_ = ~new_G2968gat_ & ~new_G1089gat_;
  assign new_G3014gat_ = ~new_G2914gat_ & ~new_G2971gat_;
  assign new_G3015gat_ = ~new_G2971gat_ & ~new_G1137gat_;
  assign new_G3016gat_ = ~new_G2797gat_ & ~new_G2971gat_;
  assign new_G3019gat_ = ~new_G2975gat_ & ~new_G2976gat_;
  assign new_G3022gat_ = ~new_G2980gat_ & ~new_G2977gat_;
  assign new_G3026gat_ = ~new_G1281gat_ & ~new_G2983gat_;
  assign new_G3027gat_ = ~new_G2983gat_ & ~new_G2923gat_;
  assign new_G3028gat_ = ~new_G2987gat_ & ~new_G2988gat_;
  assign new_G3031gat_ = ~new_G2989gat_ & ~new_G2990gat_;
  assign new_G3034gat_ = ~new_G2991gat_ & ~new_G2992gat_;
  assign new_G3037gat_ = ~new_G2993gat_ & ~new_G2994gat_;
  assign new_G3040gat_ = ~new_G2995gat_ & ~new_G2996gat_;
  assign new_G3043gat_ = ~new_G2997gat_ & ~new_G2998gat_;
  assign new_G3046gat_ = ~new_G2999gat_ & ~new_G3000gat_;
  assign new_G3049gat_ = ~new_G3001gat_ & ~new_G3002gat_;
  assign new_G3052gat_ = ~new_G3003gat_ & ~new_G3004gat_;
  assign new_G3055gat_ = ~new_G3005gat_ & ~new_G3006gat_;
  assign new_G3058gat_ = ~new_G3007gat_ & ~new_G1041gat_;
  assign new_G3062gat_ = ~new_G2968gat_ & ~new_G3010gat_;
  assign new_G3063gat_ = ~new_G3010gat_ & ~new_G1089gat_;
  assign new_G3064gat_ = ~new_G2864gat_ & ~new_G3010gat_;
  assign new_G3067gat_ = ~new_G3014gat_ & ~new_G3015gat_;
  assign new_G3070gat_ = ~new_G3019gat_ & ~new_G3016gat_;
  assign new_G3074gat_ = ~new_G2980gat_ & ~new_G3022gat_;
  assign new_G3075gat_ = ~new_G3022gat_ & ~new_G2977gat_;
  assign new_G3076gat_ = ~new_G3026gat_ & ~new_G3027gat_;
  assign new_G3079gat_ = ~new_G3028gat_ & ~new_G561gat_;
  assign new_G3083gat_ = ~new_G3031gat_ & ~new_G609gat_;
  assign new_G3087gat_ = ~new_G3034gat_ & ~new_G657gat_;
  assign new_G3091gat_ = ~new_G3037gat_ & ~new_G705gat_;
  assign new_G3095gat_ = ~new_G3040gat_ & ~new_G753gat_;
  assign new_G3099gat_ = ~new_G3043gat_ & ~new_G801gat_;
  assign new_G3103gat_ = ~new_G3046gat_ & ~new_G849gat_;
  assign new_G3107gat_ = ~new_G3049gat_ & ~new_G897gat_;
  assign new_G3111gat_ = ~new_G3052gat_ & ~new_G945gat_;
  assign new_G3115gat_ = ~new_G3055gat_ & ~new_G993gat_;
  assign new_G3119gat_ = ~new_G3007gat_ & ~new_G3058gat_;
  assign new_G3120gat_ = ~new_G3058gat_ & ~new_G1041gat_;
  assign new_G3121gat_ = ~new_G2908gat_ & ~new_G3058gat_;
  assign new_G3124gat_ = ~new_G3062gat_ & ~new_G3063gat_;
  assign new_G3127gat_ = ~new_G3067gat_ & ~new_G3064gat_;
  assign new_G3131gat_ = ~new_G3019gat_ & ~new_G3070gat_;
  assign new_G3132gat_ = ~new_G3070gat_ & ~new_G3016gat_;
  assign new_G3133gat_ = ~new_G3074gat_ & ~new_G3075gat_;
  assign new_G3136gat_ = ~new_G3076gat_ & ~new_G1236gat_;
  assign new_G3140gat_ = ~new_G3028gat_ & ~new_G3079gat_;
  assign new_G3141gat_ = ~new_G3079gat_ & ~new_G561gat_;
  assign new_G3142gat_ = ~new_G2926gat_ & ~new_G3079gat_;
  assign new_G3145gat_ = ~new_G3031gat_ & ~new_G3083gat_;
  assign new_G3146gat_ = ~new_G3083gat_ & ~new_G609gat_;
  assign new_G3147gat_ = ~new_G2930gat_ & ~new_G3083gat_;
  assign new_G3150gat_ = ~new_G3034gat_ & ~new_G3087gat_;
  assign new_G3151gat_ = ~new_G3087gat_ & ~new_G657gat_;
  assign new_G3152gat_ = ~new_G2934gat_ & ~new_G3087gat_;
  assign new_G3155gat_ = ~new_G3037gat_ & ~new_G3091gat_;
  assign new_G3156gat_ = ~new_G3091gat_ & ~new_G705gat_;
  assign new_G3157gat_ = ~new_G2938gat_ & ~new_G3091gat_;
  assign new_G3160gat_ = ~new_G3040gat_ & ~new_G3095gat_;
  assign new_G3161gat_ = ~new_G3095gat_ & ~new_G753gat_;
  assign new_G3162gat_ = ~new_G2942gat_ & ~new_G3095gat_;
  assign new_G3165gat_ = ~new_G3043gat_ & ~new_G3099gat_;
  assign new_G3166gat_ = ~new_G3099gat_ & ~new_G801gat_;
  assign new_G3167gat_ = ~new_G2946gat_ & ~new_G3099gat_;
  assign new_G3170gat_ = ~new_G3046gat_ & ~new_G3103gat_;
  assign new_G3171gat_ = ~new_G3103gat_ & ~new_G849gat_;
  assign new_G3172gat_ = ~new_G2950gat_ & ~new_G3103gat_;
  assign new_G3175gat_ = ~new_G3049gat_ & ~new_G3107gat_;
  assign new_G3176gat_ = ~new_G3107gat_ & ~new_G897gat_;
  assign new_G3177gat_ = ~new_G2954gat_ & ~new_G3107gat_;
  assign new_G3180gat_ = ~new_G3052gat_ & ~new_G3111gat_;
  assign new_G3181gat_ = ~new_G3111gat_ & ~new_G945gat_;
  assign new_G3182gat_ = ~new_G2958gat_ & ~new_G3111gat_;
  assign new_G3185gat_ = ~new_G3055gat_ & ~new_G3115gat_;
  assign new_G3186gat_ = ~new_G3115gat_ & ~new_G993gat_;
  assign new_G3187gat_ = ~new_G2962gat_ & ~new_G3115gat_;
  assign new_G3190gat_ = ~new_G3119gat_ & ~new_G3120gat_;
  assign new_G3193gat_ = ~new_G3124gat_ & ~new_G3121gat_;
  assign new_G3197gat_ = ~new_G3067gat_ & ~new_G3127gat_;
  assign new_G3198gat_ = ~new_G3127gat_ & ~new_G3064gat_;
  assign new_G3199gat_ = ~new_G3131gat_ & ~new_G3132gat_;
  assign new_G3202gat_ = ~new_G3133gat_ & ~new_G1188gat_;
  assign new_G3206gat_ = ~new_G3076gat_ & ~new_G3136gat_;
  assign new_G3207gat_ = ~new_G3136gat_ & ~new_G1236gat_;
  assign new_G3208gat_ = ~new_G2983gat_ & ~new_G3136gat_;
  assign G3211gat = ~new_G3140gat_ & ~new_G3141gat_;
  assign new_G3212gat_ = ~new_G3145gat_ & ~new_G3146gat_;
  assign new_G3215gat_ = ~new_G3150gat_ & ~new_G3151gat_;
  assign new_G3218gat_ = ~new_G3155gat_ & ~new_G3156gat_;
  assign new_G3221gat_ = ~new_G3160gat_ & ~new_G3161gat_;
  assign new_G3224gat_ = ~new_G3165gat_ & ~new_G3166gat_;
  assign new_G3227gat_ = ~new_G3170gat_ & ~new_G3171gat_;
  assign new_G3230gat_ = ~new_G3175gat_ & ~new_G3176gat_;
  assign new_G3233gat_ = ~new_G3180gat_ & ~new_G3181gat_;
  assign new_G3236gat_ = ~new_G3185gat_ & ~new_G3186gat_;
  assign new_G3239gat_ = ~new_G3190gat_ & ~new_G3187gat_;
  assign new_G3243gat_ = ~new_G3124gat_ & ~new_G3193gat_;
  assign new_G3244gat_ = ~new_G3193gat_ & ~new_G3121gat_;
  assign new_G3245gat_ = ~new_G3197gat_ & ~new_G3198gat_;
  assign new_G3248gat_ = ~new_G3199gat_ & ~new_G1140gat_;
  assign new_G3252gat_ = ~new_G3133gat_ & ~new_G3202gat_;
  assign new_G3253gat_ = ~new_G3202gat_ & ~new_G1188gat_;
  assign new_G3254gat_ = ~new_G3022gat_ & ~new_G3202gat_;
  assign new_G3257gat_ = ~new_G3206gat_ & ~new_G3207gat_;
  assign new_G3260gat_ = ~new_G1284gat_ & ~new_G3208gat_;
  assign new_G3264gat_ = ~new_G3212gat_ & ~new_G3142gat_;
  assign new_G3268gat_ = ~new_G3215gat_ & ~new_G3147gat_;
  assign new_G3272gat_ = ~new_G3218gat_ & ~new_G3152gat_;
  assign new_G3276gat_ = ~new_G3221gat_ & ~new_G3157gat_;
  assign new_G3280gat_ = ~new_G3224gat_ & ~new_G3162gat_;
  assign new_G3284gat_ = ~new_G3227gat_ & ~new_G3167gat_;
  assign new_G3288gat_ = ~new_G3230gat_ & ~new_G3172gat_;
  assign new_G3292gat_ = ~new_G3233gat_ & ~new_G3177gat_;
  assign new_G3296gat_ = ~new_G3236gat_ & ~new_G3182gat_;
  assign new_G3300gat_ = ~new_G3190gat_ & ~new_G3239gat_;
  assign new_G3301gat_ = ~new_G3239gat_ & ~new_G3187gat_;
  assign new_G3302gat_ = ~new_G3243gat_ & ~new_G3244gat_;
  assign new_G3305gat_ = ~new_G3245gat_ & ~new_G1092gat_;
  assign new_G3309gat_ = ~new_G3199gat_ & ~new_G3248gat_;
  assign new_G3310gat_ = ~new_G3248gat_ & ~new_G1140gat_;
  assign new_G3311gat_ = ~new_G3070gat_ & ~new_G3248gat_;
  assign new_G3314gat_ = ~new_G3252gat_ & ~new_G3253gat_;
  assign new_G3317gat_ = ~new_G3257gat_ & ~new_G3254gat_;
  assign new_G3321gat_ = ~new_G1284gat_ & ~new_G3260gat_;
  assign new_G3322gat_ = ~new_G3260gat_ & ~new_G3208gat_;
  assign new_G3323gat_ = ~new_G3212gat_ & ~new_G3264gat_;
  assign new_G3324gat_ = ~new_G3264gat_ & ~new_G3142gat_;
  assign new_G3325gat_ = ~new_G3215gat_ & ~new_G3268gat_;
  assign new_G3326gat_ = ~new_G3268gat_ & ~new_G3147gat_;
  assign new_G3327gat_ = ~new_G3218gat_ & ~new_G3272gat_;
  assign new_G3328gat_ = ~new_G3272gat_ & ~new_G3152gat_;
  assign new_G3329gat_ = ~new_G3221gat_ & ~new_G3276gat_;
  assign new_G3330gat_ = ~new_G3276gat_ & ~new_G3157gat_;
  assign new_G3331gat_ = ~new_G3224gat_ & ~new_G3280gat_;
  assign new_G3332gat_ = ~new_G3280gat_ & ~new_G3162gat_;
  assign new_G3333gat_ = ~new_G3227gat_ & ~new_G3284gat_;
  assign new_G3334gat_ = ~new_G3284gat_ & ~new_G3167gat_;
  assign new_G3335gat_ = ~new_G3230gat_ & ~new_G3288gat_;
  assign new_G3336gat_ = ~new_G3288gat_ & ~new_G3172gat_;
  assign new_G3337gat_ = ~new_G3233gat_ & ~new_G3292gat_;
  assign new_G3338gat_ = ~new_G3292gat_ & ~new_G3177gat_;
  assign new_G3339gat_ = ~new_G3236gat_ & ~new_G3296gat_;
  assign new_G3340gat_ = ~new_G3296gat_ & ~new_G3182gat_;
  assign new_G3341gat_ = ~new_G3300gat_ & ~new_G3301gat_;
  assign new_G3344gat_ = ~new_G3302gat_ & ~new_G1044gat_;
  assign new_G3348gat_ = ~new_G3245gat_ & ~new_G3305gat_;
  assign new_G3349gat_ = ~new_G3305gat_ & ~new_G1092gat_;
  assign new_G3350gat_ = ~new_G3127gat_ & ~new_G3305gat_;
  assign new_G3353gat_ = ~new_G3309gat_ & ~new_G3310gat_;
  assign new_G3356gat_ = ~new_G3314gat_ & ~new_G3311gat_;
  assign new_G3360gat_ = ~new_G3257gat_ & ~new_G3317gat_;
  assign new_G3361gat_ = ~new_G3317gat_ & ~new_G3254gat_;
  assign new_G3362gat_ = ~new_G3321gat_ & ~new_G3322gat_;
  assign new_G3365gat_ = ~new_G3323gat_ & ~new_G3324gat_;
  assign new_G3368gat_ = ~new_G3325gat_ & ~new_G3326gat_;
  assign new_G3371gat_ = ~new_G3327gat_ & ~new_G3328gat_;
  assign new_G3374gat_ = ~new_G3329gat_ & ~new_G3330gat_;
  assign new_G3377gat_ = ~new_G3331gat_ & ~new_G3332gat_;
  assign new_G3380gat_ = ~new_G3333gat_ & ~new_G3334gat_;
  assign new_G3383gat_ = ~new_G3335gat_ & ~new_G3336gat_;
  assign new_G3386gat_ = ~new_G3337gat_ & ~new_G3338gat_;
  assign new_G3389gat_ = ~new_G3339gat_ & ~new_G3340gat_;
  assign new_G3392gat_ = ~new_G3341gat_ & ~new_G996gat_;
  assign new_G3396gat_ = ~new_G3302gat_ & ~new_G3344gat_;
  assign new_G3397gat_ = ~new_G3344gat_ & ~new_G1044gat_;
  assign new_G3398gat_ = ~new_G3193gat_ & ~new_G3344gat_;
  assign new_G3401gat_ = ~new_G3348gat_ & ~new_G3349gat_;
  assign new_G3404gat_ = ~new_G3353gat_ & ~new_G3350gat_;
  assign new_G3408gat_ = ~new_G3314gat_ & ~new_G3356gat_;
  assign new_G3409gat_ = ~new_G3356gat_ & ~new_G3311gat_;
  assign new_G3410gat_ = ~new_G3360gat_ & ~new_G3361gat_;
  assign new_G3413gat_ = ~new_G3362gat_ & ~new_G1239gat_;
  assign new_G3417gat_ = ~new_G3365gat_ & ~new_G564gat_;
  assign new_G3421gat_ = ~new_G3368gat_ & ~new_G612gat_;
  assign new_G3425gat_ = ~new_G3371gat_ & ~new_G660gat_;
  assign new_G3429gat_ = ~new_G3374gat_ & ~new_G708gat_;
  assign new_G3433gat_ = ~new_G3377gat_ & ~new_G756gat_;
  assign new_G3437gat_ = ~new_G3380gat_ & ~new_G804gat_;
  assign new_G3441gat_ = ~new_G3383gat_ & ~new_G852gat_;
  assign new_G3445gat_ = ~new_G3386gat_ & ~new_G900gat_;
  assign new_G3449gat_ = ~new_G3389gat_ & ~new_G948gat_;
  assign new_G3453gat_ = ~new_G3341gat_ & ~new_G3392gat_;
  assign new_G3454gat_ = ~new_G3392gat_ & ~new_G996gat_;
  assign new_G3455gat_ = ~new_G3239gat_ & ~new_G3392gat_;
  assign new_G3458gat_ = ~new_G3396gat_ & ~new_G3397gat_;
  assign new_G3461gat_ = ~new_G3401gat_ & ~new_G3398gat_;
  assign new_G3465gat_ = ~new_G3353gat_ & ~new_G3404gat_;
  assign new_G3466gat_ = ~new_G3404gat_ & ~new_G3350gat_;
  assign new_G3467gat_ = ~new_G3408gat_ & ~new_G3409gat_;
  assign new_G3470gat_ = ~new_G3410gat_ & ~new_G1191gat_;
  assign new_G3474gat_ = ~new_G3362gat_ & ~new_G3413gat_;
  assign new_G3475gat_ = ~new_G3413gat_ & ~new_G1239gat_;
  assign new_G3476gat_ = ~new_G3260gat_ & ~new_G3413gat_;
  assign new_G3479gat_ = ~new_G3365gat_ & ~new_G3417gat_;
  assign new_G3480gat_ = ~new_G3417gat_ & ~new_G564gat_;
  assign new_G3481gat_ = ~new_G3264gat_ & ~new_G3417gat_;
  assign new_G3484gat_ = ~new_G3368gat_ & ~new_G3421gat_;
  assign new_G3485gat_ = ~new_G3421gat_ & ~new_G612gat_;
  assign new_G3486gat_ = ~new_G3268gat_ & ~new_G3421gat_;
  assign new_G3489gat_ = ~new_G3371gat_ & ~new_G3425gat_;
  assign new_G3490gat_ = ~new_G3425gat_ & ~new_G660gat_;
  assign new_G3491gat_ = ~new_G3272gat_ & ~new_G3425gat_;
  assign new_G3494gat_ = ~new_G3374gat_ & ~new_G3429gat_;
  assign new_G3495gat_ = ~new_G3429gat_ & ~new_G708gat_;
  assign new_G3496gat_ = ~new_G3276gat_ & ~new_G3429gat_;
  assign new_G3499gat_ = ~new_G3377gat_ & ~new_G3433gat_;
  assign new_G3500gat_ = ~new_G3433gat_ & ~new_G756gat_;
  assign new_G3501gat_ = ~new_G3280gat_ & ~new_G3433gat_;
  assign new_G3504gat_ = ~new_G3380gat_ & ~new_G3437gat_;
  assign new_G3505gat_ = ~new_G3437gat_ & ~new_G804gat_;
  assign new_G3506gat_ = ~new_G3284gat_ & ~new_G3437gat_;
  assign new_G3509gat_ = ~new_G3383gat_ & ~new_G3441gat_;
  assign new_G3510gat_ = ~new_G3441gat_ & ~new_G852gat_;
  assign new_G3511gat_ = ~new_G3288gat_ & ~new_G3441gat_;
  assign new_G3514gat_ = ~new_G3386gat_ & ~new_G3445gat_;
  assign new_G3515gat_ = ~new_G3445gat_ & ~new_G900gat_;
  assign new_G3516gat_ = ~new_G3292gat_ & ~new_G3445gat_;
  assign new_G3519gat_ = ~new_G3389gat_ & ~new_G3449gat_;
  assign new_G3520gat_ = ~new_G3449gat_ & ~new_G948gat_;
  assign new_G3521gat_ = ~new_G3296gat_ & ~new_G3449gat_;
  assign new_G3524gat_ = ~new_G3453gat_ & ~new_G3454gat_;
  assign new_G3527gat_ = ~new_G3458gat_ & ~new_G3455gat_;
  assign new_G3531gat_ = ~new_G3401gat_ & ~new_G3461gat_;
  assign new_G3532gat_ = ~new_G3461gat_ & ~new_G3398gat_;
  assign new_G3533gat_ = ~new_G3465gat_ & ~new_G3466gat_;
  assign new_G3536gat_ = ~new_G3467gat_ & ~new_G1143gat_;
  assign new_G3540gat_ = ~new_G3410gat_ & ~new_G3470gat_;
  assign new_G3541gat_ = ~new_G3470gat_ & ~new_G1191gat_;
  assign new_G3542gat_ = ~new_G3317gat_ & ~new_G3470gat_;
  assign new_G3545gat_ = ~new_G3474gat_ & ~new_G3475gat_;
  assign new_G3548gat_ = ~new_G1287gat_ & ~new_G3476gat_;
  assign G3552gat = ~new_G3479gat_ & ~new_G3480gat_;
  assign new_G3553gat_ = ~new_G3484gat_ & ~new_G3485gat_;
  assign new_G3556gat_ = ~new_G3489gat_ & ~new_G3490gat_;
  assign new_G3559gat_ = ~new_G3494gat_ & ~new_G3495gat_;
  assign new_G3562gat_ = ~new_G3499gat_ & ~new_G3500gat_;
  assign new_G3565gat_ = ~new_G3504gat_ & ~new_G3505gat_;
  assign new_G3568gat_ = ~new_G3509gat_ & ~new_G3510gat_;
  assign new_G3571gat_ = ~new_G3514gat_ & ~new_G3515gat_;
  assign new_G3574gat_ = ~new_G3519gat_ & ~new_G3520gat_;
  assign new_G3577gat_ = ~new_G3524gat_ & ~new_G3521gat_;
  assign new_G3581gat_ = ~new_G3458gat_ & ~new_G3527gat_;
  assign new_G3582gat_ = ~new_G3527gat_ & ~new_G3455gat_;
  assign new_G3583gat_ = ~new_G3531gat_ & ~new_G3532gat_;
  assign new_G3586gat_ = ~new_G3533gat_ & ~new_G1095gat_;
  assign new_G3590gat_ = ~new_G3467gat_ & ~new_G3536gat_;
  assign new_G3591gat_ = ~new_G3536gat_ & ~new_G1143gat_;
  assign new_G3592gat_ = ~new_G3356gat_ & ~new_G3536gat_;
  assign new_G3595gat_ = ~new_G3540gat_ & ~new_G3541gat_;
  assign new_G3598gat_ = ~new_G3545gat_ & ~new_G3542gat_;
  assign new_G3602gat_ = ~new_G1287gat_ & ~new_G3548gat_;
  assign new_G3603gat_ = ~new_G3548gat_ & ~new_G3476gat_;
  assign new_G3604gat_ = ~new_G3553gat_ & ~new_G3481gat_;
  assign new_G3608gat_ = ~new_G3556gat_ & ~new_G3486gat_;
  assign new_G3612gat_ = ~new_G3559gat_ & ~new_G3491gat_;
  assign new_G3616gat_ = ~new_G3562gat_ & ~new_G3496gat_;
  assign new_G3620gat_ = ~new_G3565gat_ & ~new_G3501gat_;
  assign new_G3624gat_ = ~new_G3568gat_ & ~new_G3506gat_;
  assign new_G3628gat_ = ~new_G3571gat_ & ~new_G3511gat_;
  assign new_G3632gat_ = ~new_G3574gat_ & ~new_G3516gat_;
  assign new_G3636gat_ = ~new_G3524gat_ & ~new_G3577gat_;
  assign new_G3637gat_ = ~new_G3577gat_ & ~new_G3521gat_;
  assign new_G3638gat_ = ~new_G3581gat_ & ~new_G3582gat_;
  assign new_G3641gat_ = ~new_G3583gat_ & ~new_G1047gat_;
  assign new_G3645gat_ = ~new_G3533gat_ & ~new_G3586gat_;
  assign new_G3646gat_ = ~new_G3586gat_ & ~new_G1095gat_;
  assign new_G3647gat_ = ~new_G3404gat_ & ~new_G3586gat_;
  assign new_G3650gat_ = ~new_G3590gat_ & ~new_G3591gat_;
  assign new_G3653gat_ = ~new_G3595gat_ & ~new_G3592gat_;
  assign new_G3657gat_ = ~new_G3545gat_ & ~new_G3598gat_;
  assign new_G3658gat_ = ~new_G3598gat_ & ~new_G3542gat_;
  assign new_G3659gat_ = ~new_G3602gat_ & ~new_G3603gat_;
  assign new_G3662gat_ = ~new_G3553gat_ & ~new_G3604gat_;
  assign new_G3663gat_ = ~new_G3604gat_ & ~new_G3481gat_;
  assign new_G3664gat_ = ~new_G3556gat_ & ~new_G3608gat_;
  assign new_G3665gat_ = ~new_G3608gat_ & ~new_G3486gat_;
  assign new_G3666gat_ = ~new_G3559gat_ & ~new_G3612gat_;
  assign new_G3667gat_ = ~new_G3612gat_ & ~new_G3491gat_;
  assign new_G3668gat_ = ~new_G3562gat_ & ~new_G3616gat_;
  assign new_G3669gat_ = ~new_G3616gat_ & ~new_G3496gat_;
  assign new_G3670gat_ = ~new_G3565gat_ & ~new_G3620gat_;
  assign new_G3671gat_ = ~new_G3620gat_ & ~new_G3501gat_;
  assign new_G3672gat_ = ~new_G3568gat_ & ~new_G3624gat_;
  assign new_G3673gat_ = ~new_G3624gat_ & ~new_G3506gat_;
  assign new_G3674gat_ = ~new_G3571gat_ & ~new_G3628gat_;
  assign new_G3675gat_ = ~new_G3628gat_ & ~new_G3511gat_;
  assign new_G3676gat_ = ~new_G3574gat_ & ~new_G3632gat_;
  assign new_G3677gat_ = ~new_G3632gat_ & ~new_G3516gat_;
  assign new_G3678gat_ = ~new_G3636gat_ & ~new_G3637gat_;
  assign new_G3681gat_ = ~new_G3638gat_ & ~new_G999gat_;
  assign new_G3685gat_ = ~new_G3583gat_ & ~new_G3641gat_;
  assign new_G3686gat_ = ~new_G3641gat_ & ~new_G1047gat_;
  assign new_G3687gat_ = ~new_G3461gat_ & ~new_G3641gat_;
  assign new_G3690gat_ = ~new_G3645gat_ & ~new_G3646gat_;
  assign new_G3693gat_ = ~new_G3650gat_ & ~new_G3647gat_;
  assign new_G3697gat_ = ~new_G3595gat_ & ~new_G3653gat_;
  assign new_G3698gat_ = ~new_G3653gat_ & ~new_G3592gat_;
  assign new_G3699gat_ = ~new_G3657gat_ & ~new_G3658gat_;
  assign new_G3702gat_ = ~new_G3659gat_ & ~new_G1242gat_;
  assign new_G3706gat_ = ~new_G3662gat_ & ~new_G3663gat_;
  assign new_G3709gat_ = ~new_G3664gat_ & ~new_G3665gat_;
  assign new_G3712gat_ = ~new_G3666gat_ & ~new_G3667gat_;
  assign new_G3715gat_ = ~new_G3668gat_ & ~new_G3669gat_;
  assign new_G3718gat_ = ~new_G3670gat_ & ~new_G3671gat_;
  assign new_G3721gat_ = ~new_G3672gat_ & ~new_G3673gat_;
  assign new_G3724gat_ = ~new_G3674gat_ & ~new_G3675gat_;
  assign new_G3727gat_ = ~new_G3676gat_ & ~new_G3677gat_;
  assign new_G3730gat_ = ~new_G3678gat_ & ~new_G951gat_;
  assign new_G3734gat_ = ~new_G3638gat_ & ~new_G3681gat_;
  assign new_G3735gat_ = ~new_G3681gat_ & ~new_G999gat_;
  assign new_G3736gat_ = ~new_G3527gat_ & ~new_G3681gat_;
  assign new_G3739gat_ = ~new_G3685gat_ & ~new_G3686gat_;
  assign new_G3742gat_ = ~new_G3690gat_ & ~new_G3687gat_;
  assign new_G3746gat_ = ~new_G3650gat_ & ~new_G3693gat_;
  assign new_G3747gat_ = ~new_G3693gat_ & ~new_G3647gat_;
  assign new_G3748gat_ = ~new_G3697gat_ & ~new_G3698gat_;
  assign new_G3751gat_ = ~new_G3699gat_ & ~new_G1194gat_;
  assign new_G3755gat_ = ~new_G3659gat_ & ~new_G3702gat_;
  assign new_G3756gat_ = ~new_G3702gat_ & ~new_G1242gat_;
  assign new_G3757gat_ = ~new_G3548gat_ & ~new_G3702gat_;
  assign new_G3760gat_ = ~new_G3706gat_ & ~new_G567gat_;
  assign new_G3764gat_ = ~new_G3709gat_ & ~new_G615gat_;
  assign new_G3768gat_ = ~new_G3712gat_ & ~new_G663gat_;
  assign new_G3772gat_ = ~new_G3715gat_ & ~new_G711gat_;
  assign new_G3776gat_ = ~new_G3718gat_ & ~new_G759gat_;
  assign new_G3780gat_ = ~new_G3721gat_ & ~new_G807gat_;
  assign new_G3784gat_ = ~new_G3724gat_ & ~new_G855gat_;
  assign new_G3788gat_ = ~new_G3727gat_ & ~new_G903gat_;
  assign new_G3792gat_ = ~new_G3678gat_ & ~new_G3730gat_;
  assign new_G3793gat_ = ~new_G3730gat_ & ~new_G951gat_;
  assign new_G3794gat_ = ~new_G3577gat_ & ~new_G3730gat_;
  assign new_G3797gat_ = ~new_G3734gat_ & ~new_G3735gat_;
  assign new_G3800gat_ = ~new_G3739gat_ & ~new_G3736gat_;
  assign new_G3804gat_ = ~new_G3690gat_ & ~new_G3742gat_;
  assign new_G3805gat_ = ~new_G3742gat_ & ~new_G3687gat_;
  assign new_G3806gat_ = ~new_G3746gat_ & ~new_G3747gat_;
  assign new_G3809gat_ = ~new_G3748gat_ & ~new_G1146gat_;
  assign new_G3813gat_ = ~new_G3699gat_ & ~new_G3751gat_;
  assign new_G3814gat_ = ~new_G3751gat_ & ~new_G1194gat_;
  assign new_G3815gat_ = ~new_G3598gat_ & ~new_G3751gat_;
  assign new_G3818gat_ = ~new_G3755gat_ & ~new_G3756gat_;
  assign new_G3821gat_ = ~new_G1290gat_ & ~new_G3757gat_;
  assign new_G3825gat_ = ~new_G3706gat_ & ~new_G3760gat_;
  assign new_G3826gat_ = ~new_G3760gat_ & ~new_G567gat_;
  assign new_G3827gat_ = ~new_G3604gat_ & ~new_G3760gat_;
  assign new_G3830gat_ = ~new_G3709gat_ & ~new_G3764gat_;
  assign new_G3831gat_ = ~new_G3764gat_ & ~new_G615gat_;
  assign new_G3832gat_ = ~new_G3608gat_ & ~new_G3764gat_;
  assign new_G3835gat_ = ~new_G3712gat_ & ~new_G3768gat_;
  assign new_G3836gat_ = ~new_G3768gat_ & ~new_G663gat_;
  assign new_G3837gat_ = ~new_G3612gat_ & ~new_G3768gat_;
  assign new_G3840gat_ = ~new_G3715gat_ & ~new_G3772gat_;
  assign new_G3841gat_ = ~new_G3772gat_ & ~new_G711gat_;
  assign new_G3842gat_ = ~new_G3616gat_ & ~new_G3772gat_;
  assign new_G3845gat_ = ~new_G3718gat_ & ~new_G3776gat_;
  assign new_G3846gat_ = ~new_G3776gat_ & ~new_G759gat_;
  assign new_G3847gat_ = ~new_G3620gat_ & ~new_G3776gat_;
  assign new_G3850gat_ = ~new_G3721gat_ & ~new_G3780gat_;
  assign new_G3851gat_ = ~new_G3780gat_ & ~new_G807gat_;
  assign new_G3852gat_ = ~new_G3624gat_ & ~new_G3780gat_;
  assign new_G3855gat_ = ~new_G3724gat_ & ~new_G3784gat_;
  assign new_G3856gat_ = ~new_G3784gat_ & ~new_G855gat_;
  assign new_G3857gat_ = ~new_G3628gat_ & ~new_G3784gat_;
  assign new_G3860gat_ = ~new_G3727gat_ & ~new_G3788gat_;
  assign new_G3861gat_ = ~new_G3788gat_ & ~new_G903gat_;
  assign new_G3862gat_ = ~new_G3632gat_ & ~new_G3788gat_;
  assign new_G3865gat_ = ~new_G3792gat_ & ~new_G3793gat_;
  assign new_G3868gat_ = ~new_G3797gat_ & ~new_G3794gat_;
  assign new_G3872gat_ = ~new_G3739gat_ & ~new_G3800gat_;
  assign new_G3873gat_ = ~new_G3800gat_ & ~new_G3736gat_;
  assign new_G3874gat_ = ~new_G3804gat_ & ~new_G3805gat_;
  assign new_G3877gat_ = ~new_G3806gat_ & ~new_G1098gat_;
  assign new_G3881gat_ = ~new_G3748gat_ & ~new_G3809gat_;
  assign new_G3882gat_ = ~new_G3809gat_ & ~new_G1146gat_;
  assign new_G3883gat_ = ~new_G3653gat_ & ~new_G3809gat_;
  assign new_G3886gat_ = ~new_G3813gat_ & ~new_G3814gat_;
  assign new_G3889gat_ = ~new_G3818gat_ & ~new_G3815gat_;
  assign new_G3893gat_ = ~new_G1290gat_ & ~new_G3821gat_;
  assign new_G3894gat_ = ~new_G3821gat_ & ~new_G3757gat_;
  assign G3895gat = ~new_G3825gat_ & ~new_G3826gat_;
  assign new_G3896gat_ = ~new_G3830gat_ & ~new_G3831gat_;
  assign new_G3899gat_ = ~new_G3835gat_ & ~new_G3836gat_;
  assign new_G3902gat_ = ~new_G3840gat_ & ~new_G3841gat_;
  assign new_G3905gat_ = ~new_G3845gat_ & ~new_G3846gat_;
  assign new_G3908gat_ = ~new_G3850gat_ & ~new_G3851gat_;
  assign new_G3911gat_ = ~new_G3855gat_ & ~new_G3856gat_;
  assign new_G3914gat_ = ~new_G3860gat_ & ~new_G3861gat_;
  assign new_G3917gat_ = ~new_G3865gat_ & ~new_G3862gat_;
  assign new_G3921gat_ = ~new_G3797gat_ & ~new_G3868gat_;
  assign new_G3922gat_ = ~new_G3868gat_ & ~new_G3794gat_;
  assign new_G3923gat_ = ~new_G3872gat_ & ~new_G3873gat_;
  assign new_G3926gat_ = ~new_G3874gat_ & ~new_G1050gat_;
  assign new_G3930gat_ = ~new_G3806gat_ & ~new_G3877gat_;
  assign new_G3931gat_ = ~new_G3877gat_ & ~new_G1098gat_;
  assign new_G3932gat_ = ~new_G3693gat_ & ~new_G3877gat_;
  assign new_G3935gat_ = ~new_G3881gat_ & ~new_G3882gat_;
  assign new_G3938gat_ = ~new_G3886gat_ & ~new_G3883gat_;
  assign new_G3942gat_ = ~new_G3818gat_ & ~new_G3889gat_;
  assign new_G3943gat_ = ~new_G3889gat_ & ~new_G3815gat_;
  assign new_G3944gat_ = ~new_G3893gat_ & ~new_G3894gat_;
  assign new_G3947gat_ = ~new_G3896gat_ & ~new_G3827gat_;
  assign new_G3951gat_ = ~new_G3899gat_ & ~new_G3832gat_;
  assign new_G3955gat_ = ~new_G3902gat_ & ~new_G3837gat_;
  assign new_G3959gat_ = ~new_G3905gat_ & ~new_G3842gat_;
  assign new_G3963gat_ = ~new_G3908gat_ & ~new_G3847gat_;
  assign new_G3967gat_ = ~new_G3911gat_ & ~new_G3852gat_;
  assign new_G3971gat_ = ~new_G3914gat_ & ~new_G3857gat_;
  assign new_G3975gat_ = ~new_G3865gat_ & ~new_G3917gat_;
  assign new_G3976gat_ = ~new_G3917gat_ & ~new_G3862gat_;
  assign new_G3977gat_ = ~new_G3921gat_ & ~new_G3922gat_;
  assign new_G3980gat_ = ~new_G3923gat_ & ~new_G1002gat_;
  assign new_G3984gat_ = ~new_G3874gat_ & ~new_G3926gat_;
  assign new_G3985gat_ = ~new_G3926gat_ & ~new_G1050gat_;
  assign new_G3986gat_ = ~new_G3742gat_ & ~new_G3926gat_;
  assign new_G3989gat_ = ~new_G3930gat_ & ~new_G3931gat_;
  assign new_G3992gat_ = ~new_G3935gat_ & ~new_G3932gat_;
  assign new_G3996gat_ = ~new_G3886gat_ & ~new_G3938gat_;
  assign new_G3997gat_ = ~new_G3938gat_ & ~new_G3883gat_;
  assign new_G3998gat_ = ~new_G3942gat_ & ~new_G3943gat_;
  assign new_G4001gat_ = ~new_G3944gat_ & ~new_G1245gat_;
  assign new_G4005gat_ = ~new_G3896gat_ & ~new_G3947gat_;
  assign new_G4006gat_ = ~new_G3947gat_ & ~new_G3827gat_;
  assign new_G4007gat_ = ~new_G3899gat_ & ~new_G3951gat_;
  assign new_G4008gat_ = ~new_G3951gat_ & ~new_G3832gat_;
  assign new_G4009gat_ = ~new_G3902gat_ & ~new_G3955gat_;
  assign new_G4010gat_ = ~new_G3955gat_ & ~new_G3837gat_;
  assign new_G4011gat_ = ~new_G3905gat_ & ~new_G3959gat_;
  assign new_G4012gat_ = ~new_G3959gat_ & ~new_G3842gat_;
  assign new_G4013gat_ = ~new_G3908gat_ & ~new_G3963gat_;
  assign new_G4014gat_ = ~new_G3963gat_ & ~new_G3847gat_;
  assign new_G4015gat_ = ~new_G3911gat_ & ~new_G3967gat_;
  assign new_G4016gat_ = ~new_G3967gat_ & ~new_G3852gat_;
  assign new_G4017gat_ = ~new_G3914gat_ & ~new_G3971gat_;
  assign new_G4018gat_ = ~new_G3971gat_ & ~new_G3857gat_;
  assign new_G4019gat_ = ~new_G3975gat_ & ~new_G3976gat_;
  assign new_G4022gat_ = ~new_G3977gat_ & ~new_G954gat_;
  assign new_G4026gat_ = ~new_G3923gat_ & ~new_G3980gat_;
  assign new_G4027gat_ = ~new_G3980gat_ & ~new_G1002gat_;
  assign new_G4028gat_ = ~new_G3800gat_ & ~new_G3980gat_;
  assign new_G4031gat_ = ~new_G3984gat_ & ~new_G3985gat_;
  assign new_G4034gat_ = ~new_G3989gat_ & ~new_G3986gat_;
  assign new_G4038gat_ = ~new_G3935gat_ & ~new_G3992gat_;
  assign new_G4039gat_ = ~new_G3992gat_ & ~new_G3932gat_;
  assign new_G4040gat_ = ~new_G3996gat_ & ~new_G3997gat_;
  assign new_G4043gat_ = ~new_G3998gat_ & ~new_G1197gat_;
  assign new_G4047gat_ = ~new_G3944gat_ & ~new_G4001gat_;
  assign new_G4048gat_ = ~new_G4001gat_ & ~new_G1245gat_;
  assign new_G4049gat_ = ~new_G3821gat_ & ~new_G4001gat_;
  assign new_G4052gat_ = ~new_G4005gat_ & ~new_G4006gat_;
  assign new_G4055gat_ = ~new_G4007gat_ & ~new_G4008gat_;
  assign new_G4058gat_ = ~new_G4009gat_ & ~new_G4010gat_;
  assign new_G4061gat_ = ~new_G4011gat_ & ~new_G4012gat_;
  assign new_G4064gat_ = ~new_G4013gat_ & ~new_G4014gat_;
  assign new_G4067gat_ = ~new_G4015gat_ & ~new_G4016gat_;
  assign new_G4070gat_ = ~new_G4017gat_ & ~new_G4018gat_;
  assign new_G4073gat_ = ~new_G4019gat_ & ~new_G906gat_;
  assign new_G4077gat_ = ~new_G3977gat_ & ~new_G4022gat_;
  assign new_G4078gat_ = ~new_G4022gat_ & ~new_G954gat_;
  assign new_G4079gat_ = ~new_G3868gat_ & ~new_G4022gat_;
  assign new_G4082gat_ = ~new_G4026gat_ & ~new_G4027gat_;
  assign new_G4085gat_ = ~new_G4031gat_ & ~new_G4028gat_;
  assign new_G4089gat_ = ~new_G3989gat_ & ~new_G4034gat_;
  assign new_G4090gat_ = ~new_G4034gat_ & ~new_G3986gat_;
  assign new_G4091gat_ = ~new_G4038gat_ & ~new_G4039gat_;
  assign new_G4094gat_ = ~new_G4040gat_ & ~new_G1149gat_;
  assign new_G4098gat_ = ~new_G3998gat_ & ~new_G4043gat_;
  assign new_G4099gat_ = ~new_G4043gat_ & ~new_G1197gat_;
  assign new_G4100gat_ = ~new_G3889gat_ & ~new_G4043gat_;
  assign new_G4103gat_ = ~new_G4047gat_ & ~new_G4048gat_;
  assign new_G4106gat_ = ~new_G1293gat_ & ~new_G4049gat_;
  assign new_G4110gat_ = ~new_G4052gat_ & ~new_G570gat_;
  assign new_G4114gat_ = ~new_G4055gat_ & ~new_G618gat_;
  assign new_G4118gat_ = ~new_G4058gat_ & ~new_G666gat_;
  assign new_G4122gat_ = ~new_G4061gat_ & ~new_G714gat_;
  assign new_G4126gat_ = ~new_G4064gat_ & ~new_G762gat_;
  assign new_G4130gat_ = ~new_G4067gat_ & ~new_G810gat_;
  assign new_G4134gat_ = ~new_G4070gat_ & ~new_G858gat_;
  assign new_G4138gat_ = ~new_G4019gat_ & ~new_G4073gat_;
  assign new_G4139gat_ = ~new_G4073gat_ & ~new_G906gat_;
  assign new_G4140gat_ = ~new_G3917gat_ & ~new_G4073gat_;
  assign new_G4143gat_ = ~new_G4077gat_ & ~new_G4078gat_;
  assign new_G4146gat_ = ~new_G4082gat_ & ~new_G4079gat_;
  assign new_G4150gat_ = ~new_G4031gat_ & ~new_G4085gat_;
  assign new_G4151gat_ = ~new_G4085gat_ & ~new_G4028gat_;
  assign new_G4152gat_ = ~new_G4089gat_ & ~new_G4090gat_;
  assign new_G4155gat_ = ~new_G4091gat_ & ~new_G1101gat_;
  assign new_G4159gat_ = ~new_G4040gat_ & ~new_G4094gat_;
  assign new_G4160gat_ = ~new_G4094gat_ & ~new_G1149gat_;
  assign new_G4161gat_ = ~new_G3938gat_ & ~new_G4094gat_;
  assign new_G4164gat_ = ~new_G4098gat_ & ~new_G4099gat_;
  assign new_G4167gat_ = ~new_G4103gat_ & ~new_G4100gat_;
  assign new_G4171gat_ = ~new_G1293gat_ & ~new_G4106gat_;
  assign new_G4172gat_ = ~new_G4106gat_ & ~new_G4049gat_;
  assign new_G4173gat_ = ~new_G4052gat_ & ~new_G4110gat_;
  assign new_G4174gat_ = ~new_G4110gat_ & ~new_G570gat_;
  assign new_G4175gat_ = ~new_G3947gat_ & ~new_G4110gat_;
  assign new_G4178gat_ = ~new_G4055gat_ & ~new_G4114gat_;
  assign new_G4179gat_ = ~new_G4114gat_ & ~new_G618gat_;
  assign new_G4180gat_ = ~new_G3951gat_ & ~new_G4114gat_;
  assign new_G4183gat_ = ~new_G4058gat_ & ~new_G4118gat_;
  assign new_G4184gat_ = ~new_G4118gat_ & ~new_G666gat_;
  assign new_G4185gat_ = ~new_G3955gat_ & ~new_G4118gat_;
  assign new_G4188gat_ = ~new_G4061gat_ & ~new_G4122gat_;
  assign new_G4189gat_ = ~new_G4122gat_ & ~new_G714gat_;
  assign new_G4190gat_ = ~new_G3959gat_ & ~new_G4122gat_;
  assign new_G4193gat_ = ~new_G4064gat_ & ~new_G4126gat_;
  assign new_G4194gat_ = ~new_G4126gat_ & ~new_G762gat_;
  assign new_G4195gat_ = ~new_G3963gat_ & ~new_G4126gat_;
  assign new_G4198gat_ = ~new_G4067gat_ & ~new_G4130gat_;
  assign new_G4199gat_ = ~new_G4130gat_ & ~new_G810gat_;
  assign new_G4200gat_ = ~new_G3967gat_ & ~new_G4130gat_;
  assign new_G4203gat_ = ~new_G4070gat_ & ~new_G4134gat_;
  assign new_G4204gat_ = ~new_G4134gat_ & ~new_G858gat_;
  assign new_G4205gat_ = ~new_G3971gat_ & ~new_G4134gat_;
  assign new_G4208gat_ = ~new_G4138gat_ & ~new_G4139gat_;
  assign new_G4211gat_ = ~new_G4143gat_ & ~new_G4140gat_;
  assign new_G4215gat_ = ~new_G4082gat_ & ~new_G4146gat_;
  assign new_G4216gat_ = ~new_G4146gat_ & ~new_G4079gat_;
  assign new_G4217gat_ = ~new_G4150gat_ & ~new_G4151gat_;
  assign new_G4220gat_ = ~new_G4152gat_ & ~new_G1053gat_;
  assign new_G4224gat_ = ~new_G4091gat_ & ~new_G4155gat_;
  assign new_G4225gat_ = ~new_G4155gat_ & ~new_G1101gat_;
  assign new_G4226gat_ = ~new_G3992gat_ & ~new_G4155gat_;
  assign new_G4229gat_ = ~new_G4159gat_ & ~new_G4160gat_;
  assign new_G4232gat_ = ~new_G4164gat_ & ~new_G4161gat_;
  assign new_G4236gat_ = ~new_G4103gat_ & ~new_G4167gat_;
  assign new_G4237gat_ = ~new_G4167gat_ & ~new_G4100gat_;
  assign new_G4238gat_ = ~new_G4171gat_ & ~new_G4172gat_;
  assign G4241gat = ~new_G4173gat_ & ~new_G4174gat_;
  assign new_G4242gat_ = ~new_G4178gat_ & ~new_G4179gat_;
  assign new_G4245gat_ = ~new_G4183gat_ & ~new_G4184gat_;
  assign new_G4248gat_ = ~new_G4188gat_ & ~new_G4189gat_;
  assign new_G4251gat_ = ~new_G4193gat_ & ~new_G4194gat_;
  assign new_G4254gat_ = ~new_G4198gat_ & ~new_G4199gat_;
  assign new_G4257gat_ = ~new_G4203gat_ & ~new_G4204gat_;
  assign new_G4260gat_ = ~new_G4208gat_ & ~new_G4205gat_;
  assign new_G4264gat_ = ~new_G4143gat_ & ~new_G4211gat_;
  assign new_G4265gat_ = ~new_G4211gat_ & ~new_G4140gat_;
  assign new_G4266gat_ = ~new_G4215gat_ & ~new_G4216gat_;
  assign new_G4269gat_ = ~new_G4217gat_ & ~new_G1005gat_;
  assign new_G4273gat_ = ~new_G4152gat_ & ~new_G4220gat_;
  assign new_G4274gat_ = ~new_G4220gat_ & ~new_G1053gat_;
  assign new_G4275gat_ = ~new_G4034gat_ & ~new_G4220gat_;
  assign new_G4278gat_ = ~new_G4224gat_ & ~new_G4225gat_;
  assign new_G4281gat_ = ~new_G4229gat_ & ~new_G4226gat_;
  assign new_G4285gat_ = ~new_G4164gat_ & ~new_G4232gat_;
  assign new_G4286gat_ = ~new_G4232gat_ & ~new_G4161gat_;
  assign new_G4287gat_ = ~new_G4236gat_ & ~new_G4237gat_;
  assign new_G4290gat_ = ~new_G4238gat_ & ~new_G1248gat_;
  assign new_G4294gat_ = ~new_G4242gat_ & ~new_G4175gat_;
  assign new_G4298gat_ = ~new_G4245gat_ & ~new_G4180gat_;
  assign new_G4302gat_ = ~new_G4248gat_ & ~new_G4185gat_;
  assign new_G4306gat_ = ~new_G4251gat_ & ~new_G4190gat_;
  assign new_G4310gat_ = ~new_G4254gat_ & ~new_G4195gat_;
  assign new_G4314gat_ = ~new_G4257gat_ & ~new_G4200gat_;
  assign new_G4318gat_ = ~new_G4208gat_ & ~new_G4260gat_;
  assign new_G4319gat_ = ~new_G4260gat_ & ~new_G4205gat_;
  assign new_G4320gat_ = ~new_G4264gat_ & ~new_G4265gat_;
  assign new_G4323gat_ = ~new_G4266gat_ & ~new_G957gat_;
  assign new_G4327gat_ = ~new_G4217gat_ & ~new_G4269gat_;
  assign new_G4328gat_ = ~new_G4269gat_ & ~new_G1005gat_;
  assign new_G4329gat_ = ~new_G4085gat_ & ~new_G4269gat_;
  assign new_G4332gat_ = ~new_G4273gat_ & ~new_G4274gat_;
  assign new_G4335gat_ = ~new_G4278gat_ & ~new_G4275gat_;
  assign new_G4339gat_ = ~new_G4229gat_ & ~new_G4281gat_;
  assign new_G4340gat_ = ~new_G4281gat_ & ~new_G4226gat_;
  assign new_G4341gat_ = ~new_G4285gat_ & ~new_G4286gat_;
  assign new_G4344gat_ = ~new_G4287gat_ & ~new_G1200gat_;
  assign new_G4348gat_ = ~new_G4238gat_ & ~new_G4290gat_;
  assign new_G4349gat_ = ~new_G4290gat_ & ~new_G1248gat_;
  assign new_G4350gat_ = ~new_G4106gat_ & ~new_G4290gat_;
  assign new_G4353gat_ = ~new_G4242gat_ & ~new_G4294gat_;
  assign new_G4354gat_ = ~new_G4294gat_ & ~new_G4175gat_;
  assign new_G4355gat_ = ~new_G4245gat_ & ~new_G4298gat_;
  assign new_G4356gat_ = ~new_G4298gat_ & ~new_G4180gat_;
  assign new_G4357gat_ = ~new_G4248gat_ & ~new_G4302gat_;
  assign new_G4358gat_ = ~new_G4302gat_ & ~new_G4185gat_;
  assign new_G4359gat_ = ~new_G4251gat_ & ~new_G4306gat_;
  assign new_G4360gat_ = ~new_G4306gat_ & ~new_G4190gat_;
  assign new_G4361gat_ = ~new_G4254gat_ & ~new_G4310gat_;
  assign new_G4362gat_ = ~new_G4310gat_ & ~new_G4195gat_;
  assign new_G4363gat_ = ~new_G4257gat_ & ~new_G4314gat_;
  assign new_G4364gat_ = ~new_G4314gat_ & ~new_G4200gat_;
  assign new_G4365gat_ = ~new_G4318gat_ & ~new_G4319gat_;
  assign new_G4368gat_ = ~new_G4320gat_ & ~new_G909gat_;
  assign new_G4372gat_ = ~new_G4266gat_ & ~new_G4323gat_;
  assign new_G4373gat_ = ~new_G4323gat_ & ~new_G957gat_;
  assign new_G4374gat_ = ~new_G4146gat_ & ~new_G4323gat_;
  assign new_G4377gat_ = ~new_G4327gat_ & ~new_G4328gat_;
  assign new_G4380gat_ = ~new_G4332gat_ & ~new_G4329gat_;
  assign new_G4384gat_ = ~new_G4278gat_ & ~new_G4335gat_;
  assign new_G4385gat_ = ~new_G4335gat_ & ~new_G4275gat_;
  assign new_G4386gat_ = ~new_G4339gat_ & ~new_G4340gat_;
  assign new_G4389gat_ = ~new_G4341gat_ & ~new_G1152gat_;
  assign new_G4393gat_ = ~new_G4287gat_ & ~new_G4344gat_;
  assign new_G4394gat_ = ~new_G4344gat_ & ~new_G1200gat_;
  assign new_G4395gat_ = ~new_G4167gat_ & ~new_G4344gat_;
  assign new_G4398gat_ = ~new_G4348gat_ & ~new_G4349gat_;
  assign new_G4401gat_ = ~new_G1296gat_ & ~new_G4350gat_;
  assign new_G4405gat_ = ~new_G4353gat_ & ~new_G4354gat_;
  assign new_G4408gat_ = ~new_G4355gat_ & ~new_G4356gat_;
  assign new_G4411gat_ = ~new_G4357gat_ & ~new_G4358gat_;
  assign new_G4414gat_ = ~new_G4359gat_ & ~new_G4360gat_;
  assign new_G4417gat_ = ~new_G4361gat_ & ~new_G4362gat_;
  assign new_G4420gat_ = ~new_G4363gat_ & ~new_G4364gat_;
  assign new_G4423gat_ = ~new_G4365gat_ & ~new_G861gat_;
  assign new_G4427gat_ = ~new_G4320gat_ & ~new_G4368gat_;
  assign new_G4428gat_ = ~new_G4368gat_ & ~new_G909gat_;
  assign new_G4429gat_ = ~new_G4211gat_ & ~new_G4368gat_;
  assign new_G4432gat_ = ~new_G4372gat_ & ~new_G4373gat_;
  assign new_G4435gat_ = ~new_G4377gat_ & ~new_G4374gat_;
  assign new_G4439gat_ = ~new_G4332gat_ & ~new_G4380gat_;
  assign new_G4440gat_ = ~new_G4380gat_ & ~new_G4329gat_;
  assign new_G4441gat_ = ~new_G4384gat_ & ~new_G4385gat_;
  assign new_G4444gat_ = ~new_G4386gat_ & ~new_G1104gat_;
  assign new_G4448gat_ = ~new_G4341gat_ & ~new_G4389gat_;
  assign new_G4449gat_ = ~new_G4389gat_ & ~new_G1152gat_;
  assign new_G4450gat_ = ~new_G4232gat_ & ~new_G4389gat_;
  assign new_G4453gat_ = ~new_G4393gat_ & ~new_G4394gat_;
  assign new_G4456gat_ = ~new_G4398gat_ & ~new_G4395gat_;
  assign new_G4460gat_ = ~new_G1296gat_ & ~new_G4401gat_;
  assign new_G4461gat_ = ~new_G4401gat_ & ~new_G4350gat_;
  assign new_G4462gat_ = ~new_G4405gat_ & ~new_G573gat_;
  assign new_G4466gat_ = ~new_G4408gat_ & ~new_G621gat_;
  assign new_G4470gat_ = ~new_G4411gat_ & ~new_G669gat_;
  assign new_G4474gat_ = ~new_G4414gat_ & ~new_G717gat_;
  assign new_G4478gat_ = ~new_G4417gat_ & ~new_G765gat_;
  assign new_G4482gat_ = ~new_G4420gat_ & ~new_G813gat_;
  assign new_G4486gat_ = ~new_G4365gat_ & ~new_G4423gat_;
  assign new_G4487gat_ = ~new_G4423gat_ & ~new_G861gat_;
  assign new_G4488gat_ = ~new_G4260gat_ & ~new_G4423gat_;
  assign new_G4491gat_ = ~new_G4427gat_ & ~new_G4428gat_;
  assign new_G4494gat_ = ~new_G4432gat_ & ~new_G4429gat_;
  assign new_G4498gat_ = ~new_G4377gat_ & ~new_G4435gat_;
  assign new_G4499gat_ = ~new_G4435gat_ & ~new_G4374gat_;
  assign new_G4500gat_ = ~new_G4439gat_ & ~new_G4440gat_;
  assign new_G4503gat_ = ~new_G4441gat_ & ~new_G1056gat_;
  assign new_G4507gat_ = ~new_G4386gat_ & ~new_G4444gat_;
  assign new_G4508gat_ = ~new_G4444gat_ & ~new_G1104gat_;
  assign new_G4509gat_ = ~new_G4281gat_ & ~new_G4444gat_;
  assign new_G4512gat_ = ~new_G4448gat_ & ~new_G4449gat_;
  assign new_G4515gat_ = ~new_G4453gat_ & ~new_G4450gat_;
  assign new_G4519gat_ = ~new_G4398gat_ & ~new_G4456gat_;
  assign new_G4520gat_ = ~new_G4456gat_ & ~new_G4395gat_;
  assign new_G4521gat_ = ~new_G4460gat_ & ~new_G4461gat_;
  assign new_G4524gat_ = ~new_G4405gat_ & ~new_G4462gat_;
  assign new_G4525gat_ = ~new_G4462gat_ & ~new_G573gat_;
  assign new_G4526gat_ = ~new_G4294gat_ & ~new_G4462gat_;
  assign new_G4529gat_ = ~new_G4408gat_ & ~new_G4466gat_;
  assign new_G4530gat_ = ~new_G4466gat_ & ~new_G621gat_;
  assign new_G4531gat_ = ~new_G4298gat_ & ~new_G4466gat_;
  assign new_G4534gat_ = ~new_G4411gat_ & ~new_G4470gat_;
  assign new_G4535gat_ = ~new_G4470gat_ & ~new_G669gat_;
  assign new_G4536gat_ = ~new_G4302gat_ & ~new_G4470gat_;
  assign new_G4539gat_ = ~new_G4414gat_ & ~new_G4474gat_;
  assign new_G4540gat_ = ~new_G4474gat_ & ~new_G717gat_;
  assign new_G4541gat_ = ~new_G4306gat_ & ~new_G4474gat_;
  assign new_G4544gat_ = ~new_G4417gat_ & ~new_G4478gat_;
  assign new_G4545gat_ = ~new_G4478gat_ & ~new_G765gat_;
  assign new_G4546gat_ = ~new_G4310gat_ & ~new_G4478gat_;
  assign new_G4549gat_ = ~new_G4420gat_ & ~new_G4482gat_;
  assign new_G4550gat_ = ~new_G4482gat_ & ~new_G813gat_;
  assign new_G4551gat_ = ~new_G4314gat_ & ~new_G4482gat_;
  assign new_G4554gat_ = ~new_G4486gat_ & ~new_G4487gat_;
  assign new_G4557gat_ = ~new_G4491gat_ & ~new_G4488gat_;
  assign new_G4561gat_ = ~new_G4432gat_ & ~new_G4494gat_;
  assign new_G4562gat_ = ~new_G4494gat_ & ~new_G4429gat_;
  assign new_G4563gat_ = ~new_G4498gat_ & ~new_G4499gat_;
  assign new_G4566gat_ = ~new_G4500gat_ & ~new_G1008gat_;
  assign new_G4570gat_ = ~new_G4441gat_ & ~new_G4503gat_;
  assign new_G4571gat_ = ~new_G4503gat_ & ~new_G1056gat_;
  assign new_G4572gat_ = ~new_G4335gat_ & ~new_G4503gat_;
  assign new_G4575gat_ = ~new_G4507gat_ & ~new_G4508gat_;
  assign new_G4578gat_ = ~new_G4512gat_ & ~new_G4509gat_;
  assign new_G4582gat_ = ~new_G4453gat_ & ~new_G4515gat_;
  assign new_G4583gat_ = ~new_G4515gat_ & ~new_G4450gat_;
  assign new_G4584gat_ = ~new_G4519gat_ & ~new_G4520gat_;
  assign new_G4587gat_ = ~new_G4521gat_ & ~new_G1251gat_;
  assign G4591gat = ~new_G4524gat_ & ~new_G4525gat_;
  assign new_G4592gat_ = ~new_G4529gat_ & ~new_G4530gat_;
  assign new_G4595gat_ = ~new_G4534gat_ & ~new_G4535gat_;
  assign new_G4598gat_ = ~new_G4539gat_ & ~new_G4540gat_;
  assign new_G4601gat_ = ~new_G4544gat_ & ~new_G4545gat_;
  assign new_G4604gat_ = ~new_G4549gat_ & ~new_G4550gat_;
  assign new_G4607gat_ = ~new_G4554gat_ & ~new_G4551gat_;
  assign new_G4611gat_ = ~new_G4491gat_ & ~new_G4557gat_;
  assign new_G4612gat_ = ~new_G4557gat_ & ~new_G4488gat_;
  assign new_G4613gat_ = ~new_G4561gat_ & ~new_G4562gat_;
  assign new_G4616gat_ = ~new_G4563gat_ & ~new_G960gat_;
  assign new_G4620gat_ = ~new_G4500gat_ & ~new_G4566gat_;
  assign new_G4621gat_ = ~new_G4566gat_ & ~new_G1008gat_;
  assign new_G4622gat_ = ~new_G4380gat_ & ~new_G4566gat_;
  assign new_G4625gat_ = ~new_G4570gat_ & ~new_G4571gat_;
  assign new_G4628gat_ = ~new_G4575gat_ & ~new_G4572gat_;
  assign new_G4632gat_ = ~new_G4512gat_ & ~new_G4578gat_;
  assign new_G4633gat_ = ~new_G4578gat_ & ~new_G4509gat_;
  assign new_G4634gat_ = ~new_G4582gat_ & ~new_G4583gat_;
  assign new_G4637gat_ = ~new_G4584gat_ & ~new_G1203gat_;
  assign new_G4641gat_ = ~new_G4521gat_ & ~new_G4587gat_;
  assign new_G4642gat_ = ~new_G4587gat_ & ~new_G1251gat_;
  assign new_G4643gat_ = ~new_G4401gat_ & ~new_G4587gat_;
  assign new_G4646gat_ = ~new_G4592gat_ & ~new_G4526gat_;
  assign new_G4650gat_ = ~new_G4595gat_ & ~new_G4531gat_;
  assign new_G4654gat_ = ~new_G4598gat_ & ~new_G4536gat_;
  assign new_G4658gat_ = ~new_G4601gat_ & ~new_G4541gat_;
  assign new_G4662gat_ = ~new_G4604gat_ & ~new_G4546gat_;
  assign new_G4666gat_ = ~new_G4554gat_ & ~new_G4607gat_;
  assign new_G4667gat_ = ~new_G4607gat_ & ~new_G4551gat_;
  assign new_G4668gat_ = ~new_G4611gat_ & ~new_G4612gat_;
  assign new_G4671gat_ = ~new_G4613gat_ & ~new_G912gat_;
  assign new_G4675gat_ = ~new_G4563gat_ & ~new_G4616gat_;
  assign new_G4676gat_ = ~new_G4616gat_ & ~new_G960gat_;
  assign new_G4677gat_ = ~new_G4435gat_ & ~new_G4616gat_;
  assign new_G4680gat_ = ~new_G4620gat_ & ~new_G4621gat_;
  assign new_G4683gat_ = ~new_G4625gat_ & ~new_G4622gat_;
  assign new_G4687gat_ = ~new_G4575gat_ & ~new_G4628gat_;
  assign new_G4688gat_ = ~new_G4628gat_ & ~new_G4572gat_;
  assign new_G4689gat_ = ~new_G4632gat_ & ~new_G4633gat_;
  assign new_G4692gat_ = ~new_G4634gat_ & ~new_G1155gat_;
  assign new_G4696gat_ = ~new_G4584gat_ & ~new_G4637gat_;
  assign new_G4697gat_ = ~new_G4637gat_ & ~new_G1203gat_;
  assign new_G4698gat_ = ~new_G4456gat_ & ~new_G4637gat_;
  assign new_G4701gat_ = ~new_G4641gat_ & ~new_G4642gat_;
  assign new_G4704gat_ = ~new_G1299gat_ & ~new_G4643gat_;
  assign new_G4708gat_ = ~new_G4592gat_ & ~new_G4646gat_;
  assign new_G4709gat_ = ~new_G4646gat_ & ~new_G4526gat_;
  assign new_G4710gat_ = ~new_G4595gat_ & ~new_G4650gat_;
  assign new_G4711gat_ = ~new_G4650gat_ & ~new_G4531gat_;
  assign new_G4712gat_ = ~new_G4598gat_ & ~new_G4654gat_;
  assign new_G4713gat_ = ~new_G4654gat_ & ~new_G4536gat_;
  assign new_G4714gat_ = ~new_G4601gat_ & ~new_G4658gat_;
  assign new_G4715gat_ = ~new_G4658gat_ & ~new_G4541gat_;
  assign new_G4716gat_ = ~new_G4604gat_ & ~new_G4662gat_;
  assign new_G4717gat_ = ~new_G4662gat_ & ~new_G4546gat_;
  assign new_G4718gat_ = ~new_G4666gat_ & ~new_G4667gat_;
  assign new_G4721gat_ = ~new_G4668gat_ & ~new_G864gat_;
  assign new_G4725gat_ = ~new_G4613gat_ & ~new_G4671gat_;
  assign new_G4726gat_ = ~new_G4671gat_ & ~new_G912gat_;
  assign new_G4727gat_ = ~new_G4494gat_ & ~new_G4671gat_;
  assign new_G4730gat_ = ~new_G4675gat_ & ~new_G4676gat_;
  assign new_G4733gat_ = ~new_G4680gat_ & ~new_G4677gat_;
  assign new_G4737gat_ = ~new_G4625gat_ & ~new_G4683gat_;
  assign new_G4738gat_ = ~new_G4683gat_ & ~new_G4622gat_;
  assign new_G4739gat_ = ~new_G4687gat_ & ~new_G4688gat_;
  assign new_G4742gat_ = ~new_G4689gat_ & ~new_G1107gat_;
  assign new_G4746gat_ = ~new_G4634gat_ & ~new_G4692gat_;
  assign new_G4747gat_ = ~new_G4692gat_ & ~new_G1155gat_;
  assign new_G4748gat_ = ~new_G4515gat_ & ~new_G4692gat_;
  assign new_G4751gat_ = ~new_G4696gat_ & ~new_G4697gat_;
  assign new_G4754gat_ = ~new_G4701gat_ & ~new_G4698gat_;
  assign new_G4758gat_ = ~new_G1299gat_ & ~new_G4704gat_;
  assign new_G4759gat_ = ~new_G4704gat_ & ~new_G4643gat_;
  assign new_G4760gat_ = ~new_G4708gat_ & ~new_G4709gat_;
  assign new_G4763gat_ = ~new_G4710gat_ & ~new_G4711gat_;
  assign new_G4766gat_ = ~new_G4712gat_ & ~new_G4713gat_;
  assign new_G4769gat_ = ~new_G4714gat_ & ~new_G4715gat_;
  assign new_G4772gat_ = ~new_G4716gat_ & ~new_G4717gat_;
  assign new_G4775gat_ = ~new_G4718gat_ & ~new_G816gat_;
  assign new_G4779gat_ = ~new_G4668gat_ & ~new_G4721gat_;
  assign new_G4780gat_ = ~new_G4721gat_ & ~new_G864gat_;
  assign new_G4781gat_ = ~new_G4557gat_ & ~new_G4721gat_;
  assign new_G4784gat_ = ~new_G4725gat_ & ~new_G4726gat_;
  assign new_G4787gat_ = ~new_G4730gat_ & ~new_G4727gat_;
  assign new_G4791gat_ = ~new_G4680gat_ & ~new_G4733gat_;
  assign new_G4792gat_ = ~new_G4733gat_ & ~new_G4677gat_;
  assign new_G4793gat_ = ~new_G4737gat_ & ~new_G4738gat_;
  assign new_G4796gat_ = ~new_G4739gat_ & ~new_G1059gat_;
  assign new_G4800gat_ = ~new_G4689gat_ & ~new_G4742gat_;
  assign new_G4801gat_ = ~new_G4742gat_ & ~new_G1107gat_;
  assign new_G4802gat_ = ~new_G4578gat_ & ~new_G4742gat_;
  assign new_G4805gat_ = ~new_G4746gat_ & ~new_G4747gat_;
  assign new_G4808gat_ = ~new_G4751gat_ & ~new_G4748gat_;
  assign new_G4812gat_ = ~new_G4701gat_ & ~new_G4754gat_;
  assign new_G4813gat_ = ~new_G4754gat_ & ~new_G4698gat_;
  assign new_G4814gat_ = ~new_G4758gat_ & ~new_G4759gat_;
  assign new_G4817gat_ = ~new_G4760gat_ & ~new_G576gat_;
  assign new_G4821gat_ = ~new_G4763gat_ & ~new_G624gat_;
  assign new_G4825gat_ = ~new_G4766gat_ & ~new_G672gat_;
  assign new_G4829gat_ = ~new_G4769gat_ & ~new_G720gat_;
  assign new_G4833gat_ = ~new_G4772gat_ & ~new_G768gat_;
  assign new_G4837gat_ = ~new_G4718gat_ & ~new_G4775gat_;
  assign new_G4838gat_ = ~new_G4775gat_ & ~new_G816gat_;
  assign new_G4839gat_ = ~new_G4607gat_ & ~new_G4775gat_;
  assign new_G4842gat_ = ~new_G4779gat_ & ~new_G4780gat_;
  assign new_G4845gat_ = ~new_G4784gat_ & ~new_G4781gat_;
  assign new_G4849gat_ = ~new_G4730gat_ & ~new_G4787gat_;
  assign new_G4850gat_ = ~new_G4787gat_ & ~new_G4727gat_;
  assign new_G4851gat_ = ~new_G4791gat_ & ~new_G4792gat_;
  assign new_G4854gat_ = ~new_G4793gat_ & ~new_G1011gat_;
  assign new_G4858gat_ = ~new_G4739gat_ & ~new_G4796gat_;
  assign new_G4859gat_ = ~new_G4796gat_ & ~new_G1059gat_;
  assign new_G4860gat_ = ~new_G4628gat_ & ~new_G4796gat_;
  assign new_G4863gat_ = ~new_G4800gat_ & ~new_G4801gat_;
  assign new_G4866gat_ = ~new_G4805gat_ & ~new_G4802gat_;
  assign new_G4870gat_ = ~new_G4751gat_ & ~new_G4808gat_;
  assign new_G4871gat_ = ~new_G4808gat_ & ~new_G4748gat_;
  assign new_G4872gat_ = ~new_G4812gat_ & ~new_G4813gat_;
  assign new_G4875gat_ = ~new_G4814gat_ & ~new_G1254gat_;
  assign new_G4879gat_ = ~new_G4760gat_ & ~new_G4817gat_;
  assign new_G4880gat_ = ~new_G4817gat_ & ~new_G576gat_;
  assign new_G4881gat_ = ~new_G4646gat_ & ~new_G4817gat_;
  assign new_G4884gat_ = ~new_G4763gat_ & ~new_G4821gat_;
  assign new_G4885gat_ = ~new_G4821gat_ & ~new_G624gat_;
  assign new_G4886gat_ = ~new_G4650gat_ & ~new_G4821gat_;
  assign new_G4889gat_ = ~new_G4766gat_ & ~new_G4825gat_;
  assign new_G4890gat_ = ~new_G4825gat_ & ~new_G672gat_;
  assign new_G4891gat_ = ~new_G4654gat_ & ~new_G4825gat_;
  assign new_G4894gat_ = ~new_G4769gat_ & ~new_G4829gat_;
  assign new_G4895gat_ = ~new_G4829gat_ & ~new_G720gat_;
  assign new_G4896gat_ = ~new_G4658gat_ & ~new_G4829gat_;
  assign new_G4899gat_ = ~new_G4772gat_ & ~new_G4833gat_;
  assign new_G4900gat_ = ~new_G4833gat_ & ~new_G768gat_;
  assign new_G4901gat_ = ~new_G4662gat_ & ~new_G4833gat_;
  assign new_G4904gat_ = ~new_G4837gat_ & ~new_G4838gat_;
  assign new_G4907gat_ = ~new_G4842gat_ & ~new_G4839gat_;
  assign new_G4911gat_ = ~new_G4784gat_ & ~new_G4845gat_;
  assign new_G4912gat_ = ~new_G4845gat_ & ~new_G4781gat_;
  assign new_G4913gat_ = ~new_G4849gat_ & ~new_G4850gat_;
  assign new_G4916gat_ = ~new_G4851gat_ & ~new_G963gat_;
  assign new_G4920gat_ = ~new_G4793gat_ & ~new_G4854gat_;
  assign new_G4921gat_ = ~new_G4854gat_ & ~new_G1011gat_;
  assign new_G4922gat_ = ~new_G4683gat_ & ~new_G4854gat_;
  assign new_G4925gat_ = ~new_G4858gat_ & ~new_G4859gat_;
  assign new_G4928gat_ = ~new_G4863gat_ & ~new_G4860gat_;
  assign new_G4932gat_ = ~new_G4805gat_ & ~new_G4866gat_;
  assign new_G4933gat_ = ~new_G4866gat_ & ~new_G4802gat_;
  assign new_G4934gat_ = ~new_G4870gat_ & ~new_G4871gat_;
  assign new_G4937gat_ = ~new_G4872gat_ & ~new_G1206gat_;
  assign new_G4941gat_ = ~new_G4814gat_ & ~new_G4875gat_;
  assign new_G4942gat_ = ~new_G4875gat_ & ~new_G1254gat_;
  assign new_G4943gat_ = ~new_G4704gat_ & ~new_G4875gat_;
  assign G4946gat = ~new_G4879gat_ & ~new_G4880gat_;
  assign new_G4947gat_ = ~new_G4884gat_ & ~new_G4885gat_;
  assign new_G4950gat_ = ~new_G4889gat_ & ~new_G4890gat_;
  assign new_G4953gat_ = ~new_G4894gat_ & ~new_G4895gat_;
  assign new_G4956gat_ = ~new_G4899gat_ & ~new_G4900gat_;
  assign new_G4959gat_ = ~new_G4904gat_ & ~new_G4901gat_;
  assign new_G4963gat_ = ~new_G4842gat_ & ~new_G4907gat_;
  assign new_G4964gat_ = ~new_G4907gat_ & ~new_G4839gat_;
  assign new_G4965gat_ = ~new_G4911gat_ & ~new_G4912gat_;
  assign new_G4968gat_ = ~new_G4913gat_ & ~new_G915gat_;
  assign new_G4972gat_ = ~new_G4851gat_ & ~new_G4916gat_;
  assign new_G4973gat_ = ~new_G4916gat_ & ~new_G963gat_;
  assign new_G4974gat_ = ~new_G4733gat_ & ~new_G4916gat_;
  assign new_G4977gat_ = ~new_G4920gat_ & ~new_G4921gat_;
  assign new_G4980gat_ = ~new_G4925gat_ & ~new_G4922gat_;
  assign new_G4984gat_ = ~new_G4863gat_ & ~new_G4928gat_;
  assign new_G4985gat_ = ~new_G4928gat_ & ~new_G4860gat_;
  assign new_G4986gat_ = ~new_G4932gat_ & ~new_G4933gat_;
  assign new_G4989gat_ = ~new_G4934gat_ & ~new_G1158gat_;
  assign new_G4993gat_ = ~new_G4872gat_ & ~new_G4937gat_;
  assign new_G4994gat_ = ~new_G4937gat_ & ~new_G1206gat_;
  assign new_G4995gat_ = ~new_G4754gat_ & ~new_G4937gat_;
  assign new_G4998gat_ = ~new_G4941gat_ & ~new_G4942gat_;
  assign new_G5001gat_ = ~new_G1302gat_ & ~new_G4943gat_;
  assign new_G5005gat_ = ~new_G4947gat_ & ~new_G4881gat_;
  assign new_G5009gat_ = ~new_G4950gat_ & ~new_G4886gat_;
  assign new_G5013gat_ = ~new_G4953gat_ & ~new_G4891gat_;
  assign new_G5017gat_ = ~new_G4956gat_ & ~new_G4896gat_;
  assign new_G5021gat_ = ~new_G4904gat_ & ~new_G4959gat_;
  assign new_G5022gat_ = ~new_G4959gat_ & ~new_G4901gat_;
  assign new_G5023gat_ = ~new_G4963gat_ & ~new_G4964gat_;
  assign new_G5026gat_ = ~new_G4965gat_ & ~new_G867gat_;
  assign new_G5030gat_ = ~new_G4913gat_ & ~new_G4968gat_;
  assign new_G5031gat_ = ~new_G4968gat_ & ~new_G915gat_;
  assign new_G5032gat_ = ~new_G4787gat_ & ~new_G4968gat_;
  assign new_G5035gat_ = ~new_G4972gat_ & ~new_G4973gat_;
  assign new_G5038gat_ = ~new_G4977gat_ & ~new_G4974gat_;
  assign new_G5042gat_ = ~new_G4925gat_ & ~new_G4980gat_;
  assign new_G5043gat_ = ~new_G4980gat_ & ~new_G4922gat_;
  assign new_G5044gat_ = ~new_G4984gat_ & ~new_G4985gat_;
  assign new_G5047gat_ = ~new_G4986gat_ & ~new_G1110gat_;
  assign new_G5051gat_ = ~new_G4934gat_ & ~new_G4989gat_;
  assign new_G5052gat_ = ~new_G4989gat_ & ~new_G1158gat_;
  assign new_G5053gat_ = ~new_G4808gat_ & ~new_G4989gat_;
  assign new_G5056gat_ = ~new_G4993gat_ & ~new_G4994gat_;
  assign new_G5059gat_ = ~new_G4998gat_ & ~new_G4995gat_;
  assign new_G5063gat_ = ~new_G1302gat_ & ~new_G5001gat_;
  assign new_G5064gat_ = ~new_G5001gat_ & ~new_G4943gat_;
  assign new_G5065gat_ = ~new_G4947gat_ & ~new_G5005gat_;
  assign new_G5066gat_ = ~new_G5005gat_ & ~new_G4881gat_;
  assign new_G5067gat_ = ~new_G4950gat_ & ~new_G5009gat_;
  assign new_G5068gat_ = ~new_G5009gat_ & ~new_G4886gat_;
  assign new_G5069gat_ = ~new_G4953gat_ & ~new_G5013gat_;
  assign new_G5070gat_ = ~new_G5013gat_ & ~new_G4891gat_;
  assign new_G5071gat_ = ~new_G4956gat_ & ~new_G5017gat_;
  assign new_G5072gat_ = ~new_G5017gat_ & ~new_G4896gat_;
  assign new_G5073gat_ = ~new_G5021gat_ & ~new_G5022gat_;
  assign new_G5076gat_ = ~new_G5023gat_ & ~new_G819gat_;
  assign new_G5080gat_ = ~new_G4965gat_ & ~new_G5026gat_;
  assign new_G5081gat_ = ~new_G5026gat_ & ~new_G867gat_;
  assign new_G5082gat_ = ~new_G4845gat_ & ~new_G5026gat_;
  assign new_G5085gat_ = ~new_G5030gat_ & ~new_G5031gat_;
  assign new_G5088gat_ = ~new_G5035gat_ & ~new_G5032gat_;
  assign new_G5092gat_ = ~new_G4977gat_ & ~new_G5038gat_;
  assign new_G5093gat_ = ~new_G5038gat_ & ~new_G4974gat_;
  assign new_G5094gat_ = ~new_G5042gat_ & ~new_G5043gat_;
  assign new_G5097gat_ = ~new_G5044gat_ & ~new_G1062gat_;
  assign new_G5101gat_ = ~new_G4986gat_ & ~new_G5047gat_;
  assign new_G5102gat_ = ~new_G5047gat_ & ~new_G1110gat_;
  assign new_G5103gat_ = ~new_G4866gat_ & ~new_G5047gat_;
  assign new_G5106gat_ = ~new_G5051gat_ & ~new_G5052gat_;
  assign new_G5109gat_ = ~new_G5056gat_ & ~new_G5053gat_;
  assign new_G5113gat_ = ~new_G4998gat_ & ~new_G5059gat_;
  assign new_G5114gat_ = ~new_G5059gat_ & ~new_G4995gat_;
  assign new_G5115gat_ = ~new_G5063gat_ & ~new_G5064gat_;
  assign new_G5118gat_ = ~new_G5065gat_ & ~new_G5066gat_;
  assign new_G5121gat_ = ~new_G5067gat_ & ~new_G5068gat_;
  assign new_G5124gat_ = ~new_G5069gat_ & ~new_G5070gat_;
  assign new_G5127gat_ = ~new_G5071gat_ & ~new_G5072gat_;
  assign new_G5130gat_ = ~new_G5073gat_ & ~new_G771gat_;
  assign new_G5134gat_ = ~new_G5023gat_ & ~new_G5076gat_;
  assign new_G5135gat_ = ~new_G5076gat_ & ~new_G819gat_;
  assign new_G5136gat_ = ~new_G4907gat_ & ~new_G5076gat_;
  assign new_G5139gat_ = ~new_G5080gat_ & ~new_G5081gat_;
  assign new_G5142gat_ = ~new_G5085gat_ & ~new_G5082gat_;
  assign new_G5146gat_ = ~new_G5035gat_ & ~new_G5088gat_;
  assign new_G5147gat_ = ~new_G5088gat_ & ~new_G5032gat_;
  assign new_G5148gat_ = ~new_G5092gat_ & ~new_G5093gat_;
  assign new_G5151gat_ = ~new_G5094gat_ & ~new_G1014gat_;
  assign new_G5155gat_ = ~new_G5044gat_ & ~new_G5097gat_;
  assign new_G5156gat_ = ~new_G5097gat_ & ~new_G1062gat_;
  assign new_G5157gat_ = ~new_G4928gat_ & ~new_G5097gat_;
  assign new_G5160gat_ = ~new_G5101gat_ & ~new_G5102gat_;
  assign new_G5163gat_ = ~new_G5106gat_ & ~new_G5103gat_;
  assign new_G5167gat_ = ~new_G5056gat_ & ~new_G5109gat_;
  assign new_G5168gat_ = ~new_G5109gat_ & ~new_G5053gat_;
  assign new_G5169gat_ = ~new_G5113gat_ & ~new_G5114gat_;
  assign new_G5172gat_ = ~new_G5115gat_ & ~new_G1257gat_;
  assign new_G5176gat_ = ~new_G5118gat_ & ~new_G579gat_;
  assign new_G5180gat_ = ~new_G5121gat_ & ~new_G627gat_;
  assign new_G5184gat_ = ~new_G5124gat_ & ~new_G675gat_;
  assign new_G5188gat_ = ~new_G5127gat_ & ~new_G723gat_;
  assign new_G5192gat_ = ~new_G5073gat_ & ~new_G5130gat_;
  assign new_G5193gat_ = ~new_G5130gat_ & ~new_G771gat_;
  assign new_G5194gat_ = ~new_G4959gat_ & ~new_G5130gat_;
  assign new_G5197gat_ = ~new_G5134gat_ & ~new_G5135gat_;
  assign new_G5200gat_ = ~new_G5139gat_ & ~new_G5136gat_;
  assign new_G5204gat_ = ~new_G5085gat_ & ~new_G5142gat_;
  assign new_G5205gat_ = ~new_G5142gat_ & ~new_G5082gat_;
  assign new_G5206gat_ = ~new_G5146gat_ & ~new_G5147gat_;
  assign new_G5209gat_ = ~new_G5148gat_ & ~new_G966gat_;
  assign new_G5213gat_ = ~new_G5094gat_ & ~new_G5151gat_;
  assign new_G5214gat_ = ~new_G5151gat_ & ~new_G1014gat_;
  assign new_G5215gat_ = ~new_G4980gat_ & ~new_G5151gat_;
  assign new_G5218gat_ = ~new_G5155gat_ & ~new_G5156gat_;
  assign new_G5221gat_ = ~new_G5160gat_ & ~new_G5157gat_;
  assign new_G5225gat_ = ~new_G5106gat_ & ~new_G5163gat_;
  assign new_G5226gat_ = ~new_G5163gat_ & ~new_G5103gat_;
  assign new_G5227gat_ = ~new_G5167gat_ & ~new_G5168gat_;
  assign new_G5230gat_ = ~new_G5169gat_ & ~new_G1209gat_;
  assign new_G5234gat_ = ~new_G5115gat_ & ~new_G5172gat_;
  assign new_G5235gat_ = ~new_G5172gat_ & ~new_G1257gat_;
  assign new_G5236gat_ = ~new_G5001gat_ & ~new_G5172gat_;
  assign new_G5239gat_ = ~new_G5118gat_ & ~new_G5176gat_;
  assign new_G5240gat_ = ~new_G5176gat_ & ~new_G579gat_;
  assign new_G5241gat_ = ~new_G5005gat_ & ~new_G5176gat_;
  assign new_G5244gat_ = ~new_G5121gat_ & ~new_G5180gat_;
  assign new_G5245gat_ = ~new_G5180gat_ & ~new_G627gat_;
  assign new_G5246gat_ = ~new_G5009gat_ & ~new_G5180gat_;
  assign new_G5249gat_ = ~new_G5124gat_ & ~new_G5184gat_;
  assign new_G5250gat_ = ~new_G5184gat_ & ~new_G675gat_;
  assign new_G5251gat_ = ~new_G5013gat_ & ~new_G5184gat_;
  assign new_G5254gat_ = ~new_G5127gat_ & ~new_G5188gat_;
  assign new_G5255gat_ = ~new_G5188gat_ & ~new_G723gat_;
  assign new_G5256gat_ = ~new_G5017gat_ & ~new_G5188gat_;
  assign new_G5259gat_ = ~new_G5192gat_ & ~new_G5193gat_;
  assign new_G5262gat_ = ~new_G5197gat_ & ~new_G5194gat_;
  assign new_G5266gat_ = ~new_G5139gat_ & ~new_G5200gat_;
  assign new_G5267gat_ = ~new_G5200gat_ & ~new_G5136gat_;
  assign new_G5268gat_ = ~new_G5204gat_ & ~new_G5205gat_;
  assign new_G5271gat_ = ~new_G5206gat_ & ~new_G918gat_;
  assign new_G5275gat_ = ~new_G5148gat_ & ~new_G5209gat_;
  assign new_G5276gat_ = ~new_G5209gat_ & ~new_G966gat_;
  assign new_G5277gat_ = ~new_G5038gat_ & ~new_G5209gat_;
  assign new_G5280gat_ = ~new_G5213gat_ & ~new_G5214gat_;
  assign new_G5283gat_ = ~new_G5218gat_ & ~new_G5215gat_;
  assign new_G5287gat_ = ~new_G5160gat_ & ~new_G5221gat_;
  assign new_G5288gat_ = ~new_G5221gat_ & ~new_G5157gat_;
  assign new_G5289gat_ = ~new_G5225gat_ & ~new_G5226gat_;
  assign new_G5292gat_ = ~new_G5227gat_ & ~new_G1161gat_;
  assign new_G5296gat_ = ~new_G5169gat_ & ~new_G5230gat_;
  assign new_G5297gat_ = ~new_G5230gat_ & ~new_G1209gat_;
  assign new_G5298gat_ = ~new_G5059gat_ & ~new_G5230gat_;
  assign new_G5301gat_ = ~new_G5234gat_ & ~new_G5235gat_;
  assign new_G5304gat_ = ~new_G1305gat_ & ~new_G5236gat_;
  assign G5308gat = ~new_G5239gat_ & ~new_G5240gat_;
  assign new_G5309gat_ = ~new_G5244gat_ & ~new_G5245gat_;
  assign new_G5312gat_ = ~new_G5249gat_ & ~new_G5250gat_;
  assign new_G5315gat_ = ~new_G5254gat_ & ~new_G5255gat_;
  assign new_G5318gat_ = ~new_G5259gat_ & ~new_G5256gat_;
  assign new_G5322gat_ = ~new_G5197gat_ & ~new_G5262gat_;
  assign new_G5323gat_ = ~new_G5262gat_ & ~new_G5194gat_;
  assign new_G5324gat_ = ~new_G5266gat_ & ~new_G5267gat_;
  assign new_G5327gat_ = ~new_G5268gat_ & ~new_G870gat_;
  assign new_G5331gat_ = ~new_G5206gat_ & ~new_G5271gat_;
  assign new_G5332gat_ = ~new_G5271gat_ & ~new_G918gat_;
  assign new_G5333gat_ = ~new_G5088gat_ & ~new_G5271gat_;
  assign new_G5336gat_ = ~new_G5275gat_ & ~new_G5276gat_;
  assign new_G5339gat_ = ~new_G5280gat_ & ~new_G5277gat_;
  assign new_G5343gat_ = ~new_G5218gat_ & ~new_G5283gat_;
  assign new_G5344gat_ = ~new_G5283gat_ & ~new_G5215gat_;
  assign new_G5345gat_ = ~new_G5287gat_ & ~new_G5288gat_;
  assign new_G5348gat_ = ~new_G5289gat_ & ~new_G1113gat_;
  assign new_G5352gat_ = ~new_G5227gat_ & ~new_G5292gat_;
  assign new_G5353gat_ = ~new_G5292gat_ & ~new_G1161gat_;
  assign new_G5354gat_ = ~new_G5109gat_ & ~new_G5292gat_;
  assign new_G5357gat_ = ~new_G5296gat_ & ~new_G5297gat_;
  assign new_G5360gat_ = ~new_G5301gat_ & ~new_G5298gat_;
  assign new_G5364gat_ = ~new_G1305gat_ & ~new_G5304gat_;
  assign new_G5365gat_ = ~new_G5304gat_ & ~new_G5236gat_;
  assign new_G5366gat_ = ~new_G5309gat_ & ~new_G5241gat_;
  assign new_G5370gat_ = ~new_G5312gat_ & ~new_G5246gat_;
  assign new_G5374gat_ = ~new_G5315gat_ & ~new_G5251gat_;
  assign new_G5378gat_ = ~new_G5259gat_ & ~new_G5318gat_;
  assign new_G5379gat_ = ~new_G5318gat_ & ~new_G5256gat_;
  assign new_G5380gat_ = ~new_G5322gat_ & ~new_G5323gat_;
  assign new_G5383gat_ = ~new_G5324gat_ & ~new_G822gat_;
  assign new_G5387gat_ = ~new_G5268gat_ & ~new_G5327gat_;
  assign new_G5388gat_ = ~new_G5327gat_ & ~new_G870gat_;
  assign new_G5389gat_ = ~new_G5142gat_ & ~new_G5327gat_;
  assign new_G5392gat_ = ~new_G5331gat_ & ~new_G5332gat_;
  assign new_G5395gat_ = ~new_G5336gat_ & ~new_G5333gat_;
  assign new_G5399gat_ = ~new_G5280gat_ & ~new_G5339gat_;
  assign new_G5400gat_ = ~new_G5339gat_ & ~new_G5277gat_;
  assign new_G5401gat_ = ~new_G5343gat_ & ~new_G5344gat_;
  assign new_G5404gat_ = ~new_G5345gat_ & ~new_G1065gat_;
  assign new_G5408gat_ = ~new_G5289gat_ & ~new_G5348gat_;
  assign new_G5409gat_ = ~new_G5348gat_ & ~new_G1113gat_;
  assign new_G5410gat_ = ~new_G5163gat_ & ~new_G5348gat_;
  assign new_G5413gat_ = ~new_G5352gat_ & ~new_G5353gat_;
  assign new_G5416gat_ = ~new_G5357gat_ & ~new_G5354gat_;
  assign new_G5420gat_ = ~new_G5301gat_ & ~new_G5360gat_;
  assign new_G5421gat_ = ~new_G5360gat_ & ~new_G5298gat_;
  assign new_G5422gat_ = ~new_G5364gat_ & ~new_G5365gat_;
  assign new_G5425gat_ = ~new_G5309gat_ & ~new_G5366gat_;
  assign new_G5426gat_ = ~new_G5366gat_ & ~new_G5241gat_;
  assign new_G5427gat_ = ~new_G5312gat_ & ~new_G5370gat_;
  assign new_G5428gat_ = ~new_G5370gat_ & ~new_G5246gat_;
  assign new_G5429gat_ = ~new_G5315gat_ & ~new_G5374gat_;
  assign new_G5430gat_ = ~new_G5374gat_ & ~new_G5251gat_;
  assign new_G5431gat_ = ~new_G5378gat_ & ~new_G5379gat_;
  assign new_G5434gat_ = ~new_G5380gat_ & ~new_G774gat_;
  assign new_G5438gat_ = ~new_G5324gat_ & ~new_G5383gat_;
  assign new_G5439gat_ = ~new_G5383gat_ & ~new_G822gat_;
  assign new_G5440gat_ = ~new_G5200gat_ & ~new_G5383gat_;
  assign new_G5443gat_ = ~new_G5387gat_ & ~new_G5388gat_;
  assign new_G5446gat_ = ~new_G5392gat_ & ~new_G5389gat_;
  assign new_G5450gat_ = ~new_G5336gat_ & ~new_G5395gat_;
  assign new_G5451gat_ = ~new_G5395gat_ & ~new_G5333gat_;
  assign new_G5452gat_ = ~new_G5399gat_ & ~new_G5400gat_;
  assign new_G5455gat_ = ~new_G5401gat_ & ~new_G1017gat_;
  assign new_G5459gat_ = ~new_G5345gat_ & ~new_G5404gat_;
  assign new_G5460gat_ = ~new_G5404gat_ & ~new_G1065gat_;
  assign new_G5461gat_ = ~new_G5221gat_ & ~new_G5404gat_;
  assign new_G5464gat_ = ~new_G5408gat_ & ~new_G5409gat_;
  assign new_G5467gat_ = ~new_G5413gat_ & ~new_G5410gat_;
  assign new_G5471gat_ = ~new_G5357gat_ & ~new_G5416gat_;
  assign new_G5472gat_ = ~new_G5416gat_ & ~new_G5354gat_;
  assign new_G5473gat_ = ~new_G5420gat_ & ~new_G5421gat_;
  assign new_G5476gat_ = ~new_G5422gat_ & ~new_G1260gat_;
  assign new_G5480gat_ = ~new_G5425gat_ & ~new_G5426gat_;
  assign new_G5483gat_ = ~new_G5427gat_ & ~new_G5428gat_;
  assign new_G5486gat_ = ~new_G5429gat_ & ~new_G5430gat_;
  assign new_G5489gat_ = ~new_G5431gat_ & ~new_G726gat_;
  assign new_G5493gat_ = ~new_G5380gat_ & ~new_G5434gat_;
  assign new_G5494gat_ = ~new_G5434gat_ & ~new_G774gat_;
  assign new_G5495gat_ = ~new_G5262gat_ & ~new_G5434gat_;
  assign new_G5498gat_ = ~new_G5438gat_ & ~new_G5439gat_;
  assign new_G5501gat_ = ~new_G5443gat_ & ~new_G5440gat_;
  assign new_G5505gat_ = ~new_G5392gat_ & ~new_G5446gat_;
  assign new_G5506gat_ = ~new_G5446gat_ & ~new_G5389gat_;
  assign new_G5507gat_ = ~new_G5450gat_ & ~new_G5451gat_;
  assign new_G5510gat_ = ~new_G5452gat_ & ~new_G969gat_;
  assign new_G5514gat_ = ~new_G5401gat_ & ~new_G5455gat_;
  assign new_G5515gat_ = ~new_G5455gat_ & ~new_G1017gat_;
  assign new_G5516gat_ = ~new_G5283gat_ & ~new_G5455gat_;
  assign new_G5519gat_ = ~new_G5459gat_ & ~new_G5460gat_;
  assign new_G5522gat_ = ~new_G5464gat_ & ~new_G5461gat_;
  assign new_G5526gat_ = ~new_G5413gat_ & ~new_G5467gat_;
  assign new_G5527gat_ = ~new_G5467gat_ & ~new_G5410gat_;
  assign new_G5528gat_ = ~new_G5471gat_ & ~new_G5472gat_;
  assign new_G5531gat_ = ~new_G5473gat_ & ~new_G1212gat_;
  assign new_G5535gat_ = ~new_G5422gat_ & ~new_G5476gat_;
  assign new_G5536gat_ = ~new_G5476gat_ & ~new_G1260gat_;
  assign new_G5537gat_ = ~new_G5304gat_ & ~new_G5476gat_;
  assign new_G5540gat_ = ~new_G5480gat_ & ~new_G582gat_;
  assign new_G5544gat_ = ~new_G5483gat_ & ~new_G630gat_;
  assign new_G5548gat_ = ~new_G5486gat_ & ~new_G678gat_;
  assign new_G5552gat_ = ~new_G5431gat_ & ~new_G5489gat_;
  assign new_G5553gat_ = ~new_G5489gat_ & ~new_G726gat_;
  assign new_G5554gat_ = ~new_G5318gat_ & ~new_G5489gat_;
  assign new_G5557gat_ = ~new_G5493gat_ & ~new_G5494gat_;
  assign new_G5560gat_ = ~new_G5498gat_ & ~new_G5495gat_;
  assign new_G5564gat_ = ~new_G5443gat_ & ~new_G5501gat_;
  assign new_G5565gat_ = ~new_G5501gat_ & ~new_G5440gat_;
  assign new_G5566gat_ = ~new_G5505gat_ & ~new_G5506gat_;
  assign new_G5569gat_ = ~new_G5507gat_ & ~new_G921gat_;
  assign new_G5573gat_ = ~new_G5452gat_ & ~new_G5510gat_;
  assign new_G5574gat_ = ~new_G5510gat_ & ~new_G969gat_;
  assign new_G5575gat_ = ~new_G5339gat_ & ~new_G5510gat_;
  assign new_G5578gat_ = ~new_G5514gat_ & ~new_G5515gat_;
  assign new_G5581gat_ = ~new_G5519gat_ & ~new_G5516gat_;
  assign new_G5585gat_ = ~new_G5464gat_ & ~new_G5522gat_;
  assign new_G5586gat_ = ~new_G5522gat_ & ~new_G5461gat_;
  assign new_G5587gat_ = ~new_G5526gat_ & ~new_G5527gat_;
  assign new_G5590gat_ = ~new_G5528gat_ & ~new_G1164gat_;
  assign new_G5594gat_ = ~new_G5473gat_ & ~new_G5531gat_;
  assign new_G5595gat_ = ~new_G5531gat_ & ~new_G1212gat_;
  assign new_G5596gat_ = ~new_G5360gat_ & ~new_G5531gat_;
  assign new_G5599gat_ = ~new_G5535gat_ & ~new_G5536gat_;
  assign new_G5602gat_ = ~new_G1308gat_ & ~new_G5537gat_;
  assign new_G5606gat_ = ~new_G5480gat_ & ~new_G5540gat_;
  assign new_G5607gat_ = ~new_G5540gat_ & ~new_G582gat_;
  assign new_G5608gat_ = ~new_G5366gat_ & ~new_G5540gat_;
  assign new_G5611gat_ = ~new_G5483gat_ & ~new_G5544gat_;
  assign new_G5612gat_ = ~new_G5544gat_ & ~new_G630gat_;
  assign new_G5613gat_ = ~new_G5370gat_ & ~new_G5544gat_;
  assign new_G5616gat_ = ~new_G5486gat_ & ~new_G5548gat_;
  assign new_G5617gat_ = ~new_G5548gat_ & ~new_G678gat_;
  assign new_G5618gat_ = ~new_G5374gat_ & ~new_G5548gat_;
  assign new_G5621gat_ = ~new_G5552gat_ & ~new_G5553gat_;
  assign new_G5624gat_ = ~new_G5557gat_ & ~new_G5554gat_;
  assign new_G5628gat_ = ~new_G5498gat_ & ~new_G5560gat_;
  assign new_G5629gat_ = ~new_G5560gat_ & ~new_G5495gat_;
  assign new_G5630gat_ = ~new_G5564gat_ & ~new_G5565gat_;
  assign new_G5633gat_ = ~new_G5566gat_ & ~new_G873gat_;
  assign new_G5637gat_ = ~new_G5507gat_ & ~new_G5569gat_;
  assign new_G5638gat_ = ~new_G5569gat_ & ~new_G921gat_;
  assign new_G5639gat_ = ~new_G5395gat_ & ~new_G5569gat_;
  assign new_G5642gat_ = ~new_G5573gat_ & ~new_G5574gat_;
  assign new_G5645gat_ = ~new_G5578gat_ & ~new_G5575gat_;
  assign new_G5649gat_ = ~new_G5519gat_ & ~new_G5581gat_;
  assign new_G5650gat_ = ~new_G5581gat_ & ~new_G5516gat_;
  assign new_G5651gat_ = ~new_G5585gat_ & ~new_G5586gat_;
  assign new_G5654gat_ = ~new_G5587gat_ & ~new_G1116gat_;
  assign new_G5658gat_ = ~new_G5528gat_ & ~new_G5590gat_;
  assign new_G5659gat_ = ~new_G5590gat_ & ~new_G1164gat_;
  assign new_G5660gat_ = ~new_G5416gat_ & ~new_G5590gat_;
  assign new_G5663gat_ = ~new_G5594gat_ & ~new_G5595gat_;
  assign new_G5666gat_ = ~new_G5599gat_ & ~new_G5596gat_;
  assign new_G5670gat_ = ~new_G1308gat_ & ~new_G5602gat_;
  assign new_G5671gat_ = ~new_G5602gat_ & ~new_G5537gat_;
  assign G5672gat = ~new_G5606gat_ & ~new_G5607gat_;
  assign new_G5673gat_ = ~new_G5611gat_ & ~new_G5612gat_;
  assign new_G5676gat_ = ~new_G5616gat_ & ~new_G5617gat_;
  assign new_G5679gat_ = ~new_G5621gat_ & ~new_G5618gat_;
  assign new_G5683gat_ = ~new_G5557gat_ & ~new_G5624gat_;
  assign new_G5684gat_ = ~new_G5624gat_ & ~new_G5554gat_;
  assign new_G5685gat_ = ~new_G5628gat_ & ~new_G5629gat_;
  assign new_G5688gat_ = ~new_G5630gat_ & ~new_G825gat_;
  assign new_G5692gat_ = ~new_G5566gat_ & ~new_G5633gat_;
  assign new_G5693gat_ = ~new_G5633gat_ & ~new_G873gat_;
  assign new_G5694gat_ = ~new_G5446gat_ & ~new_G5633gat_;
  assign new_G5697gat_ = ~new_G5637gat_ & ~new_G5638gat_;
  assign new_G5700gat_ = ~new_G5642gat_ & ~new_G5639gat_;
  assign new_G5704gat_ = ~new_G5578gat_ & ~new_G5645gat_;
  assign new_G5705gat_ = ~new_G5645gat_ & ~new_G5575gat_;
  assign new_G5706gat_ = ~new_G5649gat_ & ~new_G5650gat_;
  assign new_G5709gat_ = ~new_G5651gat_ & ~new_G1068gat_;
  assign new_G5713gat_ = ~new_G5587gat_ & ~new_G5654gat_;
  assign new_G5714gat_ = ~new_G5654gat_ & ~new_G1116gat_;
  assign new_G5715gat_ = ~new_G5467gat_ & ~new_G5654gat_;
  assign new_G5718gat_ = ~new_G5658gat_ & ~new_G5659gat_;
  assign new_G5721gat_ = ~new_G5663gat_ & ~new_G5660gat_;
  assign new_G5725gat_ = ~new_G5599gat_ & ~new_G5666gat_;
  assign new_G5726gat_ = ~new_G5666gat_ & ~new_G5596gat_;
  assign new_G5727gat_ = ~new_G5670gat_ & ~new_G5671gat_;
  assign new_G5730gat_ = ~new_G5673gat_ & ~new_G5608gat_;
  assign new_G5734gat_ = ~new_G5676gat_ & ~new_G5613gat_;
  assign new_G5738gat_ = ~new_G5621gat_ & ~new_G5679gat_;
  assign new_G5739gat_ = ~new_G5679gat_ & ~new_G5618gat_;
  assign new_G5740gat_ = ~new_G5683gat_ & ~new_G5684gat_;
  assign new_G5743gat_ = ~new_G5685gat_ & ~new_G777gat_;
  assign new_G5747gat_ = ~new_G5630gat_ & ~new_G5688gat_;
  assign new_G5748gat_ = ~new_G5688gat_ & ~new_G825gat_;
  assign new_G5749gat_ = ~new_G5501gat_ & ~new_G5688gat_;
  assign new_G5752gat_ = ~new_G5692gat_ & ~new_G5693gat_;
  assign new_G5755gat_ = ~new_G5697gat_ & ~new_G5694gat_;
  assign new_G5759gat_ = ~new_G5642gat_ & ~new_G5700gat_;
  assign new_G5760gat_ = ~new_G5700gat_ & ~new_G5639gat_;
  assign new_G5761gat_ = ~new_G5704gat_ & ~new_G5705gat_;
  assign new_G5764gat_ = ~new_G5706gat_ & ~new_G1020gat_;
  assign new_G5768gat_ = ~new_G5651gat_ & ~new_G5709gat_;
  assign new_G5769gat_ = ~new_G5709gat_ & ~new_G1068gat_;
  assign new_G5770gat_ = ~new_G5522gat_ & ~new_G5709gat_;
  assign new_G5773gat_ = ~new_G5713gat_ & ~new_G5714gat_;
  assign new_G5776gat_ = ~new_G5718gat_ & ~new_G5715gat_;
  assign new_G5780gat_ = ~new_G5663gat_ & ~new_G5721gat_;
  assign new_G5781gat_ = ~new_G5721gat_ & ~new_G5660gat_;
  assign new_G5782gat_ = ~new_G5725gat_ & ~new_G5726gat_;
  assign new_G5785gat_ = ~new_G5673gat_ & ~new_G5730gat_;
  assign new_G5786gat_ = ~new_G5730gat_ & ~new_G5608gat_;
  assign new_G5787gat_ = ~new_G5676gat_ & ~new_G5734gat_;
  assign new_G5788gat_ = ~new_G5734gat_ & ~new_G5613gat_;
  assign new_G5789gat_ = ~new_G5738gat_ & ~new_G5739gat_;
  assign new_G5792gat_ = ~new_G5740gat_ & ~new_G729gat_;
  assign new_G5796gat_ = ~new_G5685gat_ & ~new_G5743gat_;
  assign new_G5797gat_ = ~new_G5743gat_ & ~new_G777gat_;
  assign new_G5798gat_ = ~new_G5560gat_ & ~new_G5743gat_;
  assign new_G5801gat_ = ~new_G5747gat_ & ~new_G5748gat_;
  assign new_G5804gat_ = ~new_G5752gat_ & ~new_G5749gat_;
  assign new_G5808gat_ = ~new_G5697gat_ & ~new_G5755gat_;
  assign new_G5809gat_ = ~new_G5755gat_ & ~new_G5694gat_;
  assign new_G5810gat_ = ~new_G5759gat_ & ~new_G5760gat_;
  assign new_G5813gat_ = ~new_G5761gat_ & ~new_G972gat_;
  assign new_G5817gat_ = ~new_G5706gat_ & ~new_G5764gat_;
  assign new_G5818gat_ = ~new_G5764gat_ & ~new_G1020gat_;
  assign new_G5819gat_ = ~new_G5581gat_ & ~new_G5764gat_;
  assign new_G5822gat_ = ~new_G5768gat_ & ~new_G5769gat_;
  assign new_G5825gat_ = ~new_G5773gat_ & ~new_G5770gat_;
  assign new_G5829gat_ = ~new_G5718gat_ & ~new_G5776gat_;
  assign new_G5830gat_ = ~new_G5776gat_ & ~new_G5715gat_;
  assign new_G5831gat_ = ~new_G5780gat_ & ~new_G5781gat_;
  assign new_G5834gat_ = ~new_G5785gat_ & ~new_G5786gat_;
  assign new_G5837gat_ = ~new_G5787gat_ & ~new_G5788gat_;
  assign new_G5840gat_ = ~new_G5789gat_ & ~new_G681gat_;
  assign new_G5844gat_ = ~new_G5740gat_ & ~new_G5792gat_;
  assign new_G5845gat_ = ~new_G5792gat_ & ~new_G729gat_;
  assign new_G5846gat_ = ~new_G5624gat_ & ~new_G5792gat_;
  assign new_G5849gat_ = ~new_G5796gat_ & ~new_G5797gat_;
  assign new_G5852gat_ = ~new_G5801gat_ & ~new_G5798gat_;
  assign new_G5856gat_ = ~new_G5752gat_ & ~new_G5804gat_;
  assign new_G5857gat_ = ~new_G5804gat_ & ~new_G5749gat_;
  assign new_G5858gat_ = ~new_G5808gat_ & ~new_G5809gat_;
  assign new_G5861gat_ = ~new_G5810gat_ & ~new_G924gat_;
  assign new_G5865gat_ = ~new_G5761gat_ & ~new_G5813gat_;
  assign new_G5866gat_ = ~new_G5813gat_ & ~new_G972gat_;
  assign new_G5867gat_ = ~new_G5645gat_ & ~new_G5813gat_;
  assign new_G5870gat_ = ~new_G5817gat_ & ~new_G5818gat_;
  assign new_G5873gat_ = ~new_G5822gat_ & ~new_G5819gat_;
  assign new_G5877gat_ = ~new_G5773gat_ & ~new_G5825gat_;
  assign new_G5878gat_ = ~new_G5825gat_ & ~new_G5770gat_;
  assign new_G5879gat_ = ~new_G5829gat_ & ~new_G5830gat_;
  assign new_G5882gat_ = ~new_G5834gat_ & ~new_G585gat_;
  assign new_G5886gat_ = ~new_G5837gat_ & ~new_G633gat_;
  assign new_G5890gat_ = ~new_G5789gat_ & ~new_G5840gat_;
  assign new_G5891gat_ = ~new_G5840gat_ & ~new_G681gat_;
  assign new_G5892gat_ = ~new_G5679gat_ & ~new_G5840gat_;
  assign new_G5895gat_ = ~new_G5844gat_ & ~new_G5845gat_;
  assign new_G5898gat_ = ~new_G5849gat_ & ~new_G5846gat_;
  assign new_G5902gat_ = ~new_G5801gat_ & ~new_G5852gat_;
  assign new_G5903gat_ = ~new_G5852gat_ & ~new_G5798gat_;
  assign new_G5904gat_ = ~new_G5856gat_ & ~new_G5857gat_;
  assign new_G5907gat_ = ~new_G5858gat_ & ~new_G876gat_;
  assign new_G5911gat_ = ~new_G5810gat_ & ~new_G5861gat_;
  assign new_G5912gat_ = ~new_G5861gat_ & ~new_G924gat_;
  assign new_G5913gat_ = ~new_G5700gat_ & ~new_G5861gat_;
  assign new_G5916gat_ = ~new_G5865gat_ & ~new_G5866gat_;
  assign new_G5919gat_ = ~new_G5870gat_ & ~new_G5867gat_;
  assign new_G5923gat_ = ~new_G5822gat_ & ~new_G5873gat_;
  assign new_G5924gat_ = ~new_G5873gat_ & ~new_G5819gat_;
  assign new_G5925gat_ = ~new_G5877gat_ & ~new_G5878gat_;
  assign new_G5928gat_ = ~new_G5834gat_ & ~new_G5882gat_;
  assign new_G5929gat_ = ~new_G5882gat_ & ~new_G585gat_;
  assign new_G5930gat_ = ~new_G5730gat_ & ~new_G5882gat_;
  assign new_G5933gat_ = ~new_G5837gat_ & ~new_G5886gat_;
  assign new_G5934gat_ = ~new_G5886gat_ & ~new_G633gat_;
  assign new_G5935gat_ = ~new_G5734gat_ & ~new_G5886gat_;
  assign new_G5938gat_ = ~new_G5890gat_ & ~new_G5891gat_;
  assign new_G5941gat_ = ~new_G5895gat_ & ~new_G5892gat_;
  assign new_G5945gat_ = ~new_G5849gat_ & ~new_G5898gat_;
  assign new_G5946gat_ = ~new_G5898gat_ & ~new_G5846gat_;
  assign new_G5947gat_ = ~new_G5902gat_ & ~new_G5903gat_;
  assign new_G5950gat_ = ~new_G5904gat_ & ~new_G828gat_;
  assign new_G5954gat_ = ~new_G5858gat_ & ~new_G5907gat_;
  assign new_G5955gat_ = ~new_G5907gat_ & ~new_G876gat_;
  assign new_G5956gat_ = ~new_G5755gat_ & ~new_G5907gat_;
  assign new_G5959gat_ = ~new_G5911gat_ & ~new_G5912gat_;
  assign new_G5962gat_ = ~new_G5916gat_ & ~new_G5913gat_;
  assign new_G5966gat_ = ~new_G5870gat_ & ~new_G5919gat_;
  assign new_G5967gat_ = ~new_G5919gat_ & ~new_G5867gat_;
  assign new_G5968gat_ = ~new_G5923gat_ & ~new_G5924gat_;
  assign G5971gat = ~new_G5928gat_ & ~new_G5929gat_;
  assign new_G5972gat_ = ~new_G5933gat_ & ~new_G5934gat_;
  assign new_G5975gat_ = ~new_G5938gat_ & ~new_G5935gat_;
  assign new_G5979gat_ = ~new_G5895gat_ & ~new_G5941gat_;
  assign new_G5980gat_ = ~new_G5941gat_ & ~new_G5892gat_;
  assign new_G5981gat_ = ~new_G5945gat_ & ~new_G5946gat_;
  assign new_G5984gat_ = ~new_G5947gat_ & ~new_G780gat_;
  assign new_G5988gat_ = ~new_G5904gat_ & ~new_G5950gat_;
  assign new_G5989gat_ = ~new_G5950gat_ & ~new_G828gat_;
  assign new_G5990gat_ = ~new_G5804gat_ & ~new_G5950gat_;
  assign new_G5993gat_ = ~new_G5954gat_ & ~new_G5955gat_;
  assign new_G5996gat_ = ~new_G5959gat_ & ~new_G5956gat_;
  assign new_G6000gat_ = ~new_G5916gat_ & ~new_G5962gat_;
  assign new_G6001gat_ = ~new_G5962gat_ & ~new_G5913gat_;
  assign new_G6002gat_ = ~new_G5966gat_ & ~new_G5967gat_;
  assign new_G6005gat_ = ~new_G5972gat_ & ~new_G5930gat_;
  assign new_G6009gat_ = ~new_G5938gat_ & ~new_G5975gat_;
  assign new_G6010gat_ = ~new_G5975gat_ & ~new_G5935gat_;
  assign new_G6011gat_ = ~new_G5979gat_ & ~new_G5980gat_;
  assign new_G6014gat_ = ~new_G5981gat_ & ~new_G732gat_;
  assign new_G6018gat_ = ~new_G5947gat_ & ~new_G5984gat_;
  assign new_G6019gat_ = ~new_G5984gat_ & ~new_G780gat_;
  assign new_G6020gat_ = ~new_G5852gat_ & ~new_G5984gat_;
  assign new_G6023gat_ = ~new_G5988gat_ & ~new_G5989gat_;
  assign new_G6026gat_ = ~new_G5993gat_ & ~new_G5990gat_;
  assign new_G6030gat_ = ~new_G5959gat_ & ~new_G5996gat_;
  assign new_G6031gat_ = ~new_G5996gat_ & ~new_G5956gat_;
  assign new_G6032gat_ = ~new_G6000gat_ & ~new_G6001gat_;
  assign new_G6035gat_ = ~new_G5972gat_ & ~new_G6005gat_;
  assign new_G6036gat_ = ~new_G6005gat_ & ~new_G5930gat_;
  assign new_G6037gat_ = ~new_G6009gat_ & ~new_G6010gat_;
  assign new_G6040gat_ = ~new_G6011gat_ & ~new_G684gat_;
  assign new_G6044gat_ = ~new_G5981gat_ & ~new_G6014gat_;
  assign new_G6045gat_ = ~new_G6014gat_ & ~new_G732gat_;
  assign new_G6046gat_ = ~new_G5898gat_ & ~new_G6014gat_;
  assign new_G6049gat_ = ~new_G6018gat_ & ~new_G6019gat_;
  assign new_G6052gat_ = ~new_G6023gat_ & ~new_G6020gat_;
  assign new_G6056gat_ = ~new_G5993gat_ & ~new_G6026gat_;
  assign new_G6057gat_ = ~new_G6026gat_ & ~new_G5990gat_;
  assign new_G6058gat_ = ~new_G6030gat_ & ~new_G6031gat_;
  assign new_G6061gat_ = ~new_G6035gat_ & ~new_G6036gat_;
  assign new_G6064gat_ = ~new_G6037gat_ & ~new_G636gat_;
  assign new_G6068gat_ = ~new_G6011gat_ & ~new_G6040gat_;
  assign new_G6069gat_ = ~new_G6040gat_ & ~new_G684gat_;
  assign new_G6070gat_ = ~new_G5941gat_ & ~new_G6040gat_;
  assign new_G6073gat_ = ~new_G6044gat_ & ~new_G6045gat_;
  assign new_G6076gat_ = ~new_G6049gat_ & ~new_G6046gat_;
  assign new_G6080gat_ = ~new_G6023gat_ & ~new_G6052gat_;
  assign new_G6081gat_ = ~new_G6052gat_ & ~new_G6020gat_;
  assign new_G6082gat_ = ~new_G6056gat_ & ~new_G6057gat_;
  assign new_G6085gat_ = ~new_G6061gat_ & ~new_G588gat_;
  assign new_G6089gat_ = ~new_G6037gat_ & ~new_G6064gat_;
  assign new_G6090gat_ = ~new_G6064gat_ & ~new_G636gat_;
  assign new_G6091gat_ = ~new_G5975gat_ & ~new_G6064gat_;
  assign new_G6094gat_ = ~new_G6068gat_ & ~new_G6069gat_;
  assign new_G6097gat_ = ~new_G6073gat_ & ~new_G6070gat_;
  assign new_G6101gat_ = ~new_G6049gat_ & ~new_G6076gat_;
  assign new_G6102gat_ = ~new_G6076gat_ & ~new_G6046gat_;
  assign new_G6103gat_ = ~new_G6080gat_ & ~new_G6081gat_;
  assign new_G6106gat_ = ~new_G6061gat_ & ~new_G6085gat_;
  assign new_G6107gat_ = ~new_G6085gat_ & ~new_G588gat_;
  assign new_G6108gat_ = ~new_G6005gat_ & ~new_G6085gat_;
  assign new_G6111gat_ = ~new_G6089gat_ & ~new_G6090gat_;
  assign new_G6114gat_ = ~new_G6094gat_ & ~new_G6091gat_;
  assign new_G6118gat_ = ~new_G6073gat_ & ~new_G6097gat_;
  assign new_G6119gat_ = ~new_G6097gat_ & ~new_G6070gat_;
  assign new_G6120gat_ = ~new_G6101gat_ & ~new_G6102gat_;
  assign G6123gat = ~new_G6106gat_ & ~new_G6107gat_;
  assign new_G6124gat_ = ~new_G6111gat_ & ~new_G6108gat_;
  assign new_G6128gat_ = ~new_G6094gat_ & ~new_G6114gat_;
  assign new_G6129gat_ = ~new_G6114gat_ & ~new_G6091gat_;
  assign new_G6130gat_ = ~new_G6118gat_ & ~new_G6119gat_;
  assign new_G6133gat_ = ~new_G6111gat_ & ~new_G6124gat_;
  assign new_G6134gat_ = ~new_G6124gat_ & ~new_G6108gat_;
  assign new_G6135gat_ = ~new_G6128gat_ & ~new_G6129gat_;
  assign new_G6138gat_ = ~new_G6133gat_ & ~new_G6134gat_;
  assign new_G6141gat_ = ~new_G6138gat_;
  assign new_G6145gat_ = ~new_G6138gat_ & ~new_G6141gat_;
  assign new_G6146gat_ = ~new_G6141gat_;
  assign new_G6147gat_ = ~new_G6124gat_ & ~new_G6141gat_;
  assign G6150gat = ~new_G6145gat_ & ~new_G6146gat_;
  assign new_G6151gat_ = ~new_G6135gat_ & ~new_G6147gat_;
  assign new_G6155gat_ = ~new_G6135gat_ & ~new_G6151gat_;
  assign new_G6156gat_ = ~new_G6151gat_ & ~new_G6147gat_;
  assign new_G6157gat_ = ~new_G6114gat_ & ~new_G6151gat_;
  assign G6160gat = ~new_G6155gat_ & ~new_G6156gat_;
  assign new_G6161gat_ = ~new_G6130gat_ & ~new_G6157gat_;
  assign new_G6165gat_ = ~new_G6130gat_ & ~new_G6161gat_;
  assign new_G6166gat_ = ~new_G6161gat_ & ~new_G6157gat_;
  assign new_G6167gat_ = ~new_G6097gat_ & ~new_G6161gat_;
  assign G6170gat = ~new_G6165gat_ & ~new_G6166gat_;
  assign new_G6171gat_ = ~new_G6120gat_ & ~new_G6167gat_;
  assign new_G6175gat_ = ~new_G6120gat_ & ~new_G6171gat_;
  assign new_G6176gat_ = ~new_G6171gat_ & ~new_G6167gat_;
  assign new_G6177gat_ = ~new_G6076gat_ & ~new_G6171gat_;
  assign G6180gat = ~new_G6175gat_ & ~new_G6176gat_;
  assign new_G6181gat_ = ~new_G6103gat_ & ~new_G6177gat_;
  assign new_G6185gat_ = ~new_G6103gat_ & ~new_G6181gat_;
  assign new_G6186gat_ = ~new_G6181gat_ & ~new_G6177gat_;
  assign new_G6187gat_ = ~new_G6052gat_ & ~new_G6181gat_;
  assign G6190gat = ~new_G6185gat_ & ~new_G6186gat_;
  assign new_G6191gat_ = ~new_G6082gat_ & ~new_G6187gat_;
  assign new_G6195gat_ = ~new_G6082gat_ & ~new_G6191gat_;
  assign new_G6196gat_ = ~new_G6191gat_ & ~new_G6187gat_;
  assign new_G6197gat_ = ~new_G6026gat_ & ~new_G6191gat_;
  assign G6200gat = ~new_G6195gat_ & ~new_G6196gat_;
  assign new_G6201gat_ = ~new_G6058gat_ & ~new_G6197gat_;
  assign new_G6205gat_ = ~new_G6058gat_ & ~new_G6201gat_;
  assign new_G6206gat_ = ~new_G6201gat_ & ~new_G6197gat_;
  assign new_G6207gat_ = ~new_G5996gat_ & ~new_G6201gat_;
  assign G6210gat = ~new_G6205gat_ & ~new_G6206gat_;
  assign new_G6211gat_ = ~new_G6032gat_ & ~new_G6207gat_;
  assign new_G6215gat_ = ~new_G6032gat_ & ~new_G6211gat_;
  assign new_G6216gat_ = ~new_G6211gat_ & ~new_G6207gat_;
  assign new_G6217gat_ = ~new_G5962gat_ & ~new_G6211gat_;
  assign G6220gat = ~new_G6215gat_ & ~new_G6216gat_;
  assign new_G6221gat_ = ~new_G6002gat_ & ~new_G6217gat_;
  assign new_G6225gat_ = ~new_G6002gat_ & ~new_G6221gat_;
  assign new_G6226gat_ = ~new_G6221gat_ & ~new_G6217gat_;
  assign new_G6227gat_ = ~new_G5919gat_ & ~new_G6221gat_;
  assign G6230gat = ~new_G6225gat_ & ~new_G6226gat_;
  assign new_G6231gat_ = ~new_G5968gat_ & ~new_G6227gat_;
  assign new_G6235gat_ = ~new_G5968gat_ & ~new_G6231gat_;
  assign new_G6236gat_ = ~new_G6231gat_ & ~new_G6227gat_;
  assign new_G6237gat_ = ~new_G5873gat_ & ~new_G6231gat_;
  assign G6240gat = ~new_G6235gat_ & ~new_G6236gat_;
  assign new_G6241gat_ = ~new_G5925gat_ & ~new_G6237gat_;
  assign new_G6245gat_ = ~new_G5925gat_ & ~new_G6241gat_;
  assign new_G6246gat_ = ~new_G6241gat_ & ~new_G6237gat_;
  assign new_G6247gat_ = ~new_G5825gat_ & ~new_G6241gat_;
  assign G6250gat = ~new_G6245gat_ & ~new_G6246gat_;
  assign new_G6251gat_ = ~new_G5879gat_ & ~new_G6247gat_;
  assign new_G6255gat_ = ~new_G5879gat_ & ~new_G6251gat_;
  assign new_G6256gat_ = ~new_G6251gat_ & ~new_G6247gat_;
  assign new_G6257gat_ = ~new_G5776gat_ & ~new_G6251gat_;
  assign G6260gat = ~new_G6255gat_ & ~new_G6256gat_;
  assign new_G6261gat_ = ~new_G5831gat_ & ~new_G6257gat_;
  assign new_G6265gat_ = ~new_G5831gat_ & ~new_G6261gat_;
  assign new_G6266gat_ = ~new_G6261gat_ & ~new_G6257gat_;
  assign new_G6267gat_ = ~new_G5721gat_ & ~new_G6261gat_;
  assign G6270gat = ~new_G6265gat_ & ~new_G6266gat_;
  assign new_G6271gat_ = ~new_G5782gat_ & ~new_G6267gat_;
  assign new_G6275gat_ = ~new_G5782gat_ & ~new_G6271gat_;
  assign new_G6276gat_ = ~new_G6271gat_ & ~new_G6267gat_;
  assign new_G6277gat_ = ~new_G5666gat_ & ~new_G6271gat_;
  assign G6280gat = ~new_G6275gat_ & ~new_G6276gat_;
  assign new_G6281gat_ = ~new_G5727gat_ & ~new_G6277gat_;
  assign new_G6285gat_ = ~new_G5727gat_ & ~new_G6281gat_;
  assign new_G6286gat_ = ~new_G6281gat_ & ~new_G6277gat_;
  assign G6287gat = ~new_G5602gat_ & ~new_G6281gat_;
  assign G6288gat = ~new_G6285gat_ & ~new_G6286gat_;
endmodule


