//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT71), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT36), .ZN(new_n207_));
  INV_X1    g006(.A(G85gat), .ZN(new_n208_));
  INV_X1    g007(.A(G92gat), .ZN(new_n209_));
  NOR3_X1   g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT9), .ZN(new_n210_));
  XOR2_X1   g009(.A(G85gat), .B(G92gat), .Z(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(KEYINPUT9), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT10), .B(G99gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(G106gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT6), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n219_), .A2(KEYINPUT64), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(KEYINPUT64), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n216_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n212_), .A2(new_n214_), .A3(new_n218_), .A4(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224_));
  OAI22_X1  g023(.A1(new_n224_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(KEYINPUT66), .B2(KEYINPUT7), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OAI221_X1 g026(.A(new_n224_), .B1(KEYINPUT66), .B2(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n222_), .A2(new_n218_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n211_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n229_), .B2(new_n211_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n223_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G29gat), .B(G36gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G43gat), .B(G50gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT15), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n223_), .B(new_n236_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G232gat), .A2(G233gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT34), .Z(new_n241_));
  INV_X1    g040(.A(KEYINPUT35), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT70), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n238_), .A2(new_n239_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT69), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n241_), .A2(new_n242_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n238_), .A2(new_n239_), .A3(new_n249_), .A4(new_n245_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n248_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n207_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n250_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n248_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n205_), .B(KEYINPUT36), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n251_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT72), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n254_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT37), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n257_), .A2(KEYINPUT72), .A3(new_n251_), .A4(new_n258_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n254_), .A2(new_n259_), .A3(KEYINPUT37), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT75), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G127gat), .B(G155gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT16), .ZN(new_n269_));
  XOR2_X1   g068(.A(G183gat), .B(G211gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT17), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n267_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G57gat), .B(G64gat), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT11), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT11), .ZN(new_n276_));
  XOR2_X1   g075(.A(G71gat), .B(G78gat), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n276_), .A2(new_n277_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n273_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G1gat), .B(G8gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT73), .ZN(new_n284_));
  INV_X1    g083(.A(G15gat), .ZN(new_n285_));
  INV_X1    g084(.A(G22gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G15gat), .A2(G22gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G1gat), .A2(G8gat), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n287_), .A2(new_n288_), .B1(KEYINPUT14), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n284_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n282_), .B(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G231gat), .A2(G233gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT74), .Z(new_n294_));
  OR2_X1    g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n294_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n271_), .A2(new_n272_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n266_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n233_), .A2(new_n281_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n280_), .B(new_n223_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G230gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT12), .B1(new_n233_), .B2(new_n281_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n305_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G176gat), .B(G204gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT68), .ZN(new_n311_));
  XOR2_X1   g110(.A(G120gat), .B(G148gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  OR3_X1    g115(.A1(new_n308_), .A2(new_n309_), .A3(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n317_), .A2(KEYINPUT13), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT13), .B1(new_n317_), .B2(new_n318_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n300_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT94), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G1gat), .B(G29gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G85gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT0), .B(G57gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT1), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT83), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G155gat), .ZN(new_n340_));
  INV_X1    g139(.A(G162gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(KEYINPUT82), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT82), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(G155gat), .B2(G162gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(G155gat), .A3(G162gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n333_), .B1(new_n339_), .B2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n342_), .A2(new_n344_), .A3(new_n334_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351_));
  INV_X1    g150(.A(G141gat), .ZN(new_n352_));
  INV_X1    g151(.A(G148gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT2), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n330_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .A4(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n350_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n348_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G127gat), .B(G134gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G113gat), .B(G120gat), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n363_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n348_), .A2(new_n372_), .A3(new_n360_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n364_), .A2(new_n366_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n364_), .A2(new_n366_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n376_), .A2(new_n348_), .A3(new_n372_), .A4(new_n360_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n371_), .B1(new_n378_), .B2(KEYINPUT4), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n370_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n329_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n369_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n365_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n382_), .B(new_n328_), .C1(new_n383_), .C2(new_n371_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n324_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n381_), .A2(new_n324_), .A3(new_n384_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G169gat), .ZN(new_n389_));
  INV_X1    g188(.A(G176gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(KEYINPUT24), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(G183gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT76), .B1(new_n394_), .B2(KEYINPUT25), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT25), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(G183gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(KEYINPUT25), .ZN(new_n400_));
  INV_X1    g199(.A(G190gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT26), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT26), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(G190gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n393_), .B1(new_n399_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT77), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT77), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n408_), .B(new_n393_), .C1(new_n399_), .C2(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G183gat), .A2(G190gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT23), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n412_), .B(new_n413_), .C1(new_n391_), .C2(KEYINPUT24), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(new_n409_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT22), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n418_));
  OAI21_X1  g217(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n412_), .A2(new_n413_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n394_), .A2(new_n401_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n416_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G71gat), .B(G99gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT79), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n428_), .A2(KEYINPUT79), .ZN(new_n431_));
  OAI21_X1  g230(.A(G15gat), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n428_), .A2(KEYINPUT79), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(new_n429_), .A3(new_n285_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G227gat), .A2(G233gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n436_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n432_), .A2(new_n438_), .A3(new_n434_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n414_), .B1(new_n406_), .B2(KEYINPUT77), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n423_), .B1(new_n441_), .B2(new_n409_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT30), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n427_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n432_), .A2(new_n438_), .A3(new_n434_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n438_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI211_X1 g246(.A(new_n426_), .B(new_n423_), .C1(new_n441_), .C2(new_n409_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT30), .B1(new_n416_), .B2(new_n424_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n444_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT78), .B(G43gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT80), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n374_), .B(KEYINPUT31), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(KEYINPUT81), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n444_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n454_), .A2(new_n458_), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT81), .B1(new_n460_), .B2(new_n455_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n456_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n388_), .B(new_n459_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G211gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(G218gat), .ZN(new_n465_));
  INV_X1    g264(.A(G218gat), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(G211gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT87), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(G197gat), .A2(G204gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G197gat), .A2(G204gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(KEYINPUT21), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT21), .ZN(new_n473_));
  INV_X1    g272(.A(new_n471_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n473_), .B1(new_n474_), .B2(new_n469_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n466_), .A2(G211gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n464_), .A2(G218gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n468_), .A2(new_n472_), .A3(new_n475_), .A4(new_n479_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n474_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n478_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n416_), .B2(new_n424_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G226gat), .A2(G233gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n420_), .A2(KEYINPUT90), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n412_), .A2(new_n422_), .A3(new_n413_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n418_), .A2(new_n493_), .A3(new_n419_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT24), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT89), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT24), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n391_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n397_), .A2(G183gat), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n400_), .A2(new_n402_), .A3(new_n404_), .A4(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n391_), .A2(new_n497_), .A3(new_n499_), .A4(new_n392_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n502_), .A2(new_n421_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n495_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n480_), .A2(new_n484_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT20), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n486_), .A2(new_n490_), .A3(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n416_), .A2(new_n424_), .A3(new_n485_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT20), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n489_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G8gat), .B(G36gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G64gat), .B(G92gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n510_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n490_), .B1(new_n486_), .B2(new_n509_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n511_), .A2(new_n489_), .A3(new_n513_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT27), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n520_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n519_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n511_), .A2(new_n513_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n490_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n495_), .A2(new_n506_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n512_), .B1(new_n531_), .B2(new_n485_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n532_), .B(new_n489_), .C1(new_n442_), .C2(new_n485_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n530_), .A2(new_n521_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n528_), .A2(new_n534_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n526_), .A2(new_n527_), .B1(new_n525_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n334_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT83), .B1(new_n334_), .B2(KEYINPUT1), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n342_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n542_), .A2(new_n333_), .B1(new_n359_), .B2(new_n350_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT29), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n537_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n333_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n354_), .A2(new_n358_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n356_), .A2(new_n357_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n349_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NOR4_X1   g349(.A1(new_n547_), .A2(new_n550_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT84), .B1(new_n545_), .B2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT28), .B1(new_n361_), .B2(KEYINPUT29), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n543_), .A2(new_n537_), .A3(new_n544_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT84), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n544_), .B1(new_n348_), .B2(new_n360_), .ZN(new_n557_));
  OAI21_X1  g356(.A(G78gat), .B1(new_n557_), .B2(new_n485_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT29), .B1(new_n547_), .B2(new_n550_), .ZN(new_n559_));
  INV_X1    g358(.A(G78gat), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n508_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n558_), .A2(new_n561_), .A3(G106gat), .ZN(new_n562_));
  AOI21_X1  g361(.A(G106gat), .B1(new_n558_), .B2(new_n561_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n552_), .B(new_n556_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n552_), .A2(new_n556_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n558_), .A2(new_n561_), .ZN(new_n566_));
  INV_X1    g365(.A(G106gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n558_), .A2(new_n561_), .A3(G106gat), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n565_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(KEYINPUT85), .A2(G228gat), .ZN(new_n571_));
  NOR2_X1   g370(.A1(KEYINPUT85), .A2(G228gat), .ZN(new_n572_));
  OAI21_X1  g371(.A(G233gat), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT86), .Z(new_n574_));
  XNOR2_X1  g373(.A(G22gat), .B(G50gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  AND3_X1   g375(.A1(new_n564_), .A2(new_n570_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n564_), .B2(new_n570_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n534_), .A2(KEYINPUT27), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT95), .B1(new_n580_), .B2(new_n524_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n536_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT96), .B1(new_n463_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n535_), .A2(new_n525_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n524_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n585_), .A2(new_n527_), .A3(KEYINPUT27), .A4(new_n534_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n581_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n564_), .A2(new_n570_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n576_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n564_), .A2(new_n570_), .A3(new_n576_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n594_));
  INV_X1    g393(.A(new_n459_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n444_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n452_), .B1(new_n444_), .B2(new_n450_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n455_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT81), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n595_), .B1(new_n600_), .B2(new_n456_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n593_), .A2(new_n594_), .A3(new_n601_), .A4(new_n388_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n378_), .A2(KEYINPUT4), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n369_), .A3(new_n368_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n328_), .B1(new_n378_), .B2(new_n370_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT93), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT93), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n604_), .A2(new_n608_), .A3(new_n605_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n535_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n384_), .B(KEYINPUT33), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n381_), .A2(new_n384_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n521_), .A2(KEYINPUT32), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n510_), .A2(new_n514_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n615_), .B2(new_n613_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n610_), .A2(new_n611_), .B1(new_n612_), .B2(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n381_), .A2(new_n324_), .A3(new_n384_), .ZN(new_n618_));
  OAI22_X1  g417(.A1(new_n577_), .A2(new_n578_), .B1(new_n618_), .B2(new_n385_), .ZN(new_n619_));
  OAI22_X1  g418(.A1(new_n617_), .A2(new_n592_), .B1(new_n619_), .B2(new_n587_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n601_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n583_), .A2(new_n602_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n291_), .B(new_n236_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n291_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n237_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n291_), .A2(new_n236_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n624_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G169gat), .B(G197gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n632_), .B(new_n633_), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n631_), .B(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n622_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n323_), .A2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n637_), .A2(G1gat), .A3(new_n388_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n261_), .A2(new_n263_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n622_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n321_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n643_), .A2(new_n299_), .A3(new_n635_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n618_), .A2(new_n385_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n649_), .A2(KEYINPUT99), .A3(G1gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT99), .B1(new_n649_), .B2(G1gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n640_), .B1(new_n650_), .B2(new_n651_), .ZN(G1324gat));
  INV_X1    g451(.A(new_n587_), .ZN(new_n653_));
  OR3_X1    g452(.A1(new_n637_), .A2(G8gat), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n642_), .A2(new_n587_), .A3(new_n644_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G8gat), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT100), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(KEYINPUT100), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n658_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n654_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g462(.A1(new_n647_), .A2(new_n601_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G15gat), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(KEYINPUT102), .A3(G15gat), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n637_), .A2(G15gat), .A3(new_n621_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .ZN(G1326gat));
  NAND2_X1  g472(.A1(new_n647_), .A2(new_n592_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G22gat), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT42), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT42), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n592_), .A2(new_n286_), .ZN(new_n678_));
  OAI22_X1  g477(.A1(new_n676_), .A2(new_n677_), .B1(new_n637_), .B2(new_n678_), .ZN(G1327gat));
  INV_X1    g478(.A(new_n641_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n643_), .A2(new_n680_), .A3(new_n298_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n620_), .A2(new_n621_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n463_), .A2(new_n582_), .A3(KEYINPUT96), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n462_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n684_), .A2(new_n648_), .A3(new_n595_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n594_), .B1(new_n685_), .B2(new_n593_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n683_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n635_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n681_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n636_), .A2(KEYINPUT104), .A3(new_n681_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n648_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n643_), .A2(new_n298_), .A3(new_n635_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n687_), .A2(new_n266_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT43), .B1(new_n696_), .B2(KEYINPUT103), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n264_), .A2(new_n265_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT103), .B(KEYINPUT43), .C1(new_n622_), .C2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n695_), .B1(new_n697_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT44), .B(new_n695_), .C1(new_n697_), .C2(new_n700_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n648_), .A2(G29gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n694_), .B1(new_n705_), .B2(new_n706_), .ZN(G1328gat));
  NOR2_X1   g506(.A1(new_n653_), .A2(G36gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n691_), .A2(new_n692_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n712_));
  NAND4_X1  g511(.A1(new_n691_), .A2(KEYINPUT106), .A3(new_n692_), .A4(new_n708_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n703_), .A2(new_n587_), .A3(new_n704_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(new_n718_), .A3(G36gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n717_), .B2(G36gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT46), .B(new_n716_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  NAND3_X1  g524(.A1(new_n705_), .A2(G43gat), .A3(new_n601_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n693_), .A2(new_n601_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n727_), .A2(G43gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(G1330gat));
  AOI21_X1  g530(.A(G50gat), .B1(new_n693_), .B2(new_n592_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n592_), .A2(G50gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n705_), .B2(new_n733_), .ZN(G1331gat));
  NOR2_X1   g533(.A1(new_n321_), .A2(new_n688_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(new_n299_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n642_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(G57gat), .A3(new_n648_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n740_), .A2(new_n741_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n736_), .A2(new_n622_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n300_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G57gat), .B1(new_n746_), .B2(new_n648_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n742_), .A2(new_n743_), .A3(new_n747_), .ZN(G1332gat));
  OR3_X1    g547(.A1(new_n745_), .A2(G64gat), .A3(new_n653_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n739_), .A2(new_n587_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G64gat), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  XOR2_X1   g552(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n753_), .A2(new_n754_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n749_), .B1(new_n755_), .B2(new_n756_), .ZN(G1333gat));
  OAI21_X1  g556(.A(G71gat), .B1(new_n738_), .B2(new_n621_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT49), .Z(new_n759_));
  NOR3_X1   g558(.A1(new_n745_), .A2(G71gat), .A3(new_n621_), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1334gat));
  OAI21_X1  g560(.A(G78gat), .B1(new_n738_), .B2(new_n579_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT50), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n746_), .A2(new_n560_), .A3(new_n592_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1335gat));
  OR2_X1    g564(.A1(new_n697_), .A2(new_n700_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n736_), .A2(new_n298_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n388_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n680_), .A2(new_n298_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n744_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n648_), .A2(new_n208_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n769_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT112), .Z(G1336gat));
  NOR3_X1   g573(.A1(new_n768_), .A2(new_n209_), .A3(new_n653_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n209_), .B1(new_n771_), .B2(new_n653_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT113), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n768_), .B2(new_n621_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n771_), .A2(new_n621_), .A3(new_n213_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT114), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g582(.A1(new_n766_), .A2(new_n592_), .A3(new_n767_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n592_), .A2(new_n567_), .ZN(new_n788_));
  OAI22_X1  g587(.A1(new_n786_), .A2(new_n787_), .B1(new_n771_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g589(.A1(new_n688_), .A2(G113gat), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT119), .Z(new_n792_));
  INV_X1    g591(.A(new_n317_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n631_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n628_), .A2(new_n629_), .A3(new_n625_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n634_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n794_), .A2(new_n634_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n793_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n223_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n229_), .A2(new_n211_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT8), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n229_), .A2(new_n230_), .A3(new_n211_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n800_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(new_n280_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n303_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT12), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n307_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n305_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT115), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n302_), .A2(new_n303_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n307_), .B1(new_n811_), .B2(KEYINPUT12), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n305_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n306_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n810_), .A2(new_n814_), .A3(KEYINPUT55), .A4(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(KEYINPUT55), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n813_), .B1(new_n812_), .B2(new_n305_), .ZN(new_n818_));
  NOR4_X1   g617(.A1(new_n304_), .A2(KEYINPUT115), .A3(new_n306_), .A4(new_n307_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n816_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n821_), .A2(KEYINPUT118), .A3(KEYINPUT56), .A4(new_n316_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n315_), .B1(new_n816_), .B2(new_n820_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(KEYINPUT56), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT118), .B1(new_n823_), .B2(KEYINPUT56), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n799_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT58), .B(new_n799_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n266_), .A3(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n680_), .A2(KEYINPUT57), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n317_), .A2(new_n318_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n798_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n793_), .A2(new_n635_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n821_), .A2(new_n316_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n823_), .A2(KEYINPUT56), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n836_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n834_), .B1(new_n841_), .B2(KEYINPUT116), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n823_), .A2(KEYINPUT56), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n838_), .B(new_n315_), .C1(new_n816_), .C2(new_n820_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT116), .B(new_n835_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n831_), .B1(new_n842_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n830_), .A2(new_n847_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n835_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n833_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n845_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n850_), .B1(new_n854_), .B2(new_n680_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n299_), .B1(new_n848_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT54), .B1(new_n322_), .B2(new_n688_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n300_), .A2(new_n858_), .A3(new_n635_), .A4(new_n321_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n861_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n621_), .A2(new_n582_), .A3(new_n388_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT59), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n641_), .B1(new_n853_), .B2(new_n845_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n830_), .B(new_n847_), .C1(new_n865_), .C2(new_n850_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n860_), .B1(new_n866_), .B2(new_n299_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  INV_X1    g667(.A(new_n863_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n792_), .B1(new_n864_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872_));
  INV_X1    g671(.A(G113gat), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n862_), .A2(new_n863_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n635_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n871_), .A2(new_n872_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n792_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n868_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n698_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n829_), .A2(new_n879_), .B1(new_n854_), .B2(new_n831_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n854_), .A2(new_n680_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n849_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n298_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(KEYINPUT59), .B(new_n863_), .C1(new_n883_), .C2(new_n860_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n877_), .B1(new_n878_), .B2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n867_), .A2(new_n869_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G113gat), .B1(new_n886_), .B2(new_n688_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT120), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n876_), .A2(new_n888_), .ZN(G1340gat));
  INV_X1    g688(.A(G120gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n321_), .B2(KEYINPUT60), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n886_), .B(new_n891_), .C1(KEYINPUT60), .C2(new_n890_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n321_), .B1(new_n878_), .B2(new_n884_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n890_), .ZN(G1341gat));
  INV_X1    g693(.A(G127gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n886_), .A2(new_n895_), .A3(new_n298_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n299_), .B1(new_n878_), .B2(new_n884_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n895_), .ZN(G1342gat));
  INV_X1    g697(.A(G134gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n886_), .A2(new_n899_), .A3(new_n641_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n698_), .B1(new_n878_), .B2(new_n884_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1343gat));
  NOR3_X1   g701(.A1(new_n601_), .A2(new_n388_), .A3(new_n579_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n862_), .A2(new_n653_), .A3(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n635_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n352_), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n321_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n353_), .ZN(G1345gat));
  NOR2_X1   g707(.A1(new_n904_), .A2(new_n299_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT61), .B(G155gat), .Z(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  NOR3_X1   g710(.A1(new_n904_), .A2(new_n341_), .A3(new_n698_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n341_), .B1(new_n904_), .B2(new_n680_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  OAI211_X1 g714(.A(KEYINPUT121), .B(new_n341_), .C1(new_n904_), .C2(new_n680_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n912_), .B1(new_n915_), .B2(new_n916_), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n463_), .A2(new_n653_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n862_), .A2(new_n579_), .A3(new_n688_), .A4(new_n918_), .ZN(new_n919_));
  XOR2_X1   g718(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n920_));
  AOI21_X1  g719(.A(new_n389_), .B1(new_n920_), .B2(KEYINPUT123), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n920_), .A2(KEYINPUT123), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n919_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT22), .B(G169gat), .Z(new_n926_));
  OAI22_X1  g725(.A1(new_n924_), .A2(new_n925_), .B1(new_n919_), .B2(new_n926_), .ZN(G1348gat));
  OAI211_X1 g726(.A(new_n579_), .B(new_n918_), .C1(new_n883_), .C2(new_n860_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(G176gat), .B1(new_n929_), .B2(new_n643_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n867_), .A2(new_n592_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(KEYINPUT124), .B1(new_n867_), .B2(new_n592_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NOR4_X1   g734(.A1(new_n321_), .A2(new_n390_), .A3(new_n653_), .A4(new_n463_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n930_), .B1(new_n935_), .B2(new_n936_), .ZN(G1349gat));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n400_), .A2(new_n503_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n298_), .A2(new_n939_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n938_), .B1(new_n928_), .B2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n940_), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n931_), .A2(KEYINPUT125), .A3(new_n918_), .A4(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n933_), .A2(new_n298_), .A3(new_n918_), .A4(new_n934_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n394_), .B2(new_n945_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n928_), .B2(new_n698_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n641_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n928_), .B2(new_n948_), .ZN(G1351gat));
  NOR3_X1   g748(.A1(new_n601_), .A2(new_n653_), .A3(new_n619_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n862_), .A2(KEYINPUT126), .A3(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952_));
  INV_X1    g751(.A(new_n950_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n867_), .B2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n951_), .A2(new_n954_), .ZN(new_n955_));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955_), .B2(new_n688_), .ZN(new_n956_));
  INV_X1    g755(.A(G197gat), .ZN(new_n957_));
  AOI211_X1 g756(.A(new_n957_), .B(new_n635_), .C1(new_n951_), .C2(new_n954_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n956_), .A2(new_n958_), .ZN(G1352gat));
  NAND2_X1  g758(.A1(new_n955_), .A2(new_n643_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(G204gat), .ZN(new_n961_));
  INV_X1    g760(.A(G204gat), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n955_), .A2(new_n962_), .A3(new_n643_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n963_), .ZN(G1353gat));
  NOR2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  INV_X1    g764(.A(new_n965_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n299_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(new_n955_), .B2(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(new_n967_), .ZN(new_n969_));
  AOI211_X1 g768(.A(new_n965_), .B(new_n969_), .C1(new_n951_), .C2(new_n954_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n968_), .A2(new_n970_), .ZN(G1354gat));
  NAND2_X1  g770(.A1(new_n955_), .A2(new_n641_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n266_), .A2(G218gat), .ZN(new_n973_));
  XOR2_X1   g772(.A(new_n973_), .B(KEYINPUT127), .Z(new_n974_));
  AOI22_X1  g773(.A1(new_n972_), .A2(new_n466_), .B1(new_n955_), .B2(new_n974_), .ZN(G1355gat));
endmodule


