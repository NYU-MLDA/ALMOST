//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_;
  OAI211_X1 g000(.A(G85gat), .B(G92gat), .C1(KEYINPUT64), .C2(KEYINPUT9), .ZN(new_n202_));
  OAI211_X1 g001(.A(KEYINPUT64), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n209_), .B1(new_n212_), .B2(G106gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT65), .B1(new_n204_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n213_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n202_), .B(new_n203_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT7), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n223_), .A2(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT68), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n232_));
  OAI22_X1  g031(.A1(new_n231_), .A2(new_n232_), .B1(G99gat), .B2(G106gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n228_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n209_), .A3(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G85gat), .B(G92gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n220_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(new_n209_), .A3(new_n228_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n237_), .A2(KEYINPUT8), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT67), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n244_), .A3(new_n241_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n219_), .B1(new_n239_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT69), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G29gat), .B(G36gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n252_), .B(new_n219_), .C1(new_n239_), .C2(new_n246_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n248_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n251_), .B(KEYINPUT15), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n247_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT34), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n254_), .B(new_n256_), .C1(KEYINPUT35), .C2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(KEYINPUT35), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G190gat), .B(G218gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G134gat), .B(G162gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT36), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n264_), .A2(KEYINPUT36), .ZN(new_n266_));
  OR3_X1    g065(.A1(new_n261_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n261_), .A2(new_n265_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT37), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n269_), .A2(KEYINPUT70), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(KEYINPUT70), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n272_), .B(KEYINPUT71), .Z(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G15gat), .B(G22gat), .ZN(new_n276_));
  INV_X1    g075(.A(G1gat), .ZN(new_n277_));
  INV_X1    g076(.A(G8gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT14), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G8gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G231gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G57gat), .B(G64gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT11), .ZN(new_n286_));
  XOR2_X1   g085(.A(G71gat), .B(G78gat), .Z(new_n287_));
  AND2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(KEYINPUT11), .B2(new_n285_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n286_), .A2(new_n287_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n284_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G155gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT16), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G183gat), .B(G211gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT17), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n295_), .B(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n299_), .A2(KEYINPUT17), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n293_), .B2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n303_), .B(KEYINPUT73), .Z(new_n304_));
  NAND4_X1  g103(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .A4(new_n273_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n275_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT74), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT19), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(G183gat), .A3(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT82), .ZN(new_n312_));
  INV_X1    g111(.A(G183gat), .ZN(new_n313_));
  INV_X1    g112(.A(G190gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT23), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n312_), .B(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G169gat), .ZN(new_n320_));
  INV_X1    g119(.A(G176gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT22), .B(G169gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n321_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n324_), .B2(KEYINPUT81), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n319_), .B(new_n325_), .C1(KEYINPUT81), .C2(new_n324_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n315_), .A2(new_n311_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n320_), .A2(new_n321_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n328_), .A2(KEYINPUT24), .ZN(new_n329_));
  INV_X1    g128(.A(new_n322_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(KEYINPUT24), .A3(new_n328_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT25), .B(G183gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G190gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n330_), .A2(KEYINPUT79), .A3(KEYINPUT24), .A4(new_n328_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n327_), .B(new_n329_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n338_), .A2(new_n339_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n326_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G211gat), .B(G218gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT85), .B(G197gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(G204gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT21), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(G197gat), .B2(G204gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G197gat), .A2(G204gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n344_), .B2(G204gat), .ZN(new_n350_));
  OAI221_X1 g149(.A(new_n343_), .B1(new_n345_), .B2(new_n348_), .C1(KEYINPUT21), .C2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n343_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(KEYINPUT21), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n342_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n327_), .A2(new_n318_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n330_), .B(KEYINPUT88), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n323_), .B(KEYINPUT89), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n356_), .B(new_n357_), .C1(new_n358_), .C2(G176gat), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n316_), .A2(new_n331_), .A3(new_n336_), .A4(new_n329_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n354_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT20), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n309_), .B1(new_n355_), .B2(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n364_), .A2(KEYINPUT90), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n342_), .A2(new_n354_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n366_), .B(KEYINPUT20), .C1(new_n354_), .C2(new_n361_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n364_), .B(KEYINPUT90), .C1(new_n367_), .C2(new_n309_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT18), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n369_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n369_), .A2(new_n373_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n355_), .A2(new_n363_), .ZN(new_n377_));
  MUX2_X1   g176(.A(new_n377_), .B(new_n367_), .S(new_n309_), .Z(new_n378_));
  INV_X1    g177(.A(new_n373_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n374_), .A2(new_n375_), .B1(new_n376_), .B2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384_));
  NOR3_X1   g183(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G141gat), .A2(G148gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT2), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n392_));
  NOR2_X1   g191(.A1(G141gat), .A2(G148gat), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n390_), .B(new_n391_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n383_), .B(new_n384_), .C1(new_n387_), .C2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n382_), .B1(KEYINPUT1), .B2(new_n384_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(KEYINPUT1), .B2(new_n384_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n393_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n388_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G127gat), .B(G134gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G113gat), .B(G120gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n397_), .A2(new_n401_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n405_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(KEYINPUT4), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n411_), .B(KEYINPUT91), .Z(new_n412_));
  OAI211_X1 g211(.A(new_n410_), .B(new_n412_), .C1(KEYINPUT4), .C2(new_n409_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n407_), .A2(new_n409_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n411_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G1gat), .B(G29gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(G57gat), .B(G85gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(KEYINPUT92), .B(KEYINPUT0), .Z(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n413_), .A2(new_n415_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G71gat), .B(G99gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G43gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n342_), .B(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n406_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(G15gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT30), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT31), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n426_), .A2(new_n406_), .ZN(new_n435_));
  OR3_X1    g234(.A1(new_n428_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n434_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n354_), .B1(new_n402_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n354_), .ZN(new_n441_));
  OAI211_X1 g240(.A(G228gat), .B(G233gat), .C1(new_n441_), .C2(KEYINPUT86), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G78gat), .B(G106gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n354_), .B(new_n442_), .C1(new_n402_), .C2(new_n439_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n444_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G22gat), .B(G50gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT28), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n402_), .A2(new_n452_), .A3(new_n439_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT28), .B1(new_n408_), .B2(KEYINPUT29), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n451_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n454_), .A3(new_n451_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT87), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n450_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT87), .ZN(new_n460_));
  INV_X1    g259(.A(new_n457_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(new_n461_), .B2(new_n455_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n456_), .A2(KEYINPUT87), .A3(new_n457_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n462_), .B(new_n463_), .C1(new_n449_), .C2(new_n448_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n438_), .A2(new_n459_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n438_), .B1(new_n464_), .B2(new_n459_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n381_), .B(new_n423_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n459_), .A2(new_n464_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n469_), .A2(new_n438_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT32), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n369_), .B1(new_n471_), .B2(new_n379_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n378_), .A2(KEYINPUT32), .A3(new_n373_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n472_), .B(new_n473_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n413_), .A2(KEYINPUT33), .A3(new_n415_), .A4(new_n420_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n420_), .B1(new_n414_), .B2(new_n412_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n410_), .B(new_n411_), .C1(KEYINPUT4), .C2(new_n409_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n475_), .B1(new_n421_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n474_), .B1(new_n480_), .B2(new_n374_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n470_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n468_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G230gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n248_), .A2(new_n291_), .A3(new_n253_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n291_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n485_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n247_), .A2(KEYINPUT12), .A3(new_n292_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n486_), .B(new_n490_), .C1(new_n488_), .C2(KEYINPUT12), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(new_n491_), .B2(new_n485_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G120gat), .B(G148gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT5), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G176gat), .B(G204gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  OR2_X1    g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n496_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT13), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(KEYINPUT13), .A3(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n255_), .A2(new_n282_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n251_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n504_), .B1(new_n282_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT76), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n282_), .B(new_n505_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(G229gat), .A3(G233gat), .ZN(new_n511_));
  OAI22_X1  g310(.A1(new_n506_), .A2(new_n509_), .B1(new_n511_), .B2(KEYINPUT75), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(KEYINPUT75), .B2(new_n511_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G113gat), .B(G141gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT77), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT78), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G169gat), .B(G197gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n513_), .B(new_n518_), .Z(new_n519_));
  NOR2_X1   g318(.A1(new_n503_), .A2(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n483_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n307_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n423_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(KEYINPUT93), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(KEYINPUT93), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n522_), .A2(new_n277_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT38), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n304_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n267_), .A2(new_n268_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n521_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n523_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(G1gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n528_), .A2(new_n529_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n530_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT94), .Z(G1324gat));
  INV_X1    g338(.A(new_n381_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n522_), .A2(new_n278_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n540_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(G8gat), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n543_), .A2(KEYINPUT39), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(KEYINPUT39), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n541_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g346(.A(new_n438_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n534_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(G15gat), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT41), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT41), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n522_), .A2(new_n430_), .A3(new_n548_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(G1326gat));
  INV_X1    g353(.A(G22gat), .ZN(new_n555_));
  INV_X1    g354(.A(new_n469_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n534_), .B2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT42), .Z(new_n558_));
  NAND3_X1  g357(.A1(new_n522_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(G1327gat));
  INV_X1    g359(.A(new_n532_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(new_n304_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n521_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT97), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n521_), .A2(KEYINPUT97), .A3(new_n562_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(G29gat), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n523_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n469_), .A2(new_n548_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n523_), .B1(new_n570_), .B2(new_n465_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n571_), .A2(new_n381_), .B1(new_n481_), .B2(new_n470_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n275_), .A2(new_n305_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT43), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT95), .B1(new_n275_), .B2(new_n305_), .ZN(new_n576_));
  OAI22_X1  g375(.A1(new_n572_), .A2(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n483_), .A2(KEYINPUT95), .A3(KEYINPUT43), .A4(new_n573_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n520_), .A4(new_n531_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(KEYINPUT96), .A2(KEYINPUT44), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(KEYINPUT96), .A2(KEYINPUT44), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT44), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n580_), .A3(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n526_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n569_), .B1(new_n588_), .B2(new_n568_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT98), .ZN(G1328gat));
  NOR2_X1   g389(.A1(new_n381_), .A2(G36gat), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n565_), .A2(new_n566_), .A3(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT45), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n579_), .A2(new_n580_), .A3(new_n586_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n586_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n594_), .B(new_n540_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(G36gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n583_), .A2(new_n587_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n594_), .B1(new_n599_), .B2(new_n540_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n593_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT46), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI211_X1 g402(.A(KEYINPUT46), .B(new_n593_), .C1(new_n598_), .C2(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(G1329gat));
  INV_X1    g404(.A(G43gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n567_), .A2(new_n606_), .A3(new_n548_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n438_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n607_), .B1(new_n608_), .B2(new_n606_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g409(.A(G50gat), .B1(new_n567_), .B2(new_n556_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n556_), .A2(G50gat), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n599_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(G1331gat));
  NAND2_X1  g414(.A1(new_n503_), .A2(new_n519_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n572_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n307_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(G57gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(new_n527_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n617_), .A2(new_n533_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G57gat), .B1(new_n622_), .B2(new_n423_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(G1332gat));
  INV_X1    g423(.A(G64gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n618_), .A2(new_n625_), .A3(new_n540_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G64gat), .B1(new_n622_), .B2(new_n381_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(KEYINPUT48), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(KEYINPUT48), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n626_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT101), .ZN(G1333gat));
  INV_X1    g430(.A(G71gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n621_), .B2(new_n548_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT102), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT49), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(KEYINPUT49), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n618_), .A2(new_n632_), .A3(new_n548_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(G1334gat));
  INV_X1    g437(.A(G78gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n621_), .B2(new_n556_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT50), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n618_), .A2(new_n639_), .A3(new_n556_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1335gat));
  AND2_X1   g442(.A1(new_n617_), .A2(new_n562_), .ZN(new_n644_));
  INV_X1    g443(.A(G85gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(new_n527_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n577_), .A2(new_n531_), .A3(new_n578_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n616_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT103), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n650_), .B1(new_n647_), .B2(new_n616_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n423_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n646_), .B1(new_n652_), .B2(new_n645_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT104), .ZN(G1336gat));
  INV_X1    g453(.A(G92gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n644_), .A2(new_n655_), .A3(new_n540_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n381_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(new_n655_), .ZN(G1337gat));
  NAND4_X1  g457(.A1(new_n644_), .A2(new_n210_), .A3(new_n211_), .A4(new_n548_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n438_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n225_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g461(.A1(new_n644_), .A2(new_n226_), .A3(new_n556_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT52), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n648_), .A2(new_n556_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(G106gat), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT52), .B(new_n226_), .C1(new_n648_), .C2(new_n556_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT105), .B(KEYINPUT53), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n668_), .B(new_n670_), .ZN(G1339gat));
  INV_X1    g470(.A(new_n519_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(new_n497_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n484_), .A2(KEYINPUT108), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n485_), .A2(KEYINPUT55), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n491_), .B2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n486_), .A2(new_n490_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n678_), .B(new_n674_), .C1(KEYINPUT12), .C2(new_n488_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT55), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n491_), .B2(new_n485_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT107), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n684_), .B(new_n681_), .C1(new_n491_), .C2(new_n485_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n680_), .A2(new_n683_), .A3(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(KEYINPUT56), .A3(new_n496_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT56), .B1(new_n686_), .B2(new_n496_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(KEYINPUT109), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n690_), .B(KEYINPUT56), .C1(new_n686_), .C2(new_n496_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n673_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n508_), .B1(new_n506_), .B2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(new_n693_), .B2(new_n506_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n518_), .B1(new_n510_), .B2(new_n508_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n513_), .A2(new_n518_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n499_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n532_), .B1(new_n692_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT111), .B(KEYINPUT57), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n686_), .A2(new_n496_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT56), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n687_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n497_), .A2(new_n697_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n688_), .B2(KEYINPUT112), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n705_), .A2(KEYINPUT58), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n573_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT58), .B1(new_n705_), .B2(new_n707_), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n699_), .A2(new_n700_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n692_), .A2(new_n698_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n712_), .A2(KEYINPUT57), .A3(new_n561_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n531_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n503_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(KEYINPUT106), .A2(KEYINPUT54), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n306_), .A2(new_n519_), .A3(new_n715_), .A4(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n519_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n275_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  AOI22_X1  g520(.A1(new_n718_), .A2(new_n721_), .B1(KEYINPUT106), .B2(KEYINPUT54), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n714_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n527_), .A2(new_n381_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(new_n570_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT113), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G113gat), .B1(new_n728_), .B2(new_n672_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT114), .B(KEYINPUT59), .Z(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n724_), .A2(new_n727_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(KEYINPUT59), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n519_), .A2(KEYINPUT115), .ZN(new_n737_));
  MUX2_X1   g536(.A(KEYINPUT115), .B(new_n737_), .S(G113gat), .Z(new_n738_));
  AOI21_X1  g537(.A(new_n729_), .B1(new_n736_), .B2(new_n738_), .ZN(G1340gat));
  XOR2_X1   g538(.A(KEYINPUT116), .B(G120gat), .Z(new_n740_));
  INV_X1    g539(.A(KEYINPUT60), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(new_n715_), .B2(new_n740_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n724_), .A2(new_n727_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n503_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n735_), .B2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n728_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1341gat));
  INV_X1    g546(.A(G127gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n732_), .B2(new_n531_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT117), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n731_), .A2(new_n734_), .A3(G127gat), .A4(new_n304_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n750_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .ZN(G1342gat));
  OAI21_X1  g553(.A(G134gat), .B1(new_n735_), .B2(new_n574_), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n732_), .A2(G134gat), .A3(new_n561_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1343gat));
  INV_X1    g556(.A(new_n700_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n698_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n496_), .ZN(new_n760_));
  AOI22_X1  g559(.A1(KEYINPUT107), .A2(new_n682_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n685_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n690_), .B1(new_n762_), .B2(KEYINPUT56), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n688_), .A2(KEYINPUT109), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n687_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n759_), .B1(new_n765_), .B2(new_n673_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n758_), .B1(new_n766_), .B2(new_n532_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n712_), .A2(KEYINPUT57), .A3(new_n561_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n705_), .A2(new_n707_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n573_), .A3(new_n708_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n767_), .A2(new_n768_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n722_), .B1(new_n773_), .B2(new_n531_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n774_), .A2(new_n465_), .A3(new_n725_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n672_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n503_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g578(.A1(new_n774_), .A2(new_n465_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n725_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n304_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT118), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n775_), .A2(new_n784_), .A3(new_n304_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(KEYINPUT61), .B(G155gat), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n783_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1346gat));
  INV_X1    g590(.A(G162gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n775_), .A2(new_n792_), .A3(new_n532_), .ZN(new_n793_));
  NOR4_X1   g592(.A1(new_n774_), .A2(new_n465_), .A3(new_n574_), .A4(new_n725_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n792_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT119), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n793_), .B(new_n797_), .C1(new_n794_), .C2(new_n792_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1347gat));
  NOR3_X1   g598(.A1(new_n527_), .A2(new_n381_), .A3(new_n570_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n724_), .A2(KEYINPUT120), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n802_));
  INV_X1    g601(.A(new_n800_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n774_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n519_), .A2(new_n358_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n774_), .A2(new_n803_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n320_), .B1(new_n808_), .B2(new_n672_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n809_), .A2(new_n810_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n807_), .B1(new_n811_), .B2(new_n812_), .ZN(G1348gat));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n724_), .A2(new_n814_), .A3(new_n469_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT121), .B1(new_n774_), .B2(new_n556_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n527_), .A2(new_n381_), .A3(new_n438_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n715_), .A2(new_n321_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(KEYINPUT122), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(KEYINPUT122), .ZN(new_n821_));
  AOI21_X1  g620(.A(G176gat), .B1(new_n805_), .B2(new_n503_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(G1349gat));
  NAND4_X1  g622(.A1(new_n815_), .A2(new_n816_), .A3(new_n304_), .A4(new_n817_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n531_), .A2(new_n334_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n824_), .A2(new_n313_), .B1(new_n805_), .B2(new_n825_), .ZN(G1350gat));
  NAND3_X1  g625(.A1(new_n805_), .A2(new_n335_), .A3(new_n532_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT123), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT120), .B1(new_n724_), .B2(new_n800_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n774_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n573_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n831_), .B2(G190gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n574_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n833_), .A2(KEYINPUT123), .A3(new_n314_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n827_), .B1(new_n832_), .B2(new_n834_), .ZN(G1351gat));
  NOR4_X1   g634(.A1(new_n774_), .A2(new_n381_), .A3(new_n523_), .A4(new_n465_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n672_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g637(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT124), .B(G204gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n503_), .ZN(new_n841_));
  MUX2_X1   g640(.A(new_n839_), .B(new_n840_), .S(new_n841_), .Z(G1353gat));
  NAND2_X1  g641(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n304_), .A2(new_n843_), .ZN(new_n844_));
  XOR2_X1   g643(.A(new_n844_), .B(KEYINPUT125), .Z(new_n845_));
  NAND2_X1  g644(.A1(new_n836_), .A2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n847_), .A2(KEYINPUT126), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n847_), .B(KEYINPUT126), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n846_), .B2(new_n850_), .ZN(G1354gat));
  INV_X1    g650(.A(G218gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n381_), .A2(new_n523_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n780_), .A2(new_n852_), .A3(new_n532_), .A4(new_n853_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n780_), .A2(new_n573_), .A3(new_n853_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n852_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT127), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT127), .B(new_n854_), .C1(new_n855_), .C2(new_n852_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1355gat));
endmodule


