//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT99), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G226gat), .A2(G233gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G211gat), .B(G218gat), .Z(new_n208_));
  INV_X1    g007(.A(G204gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G197gat), .ZN(new_n210_));
  INV_X1    g009(.A(G197gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G204gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(KEYINPUT21), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n209_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n217_));
  OAI211_X1 g016(.A(KEYINPUT21), .B(new_n217_), .C1(new_n213_), .C2(KEYINPUT89), .ZN(new_n218_));
  INV_X1    g017(.A(new_n208_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n218_), .B(new_n219_), .C1(KEYINPUT21), .C2(new_n213_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT92), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT25), .B(G183gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n228_), .A2(KEYINPUT24), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G183gat), .ZN(new_n232_));
  INV_X1    g031(.A(G190gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT23), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G183gat), .A3(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n226_), .A2(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n225_), .A2(new_n231_), .A3(new_n237_), .A4(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT95), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G169gat), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n242_), .A2(KEYINPUT94), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(KEYINPUT94), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n243_), .A2(new_n244_), .A3(G176gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n230_), .B(KEYINPUT93), .Z(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n241_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n242_), .B(KEYINPUT94), .ZN(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT95), .B(new_n246_), .C1(new_n249_), .C2(G176gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n236_), .B(KEYINPUT82), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n234_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n232_), .A2(new_n233_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n248_), .A2(new_n250_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n221_), .B1(new_n240_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n216_), .A2(new_n220_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n228_), .A2(new_n229_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n238_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n224_), .A2(new_n222_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n252_), .A2(new_n231_), .A3(new_n259_), .A4(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n237_), .A2(new_n253_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT84), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT84), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n237_), .A2(new_n264_), .A3(new_n253_), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT22), .ZN(new_n267_));
  AOI21_X1  g066(.A(G176gat), .B1(new_n267_), .B2(KEYINPUT83), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(KEYINPUT83), .B2(new_n242_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n263_), .A2(new_n230_), .A3(new_n265_), .A4(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n261_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT20), .B1(new_n257_), .B2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n207_), .B1(new_n256_), .B2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G8gat), .B(G36gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G64gat), .B(G92gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n255_), .A2(new_n221_), .A3(new_n240_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT20), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n257_), .B2(new_n271_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n206_), .A3(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n273_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT27), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n206_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n272_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n255_), .A2(new_n240_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n206_), .B(new_n287_), .C1(new_n288_), .C2(new_n221_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n278_), .B1(new_n286_), .B2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n203_), .B1(new_n284_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292_));
  INV_X1    g091(.A(new_n283_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n278_), .B1(new_n273_), .B2(new_n282_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n278_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n256_), .A2(new_n207_), .A3(new_n272_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n296_), .B1(new_n297_), .B2(new_n285_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n298_), .A2(KEYINPUT99), .A3(KEYINPUT27), .A4(new_n283_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n291_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G1gat), .B(G29gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G85gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT0), .B(G57gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT1), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(G155gat), .A3(G162gat), .ZN(new_n309_));
  INV_X1    g108(.A(G155gat), .ZN(new_n310_));
  INV_X1    g109(.A(G162gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n307_), .A2(new_n309_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G141gat), .B(G148gat), .Z(new_n315_));
  OAI211_X1 g114(.A(new_n314_), .B(new_n315_), .C1(new_n313_), .C2(new_n309_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317_));
  INV_X1    g116(.A(G141gat), .ZN(new_n318_));
  INV_X1    g117(.A(G148gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n320_), .A2(new_n323_), .A3(new_n324_), .A4(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(new_n306_), .A3(new_n312_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n316_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT87), .ZN(new_n329_));
  XOR2_X1   g128(.A(G127gat), .B(G134gat), .Z(new_n330_));
  INV_X1    g129(.A(KEYINPUT85), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G127gat), .B(G134gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT85), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G113gat), .B(G120gat), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n332_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT87), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n316_), .A2(new_n339_), .A3(new_n327_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n329_), .A2(new_n338_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n328_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(KEYINPUT4), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n329_), .A2(new_n338_), .A3(new_n347_), .A4(new_n340_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n344_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n341_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n305_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n350_), .A3(new_n305_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G22gat), .B(G50gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT88), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n257_), .B(new_n358_), .C1(new_n359_), .C2(new_n342_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n329_), .A2(KEYINPUT29), .A3(new_n340_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n358_), .B1(new_n362_), .B2(new_n257_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n355_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n361_), .A2(new_n363_), .A3(new_n355_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n329_), .A2(new_n340_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT28), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n359_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n369_), .B1(new_n368_), .B2(new_n359_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n367_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n367_), .ZN(new_n375_));
  OAI22_X1  g174(.A1(new_n365_), .A2(new_n366_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n366_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n375_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n373_), .A4(new_n364_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n354_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n341_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n304_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT97), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT97), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n384_), .A3(new_n304_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n344_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT98), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n273_), .A2(new_n282_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n296_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n283_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n353_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n349_), .A2(KEYINPUT33), .A3(new_n350_), .A4(new_n305_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n394_), .B(new_n395_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n354_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n278_), .A2(KEYINPUT32), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n273_), .A2(new_n398_), .A3(new_n282_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n297_), .A2(new_n285_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(new_n398_), .ZN(new_n401_));
  OAI22_X1  g200(.A1(new_n392_), .A2(new_n396_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n376_), .A2(new_n379_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n300_), .A2(new_n380_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G43gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n271_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n338_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n409_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G227gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(G15gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT30), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT31), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n412_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n410_), .A2(new_n417_), .A3(new_n411_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n202_), .B1(new_n405_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n402_), .A2(new_n404_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n380_), .A2(new_n291_), .A3(new_n295_), .A4(new_n299_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(KEYINPUT100), .A3(new_n421_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n404_), .A2(new_n291_), .A3(new_n295_), .A4(new_n299_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n421_), .A2(new_n354_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT101), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT101), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n300_), .A2(new_n432_), .A3(new_n404_), .A4(new_n429_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n423_), .A2(new_n427_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT15), .ZN(new_n435_));
  INV_X1    g234(.A(G36gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G29gat), .ZN(new_n437_));
  INV_X1    g236(.A(G29gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G36gat), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n437_), .A2(new_n439_), .A3(KEYINPUT71), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT71), .B1(new_n437_), .B2(new_n439_), .ZN(new_n441_));
  INV_X1    g240(.A(G50gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G43gat), .ZN(new_n443_));
  INV_X1    g242(.A(G43gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G50gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n440_), .A2(new_n441_), .A3(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n443_), .A2(new_n445_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT71), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n438_), .A2(G36gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n436_), .A2(G29gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n437_), .A2(new_n439_), .A3(KEYINPUT71), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n448_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n435_), .B1(new_n447_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n446_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n453_), .A3(new_n448_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT15), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT14), .ZN(new_n460_));
  INV_X1    g259(.A(G1gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT74), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT74), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G1gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n460_), .B1(new_n465_), .B2(G8gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G15gat), .B(G22gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT75), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT75), .ZN(new_n470_));
  INV_X1    g269(.A(G8gat), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n471_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n470_), .B(new_n467_), .C1(new_n472_), .C2(new_n460_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G8gat), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n469_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n459_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT78), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT78), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n459_), .B(new_n480_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n474_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n473_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT74), .B(G1gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n484_), .B2(new_n471_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n470_), .B1(new_n485_), .B2(new_n467_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n482_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n447_), .A2(new_n454_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n469_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n478_), .A2(new_n479_), .A3(new_n481_), .A4(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT79), .ZN(new_n492_));
  INV_X1    g291(.A(new_n488_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n490_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n479_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n492_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n475_), .A2(new_n476_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n477_), .A2(KEYINPUT78), .B1(new_n499_), .B2(new_n488_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n500_), .A2(new_n492_), .A3(new_n479_), .A4(new_n481_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G113gat), .B(G141gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT80), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G169gat), .B(G197gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n498_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(G85gat), .ZN(new_n510_));
  INV_X1    g309(.A(G92gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518_));
  INV_X1    g317(.A(G99gat), .ZN(new_n519_));
  INV_X1    g318(.A(G106gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n514_), .B1(new_n517_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT8), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(new_n514_), .C1(new_n517_), .C2(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT64), .ZN(new_n530_));
  NAND2_X1  g329(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT64), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT65), .B(G106gat), .Z(new_n537_));
  AOI21_X1  g336(.A(new_n517_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n512_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT66), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n512_), .A2(new_n540_), .A3(new_n513_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT9), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n512_), .A2(new_n540_), .A3(KEYINPUT9), .A4(new_n513_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n539_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n538_), .B1(new_n545_), .B2(KEYINPUT67), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT67), .ZN(new_n547_));
  AOI211_X1 g346(.A(new_n547_), .B(new_n539_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n528_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT68), .B(G71gat), .ZN(new_n550_));
  INV_X1    g349(.A(G78gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n553_), .B(KEYINPUT11), .Z(new_n556_));
  OAI21_X1  g355(.A(new_n555_), .B1(new_n556_), .B2(new_n552_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n549_), .A2(KEYINPUT12), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT69), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n549_), .A2(new_n560_), .A3(KEYINPUT12), .A4(new_n557_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G230gat), .A2(G233gat), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT12), .B1(new_n549_), .B2(new_n557_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n549_), .A2(new_n557_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n562_), .A2(new_n563_), .A3(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n549_), .B(new_n557_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(G230gat), .A3(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT5), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G176gat), .B(G204gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n567_), .A2(new_n569_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n578_));
  NAND2_X1  g377(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OAI22_X1  g379(.A1(new_n576_), .A2(new_n577_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n577_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n549_), .A2(new_n459_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n528_), .B(new_n488_), .C1(new_n546_), .C2(new_n548_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n590_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n593_), .A2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n598_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n590_), .A2(new_n600_), .A3(new_n595_), .A4(new_n596_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT72), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n589_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n589_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n599_), .A2(KEYINPUT72), .A3(new_n605_), .A4(new_n601_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(KEYINPUT36), .A3(new_n588_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n604_), .A2(new_n607_), .A3(new_n606_), .A4(new_n609_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT77), .ZN(new_n614_));
  INV_X1    g413(.A(G231gat), .ZN(new_n615_));
  INV_X1    g414(.A(G233gat), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT17), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(G127gat), .A2(G155gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G127gat), .A2(G155gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(KEYINPUT16), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT16), .B1(new_n621_), .B2(new_n622_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n620_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n623_), .A3(new_n619_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n618_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT76), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n617_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n629_), .A2(new_n630_), .A3(new_n617_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n557_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n633_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n557_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n631_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n637_), .A3(new_n499_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n626_), .A2(new_n628_), .A3(new_n618_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n499_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n614_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n641_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n643_), .A2(KEYINPUT77), .A3(new_n639_), .A4(new_n638_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n613_), .A2(new_n645_), .ZN(new_n646_));
  NOR4_X1   g445(.A1(new_n434_), .A2(new_n509_), .A3(new_n585_), .A4(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n354_), .A3(new_n484_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT38), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n431_), .A2(new_n433_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT100), .B1(new_n426_), .B2(new_n421_), .ZN(new_n651_));
  AOI211_X1 g450(.A(new_n202_), .B(new_n422_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n608_), .B(KEYINPUT102), .Z(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT103), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n640_), .A2(new_n641_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n585_), .A2(new_n657_), .A3(new_n509_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(new_n354_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n649_), .B1(new_n660_), .B2(new_n461_), .ZN(G1324gat));
  INV_X1    g460(.A(new_n300_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n647_), .A2(new_n471_), .A3(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n656_), .A2(new_n662_), .A3(new_n658_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(G8gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n664_), .B2(G8gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(G1325gat));
  NAND3_X1  g469(.A1(new_n647_), .A2(new_n414_), .A3(new_n422_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n659_), .A2(new_n422_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n672_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT41), .B1(new_n672_), .B2(G15gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n673_), .B2(new_n674_), .ZN(G1326gat));
  INV_X1    g474(.A(G22gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n647_), .A2(new_n676_), .A3(new_n403_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n659_), .A2(new_n403_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(G22gat), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT42), .B(new_n676_), .C1(new_n659_), .C2(new_n403_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(G1327gat));
  INV_X1    g481(.A(new_n654_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n645_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NOR4_X1   g484(.A1(new_n434_), .A2(new_n509_), .A3(new_n585_), .A4(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n438_), .A3(new_n354_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  INV_X1    g487(.A(new_n613_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(KEYINPUT104), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n690_), .B1(new_n434_), .B2(new_n613_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n690_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n653_), .A2(new_n689_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n509_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n584_), .A2(new_n695_), .A3(new_n684_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT44), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n699_), .B(new_n696_), .C1(new_n691_), .C2(new_n693_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n698_), .A2(new_n700_), .A3(new_n397_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n687_), .B1(new_n701_), .B2(new_n438_), .ZN(G1328gat));
  NAND2_X1  g501(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n703_));
  NOR2_X1   g502(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n686_), .A2(new_n436_), .A3(new_n662_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT45), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(KEYINPUT45), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n698_), .A2(new_n700_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT105), .B1(new_n709_), .B2(new_n662_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n434_), .A2(new_n613_), .A3(new_n690_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n692_), .B1(new_n653_), .B2(new_n689_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n697_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n699_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n694_), .A2(KEYINPUT44), .A3(new_n697_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n714_), .A2(KEYINPUT105), .A3(new_n662_), .A4(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G36gat), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n703_), .B(new_n708_), .C1(new_n710_), .C2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n714_), .A2(new_n662_), .A3(new_n715_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(G36gat), .A3(new_n716_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n703_), .B1(new_n723_), .B2(new_n708_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n719_), .A2(new_n724_), .ZN(G1329gat));
  NAND3_X1  g524(.A1(new_n709_), .A2(G43gat), .A3(new_n422_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n686_), .A2(new_n422_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(new_n444_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n709_), .A2(new_n727_), .A3(G43gat), .A4(new_n422_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n730_), .B2(new_n732_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1330gat));
  NAND2_X1  g534(.A1(new_n403_), .A2(new_n442_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT109), .Z(new_n737_));
  NAND2_X1  g536(.A1(new_n686_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n709_), .A2(new_n403_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(G50gat), .ZN(new_n741_));
  AOI211_X1 g540(.A(KEYINPUT108), .B(new_n442_), .C1(new_n709_), .C2(new_n403_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(G1331gat));
  NOR4_X1   g542(.A1(new_n434_), .A2(new_n695_), .A3(new_n584_), .A4(new_n646_), .ZN(new_n744_));
  INV_X1    g543(.A(G57gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n354_), .ZN(new_n746_));
  AND4_X1   g545(.A1(new_n656_), .A2(new_n509_), .A3(new_n585_), .A4(new_n645_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(new_n354_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n748_), .B2(new_n745_), .ZN(G1332gat));
  NOR2_X1   g548(.A1(new_n300_), .A2(G64gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT110), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n744_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n747_), .A2(new_n662_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(G64gat), .ZN(new_n755_));
  INV_X1    g554(.A(G64gat), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT48), .B(new_n756_), .C1(new_n747_), .C2(new_n662_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n752_), .B1(new_n755_), .B2(new_n757_), .ZN(G1333gat));
  NOR2_X1   g557(.A1(new_n421_), .A2(G71gat), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT112), .Z(new_n760_));
  NAND2_X1  g559(.A1(new_n744_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n747_), .A2(new_n422_), .ZN(new_n762_));
  XOR2_X1   g561(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(G71gat), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G71gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(G1334gat));
  NAND3_X1  g565(.A1(new_n744_), .A2(new_n551_), .A3(new_n403_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n747_), .A2(new_n403_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(G78gat), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT50), .B(new_n551_), .C1(new_n747_), .C2(new_n403_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(G1335gat));
  NOR3_X1   g571(.A1(new_n584_), .A2(new_n695_), .A3(new_n645_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n397_), .ZN(new_n777_));
  NOR4_X1   g576(.A1(new_n434_), .A2(new_n695_), .A3(new_n584_), .A4(new_n685_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n510_), .A3(new_n354_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1336gat));
  OAI21_X1  g579(.A(G92gat), .B1(new_n776_), .B2(new_n300_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n511_), .A3(new_n662_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n776_), .B2(new_n421_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n778_), .A2(new_n536_), .A3(new_n422_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g586(.A1(new_n778_), .A2(new_n537_), .A3(new_n403_), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n404_), .B(new_n774_), .C1(new_n691_), .C2(new_n693_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n520_), .B1(new_n789_), .B2(KEYINPUT113), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n775_), .A2(new_n403_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n790_), .A2(new_n791_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n790_), .B2(new_n794_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n788_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n788_), .B(new_n798_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1339gat));
  NOR3_X1   g601(.A1(new_n428_), .A2(new_n397_), .A3(new_n421_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n498_), .A2(new_n501_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n505_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n500_), .A2(new_n496_), .A3(new_n481_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n505_), .B1(new_n495_), .B2(new_n479_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(KEYINPUT119), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n508_), .B2(new_n809_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n576_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n563_), .B1(new_n562_), .B2(new_n566_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n567_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n562_), .A2(KEYINPUT55), .A3(new_n563_), .A4(new_n566_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n819_), .B2(new_n573_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n821_), .B(new_n574_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n814_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n814_), .B(KEYINPUT58), .C1(new_n820_), .C2(new_n822_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n689_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n582_), .A2(new_n575_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT119), .B1(new_n806_), .B2(new_n810_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n508_), .A2(new_n812_), .A3(new_n809_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n828_), .B(KEYINPUT120), .C1(new_n829_), .C2(new_n830_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n820_), .A2(new_n822_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT118), .B1(new_n509_), .B2(new_n576_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n575_), .B(new_n837_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n833_), .B(new_n834_), .C1(new_n835_), .C2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n654_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n840_), .B2(new_n654_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n827_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n657_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n645_), .A2(new_n847_), .A3(new_n509_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n498_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n806_), .A2(new_n642_), .A3(new_n644_), .A4(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT115), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n584_), .A2(new_n613_), .A3(new_n848_), .A4(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT54), .B1(new_n852_), .B2(KEYINPUT116), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855_));
  INV_X1    g654(.A(new_n852_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n852_), .A2(KEYINPUT116), .A3(KEYINPUT117), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n854_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n856_), .A2(new_n857_), .A3(new_n855_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT117), .B1(new_n852_), .B2(KEYINPUT116), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n853_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n804_), .B1(new_n846_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n695_), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n845_), .A2(new_n684_), .B1(new_n863_), .B2(new_n860_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n804_), .A2(KEYINPUT59), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n865_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n827_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n840_), .A2(new_n654_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT57), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n877_), .B2(new_n842_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n657_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n864_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n803_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n871_), .B1(new_n874_), .B2(new_n882_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n883_), .A2(new_n695_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n867_), .B1(new_n884_), .B2(new_n866_), .ZN(G1340gat));
  INV_X1    g684(.A(new_n871_), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(new_n881_), .B2(KEYINPUT59), .ZN(new_n887_));
  AOI211_X1 g686(.A(new_n872_), .B(new_n873_), .C1(new_n880_), .C2(new_n803_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n585_), .B(new_n886_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n874_), .A2(new_n882_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n892_), .A2(KEYINPUT122), .A3(new_n585_), .A4(new_n886_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(G120gat), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(G120gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n584_), .B2(KEYINPUT60), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n865_), .B(new_n896_), .C1(KEYINPUT60), .C2(new_n895_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n897_), .ZN(G1341gat));
  AOI21_X1  g697(.A(G127gat), .B1(new_n865_), .B2(new_n645_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT123), .B(G127gat), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n657_), .A2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n883_), .B2(new_n901_), .ZN(G1342gat));
  INV_X1    g701(.A(G134gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n865_), .A2(new_n903_), .A3(new_n683_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n883_), .A2(new_n689_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n903_), .ZN(G1343gat));
  NOR3_X1   g705(.A1(new_n404_), .A2(new_n422_), .A3(new_n397_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n880_), .A2(new_n300_), .A3(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n509_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n318_), .ZN(G1344gat));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n584_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT124), .B(G148gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1345gat));
  NOR2_X1   g712(.A1(new_n908_), .A2(new_n684_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT61), .B(G155gat), .Z(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n908_), .B2(new_n613_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n683_), .A2(new_n311_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n908_), .B2(new_n918_), .ZN(G1347gat));
  NOR3_X1   g718(.A1(new_n300_), .A2(new_n430_), .A3(new_n403_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n868_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n695_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n266_), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n923_), .B(new_n924_), .C1(KEYINPUT125), .C2(KEYINPUT62), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n249_), .B2(new_n923_), .ZN(new_n926_));
  AOI211_X1 g725(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n923_), .C2(G169gat), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1348gat));
  AOI21_X1  g727(.A(G176gat), .B1(new_n922_), .B2(new_n585_), .ZN(new_n929_));
  AND4_X1   g728(.A1(G176gat), .A2(new_n880_), .A3(new_n585_), .A4(new_n920_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1349gat));
  NOR2_X1   g730(.A1(new_n657_), .A2(new_n224_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n880_), .A2(new_n645_), .A3(new_n920_), .ZN(new_n933_));
  AOI22_X1  g732(.A1(new_n922_), .A2(new_n932_), .B1(new_n933_), .B2(new_n232_), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n922_), .A2(new_n683_), .A3(new_n223_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n868_), .A2(new_n613_), .A3(new_n921_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n233_), .ZN(G1351gat));
  NAND3_X1  g736(.A1(new_n662_), .A2(new_n380_), .A3(new_n421_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n846_), .B2(new_n864_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n695_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n585_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT126), .B(G204gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1353gat));
  NAND2_X1  g743(.A1(new_n939_), .A2(new_n879_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n945_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(KEYINPUT63), .B(G211gat), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n939_), .A2(new_n879_), .A3(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(new_n949_));
  XOR2_X1   g748(.A(new_n949_), .B(KEYINPUT127), .Z(G1354gat));
  INV_X1    g749(.A(G218gat), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n939_), .A2(new_n951_), .A3(new_n683_), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n939_), .A2(new_n689_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n953_), .B2(new_n951_), .ZN(G1355gat));
endmodule


