//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT85), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR3_X1   g009(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n208_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n208_), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT82), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n218_), .A2(new_n209_), .A3(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n212_), .A2(new_n217_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT81), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT26), .B(G190gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT80), .B1(new_n227_), .B2(G183gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT25), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(G183gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT80), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n225_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT26), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT26), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G190gat), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n228_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n231_), .A2(new_n232_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT80), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n239_), .A2(new_n242_), .A3(KEYINPUT81), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n224_), .B1(new_n234_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n213_), .B(KEYINPUT23), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n230_), .A2(new_n235_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(KEYINPUT84), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n215_), .A2(new_n216_), .A3(new_n246_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT84), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT83), .B(G176gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT22), .B(G169gat), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n251_), .A2(new_n252_), .B1(G169gat), .B2(G176gat), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n247_), .A2(new_n250_), .A3(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n207_), .B1(new_n244_), .B2(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n212_), .A2(new_n217_), .A3(new_n223_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT81), .B1(new_n239_), .B2(new_n242_), .ZN(new_n257_));
  NOR3_X1   g056(.A1(new_n229_), .A2(new_n233_), .A3(new_n225_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n247_), .A2(new_n250_), .A3(new_n253_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT85), .A3(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(G197gat), .A2(G204gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G197gat), .A2(G204gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT21), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(KEYINPUT21), .A3(new_n263_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n267_), .A2(new_n268_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n255_), .A2(new_n261_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n253_), .A2(new_n248_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT95), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n208_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n245_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n245_), .B2(new_n277_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT25), .B(G183gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n226_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n223_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n275_), .B1(new_n280_), .B2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n274_), .B1(new_n284_), .B2(new_n271_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n273_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G226gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT19), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n244_), .A2(new_n254_), .A3(new_n207_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT85), .B1(new_n259_), .B2(new_n260_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n271_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n272_), .B(new_n275_), .C1(new_n280_), .C2(new_n283_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n294_), .A2(KEYINPUT20), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n290_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n206_), .B1(new_n289_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n272_), .B1(new_n255_), .B2(new_n261_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(KEYINPUT20), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n299_), .A2(new_n288_), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n290_), .B1(new_n273_), .B2(new_n285_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n206_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n298_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n206_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n286_), .A2(new_n288_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n293_), .A2(new_n290_), .A3(new_n295_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(new_n304_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n297_), .A2(new_n305_), .B1(new_n310_), .B2(new_n298_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT103), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n298_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n297_), .A2(KEYINPUT27), .A3(new_n309_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT103), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT94), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT88), .ZN(new_n321_));
  INV_X1    g120(.A(G141gat), .ZN(new_n322_));
  INV_X1    g121(.A(G148gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n325_));
  AND3_X1   g124(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n324_), .B(new_n325_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n330_), .A2(new_n331_), .A3(KEYINPUT1), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n321_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n324_), .A2(new_n325_), .ZN(new_n334_));
  OR2_X1    g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n329_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT87), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n334_), .A2(new_n337_), .A3(new_n342_), .A4(KEYINPUT88), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT90), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(KEYINPUT90), .B(new_n344_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT91), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n351_), .B(KEYINPUT89), .C1(G141gat), .C2(G148gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n322_), .B(new_n323_), .C1(new_n351_), .C2(KEYINPUT89), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n351_), .A2(KEYINPUT89), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .A4(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n330_), .A2(new_n331_), .ZN(new_n357_));
  AOI221_X4 g156(.A(KEYINPUT92), .B1(new_n333_), .B2(new_n343_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT92), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n357_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n333_), .A2(new_n343_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n320_), .B1(new_n358_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT28), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n365_), .B(new_n320_), .C1(new_n358_), .C2(new_n362_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G22gat), .B(G50gat), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n319_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n360_), .A2(new_n361_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT92), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n360_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n365_), .B1(new_n375_), .B2(new_n320_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n366_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n371_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(KEYINPUT94), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G78gat), .B(G106gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT93), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n373_), .A2(KEYINPUT29), .A3(new_n374_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n385_), .B1(new_n386_), .B2(new_n271_), .ZN(new_n387_));
  AOI211_X1 g186(.A(new_n272_), .B(new_n384_), .C1(new_n372_), .C2(KEYINPUT29), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n382_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n388_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n358_), .A2(new_n362_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n272_), .B1(new_n391_), .B2(KEYINPUT29), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n381_), .B(new_n390_), .C1(new_n392_), .C2(new_n385_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n370_), .A2(new_n380_), .A3(new_n389_), .A4(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n393_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n395_), .A2(KEYINPUT94), .A3(new_n379_), .A4(new_n378_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n318_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n255_), .A2(new_n261_), .A3(KEYINPUT30), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT86), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G71gat), .B(G99gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G43gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  INV_X1    g205(.A(G15gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n405_), .B(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n403_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(G134gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(G127gat), .ZN(new_n412_));
  INV_X1    g211(.A(G127gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G134gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G120gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G113gat), .ZN(new_n417_));
  INV_X1    g216(.A(G113gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G120gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n412_), .A2(new_n414_), .A3(new_n417_), .A4(new_n419_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT31), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n402_), .A2(KEYINPUT86), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n425_), .A2(new_n403_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n410_), .B(new_n424_), .C1(new_n426_), .C2(new_n409_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n424_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n409_), .B1(new_n425_), .B2(new_n403_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n410_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT97), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n421_), .A2(new_n422_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT98), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT98), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n436_), .A2(new_n360_), .A3(new_n439_), .A4(new_n361_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n373_), .A2(new_n374_), .A3(new_n423_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G225gat), .A2(G233gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n441_), .A2(new_n442_), .A3(KEYINPUT4), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n373_), .A2(new_n446_), .A3(new_n374_), .A4(new_n423_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n443_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n444_), .B1(new_n445_), .B2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G1gat), .B(G29gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G85gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT0), .B(G57gat), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n452_), .B(new_n453_), .Z(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n444_), .B(new_n454_), .C1(new_n445_), .C2(new_n449_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(KEYINPUT101), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT101), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n450_), .A2(new_n459_), .A3(new_n455_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n432_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n398_), .A2(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n427_), .A2(new_n431_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n316_), .B1(new_n460_), .B2(new_n458_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n465_), .B2(new_n397_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT99), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n457_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT33), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n391_), .A2(new_n423_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n454_), .B1(new_n470_), .B2(new_n448_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n441_), .A2(new_n442_), .A3(KEYINPUT4), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT100), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(new_n310_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT33), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n457_), .A2(new_n467_), .A3(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT100), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n469_), .A2(new_n475_), .A3(new_n477_), .A4(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n289_), .A2(new_n296_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n304_), .A2(KEYINPUT32), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(new_n303_), .B2(new_n481_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n458_), .A2(new_n483_), .A3(new_n460_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n479_), .A2(new_n397_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT102), .B1(new_n466_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n457_), .A2(KEYINPUT101), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n472_), .A2(new_n448_), .A3(new_n447_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n454_), .B1(new_n488_), .B2(new_n444_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n460_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n311_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n394_), .A2(new_n396_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n432_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT102), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n479_), .A2(new_n397_), .A3(new_n484_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n463_), .B1(new_n486_), .B2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT72), .B(G15gat), .ZN(new_n499_));
  INV_X1    g298(.A(G22gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G1gat), .ZN(new_n502_));
  INV_X1    g301(.A(G8gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT14), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G1gat), .B(G8gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n506_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n501_), .A2(new_n508_), .A3(new_n504_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G29gat), .B(G36gat), .Z(new_n511_));
  XOR2_X1   g310(.A(G43gat), .B(G50gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT78), .B1(new_n510_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT78), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n507_), .A2(new_n516_), .A3(new_n509_), .A4(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n510_), .A2(new_n514_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT79), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n515_), .A2(new_n517_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT79), .B1(new_n525_), .B2(new_n522_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n513_), .B(KEYINPUT15), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n510_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n518_), .A2(new_n522_), .A3(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n524_), .A2(new_n526_), .A3(new_n529_), .A4(new_n533_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  XOR2_X1   g340(.A(G71gat), .B(G78gat), .Z(new_n542_));
  OR2_X1    g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n542_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n543_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT67), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT67), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n543_), .B(new_n548_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT68), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G85gat), .B(G92gat), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT9), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(KEYINPUT10), .B(G99gat), .Z(new_n556_));
  INV_X1    g355(.A(G106gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT6), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(G85gat), .A3(G92gat), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n555_), .A2(new_n558_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT64), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n553_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT8), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT7), .ZN(new_n566_));
  INV_X1    g365(.A(G99gat), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n557_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n560_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n564_), .A2(new_n565_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n569_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT65), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(KEYINPUT65), .A3(new_n569_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n560_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n565_), .B1(new_n576_), .B2(new_n564_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n562_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT12), .A4(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n578_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n547_), .A2(KEYINPUT12), .A3(new_n549_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT68), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G230gat), .A2(G233gat), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n562_), .B(new_n546_), .C1(new_n571_), .C2(new_n577_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT12), .ZN(new_n587_));
  INV_X1    g386(.A(new_n546_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n578_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n586_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n583_), .A2(new_n584_), .A3(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n585_), .A2(KEYINPUT66), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(KEYINPUT66), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(G230gat), .A3(G233gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT5), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT69), .Z(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n591_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT13), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT13), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n606_), .A3(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n578_), .A2(new_n527_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT34), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT35), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n513_), .B(new_n562_), .C1(new_n571_), .C2(new_n577_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n611_), .A2(KEYINPUT35), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n609_), .A2(new_n612_), .A3(new_n613_), .A4(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n612_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT70), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AOI211_X1 g417(.A(KEYINPUT70), .B(new_n612_), .C1(new_n609_), .C2(new_n613_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G134gat), .B(G162gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(G190gat), .B(G218gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT71), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n627_), .B(new_n615_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n624_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n626_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT37), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT73), .Z(new_n635_));
  XOR2_X1   g434(.A(new_n510_), .B(new_n635_), .Z(new_n636_));
  XNOR2_X1  g435(.A(new_n550_), .B(KEYINPUT74), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n640_));
  XOR2_X1   g439(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT76), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G127gat), .B(G155gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(G183gat), .B(G211gat), .Z(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  OR4_X1    g445(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .A4(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(KEYINPUT17), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n636_), .A2(new_n546_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n636_), .A2(new_n546_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT37), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n653_), .B(new_n626_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n608_), .A2(new_n633_), .A3(new_n652_), .A4(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n498_), .A2(new_n539_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n461_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n502_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n498_), .A2(new_n632_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n608_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n652_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n662_), .A2(new_n539_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G1gat), .B1(new_n665_), .B2(new_n461_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n658_), .A2(new_n659_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n660_), .A2(new_n666_), .A3(new_n667_), .ZN(G1324gat));
  INV_X1    g467(.A(new_n318_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n656_), .A2(new_n503_), .A3(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT104), .ZN(new_n671_));
  OAI21_X1  g470(.A(G8gat), .B1(new_n665_), .B2(new_n318_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT39), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n673_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n676_), .B(new_n678_), .ZN(G1325gat));
  OAI21_X1  g478(.A(G15gat), .B1(new_n665_), .B2(new_n464_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT41), .Z(new_n681_));
  NAND3_X1  g480(.A1(new_n656_), .A2(new_n407_), .A3(new_n432_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1326gat));
  OAI21_X1  g482(.A(G22gat), .B1(new_n665_), .B2(new_n397_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT42), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n656_), .A2(new_n500_), .A3(new_n493_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1327gat));
  NOR2_X1   g486(.A1(new_n498_), .A2(new_n539_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n632_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n662_), .A2(new_n652_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G29gat), .B1(new_n692_), .B2(new_n657_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n539_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n608_), .A2(new_n663_), .A3(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT106), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n633_), .A2(new_n654_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n498_), .A2(KEYINPUT43), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n398_), .A2(new_n462_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n492_), .A2(new_n493_), .ZN(new_n703_));
  AND4_X1   g502(.A1(new_n495_), .A2(new_n496_), .A3(new_n703_), .A4(new_n464_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n495_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n701_), .B1(new_n706_), .B2(new_n698_), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT44), .B(new_n697_), .C1(new_n700_), .C2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n498_), .B2(new_n699_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n706_), .A2(new_n701_), .A3(new_n698_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n696_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n657_), .A2(G29gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n693_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  NOR3_X1   g515(.A1(new_n691_), .A2(G36gat), .A3(new_n318_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G36gat), .B1(new_n713_), .B2(new_n318_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n719_), .A2(new_n720_), .A3(KEYINPUT46), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  NAND2_X1  g524(.A1(new_n432_), .A2(G43gat), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n691_), .A2(new_n464_), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n713_), .A2(new_n726_), .B1(G43gat), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g528(.A1(new_n691_), .A2(G50gat), .A3(new_n397_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n708_), .B(new_n493_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n731_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT108), .B1(new_n731_), .B2(G50gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n730_), .B1(new_n732_), .B2(new_n733_), .ZN(G1331gat));
  NOR3_X1   g533(.A1(new_n608_), .A2(new_n663_), .A3(new_n694_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n661_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G57gat), .B1(new_n736_), .B2(new_n461_), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT109), .B1(new_n498_), .B2(new_n694_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n706_), .A2(new_n739_), .A3(new_n539_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n698_), .A2(new_n663_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n738_), .A2(new_n740_), .A3(new_n662_), .A4(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n461_), .A2(G57gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n737_), .B1(new_n742_), .B2(new_n743_), .ZN(G1332gat));
  OAI21_X1  g543(.A(G64gat), .B1(new_n736_), .B2(new_n318_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT48), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n318_), .A2(G64gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n742_), .B2(new_n747_), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n736_), .B2(new_n464_), .ZN(new_n749_));
  XOR2_X1   g548(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n464_), .A2(G71gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n742_), .B2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n736_), .B2(new_n397_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n742_), .A2(G78gat), .A3(new_n397_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT111), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n759_), .A3(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1335gat));
  NOR2_X1   g560(.A1(new_n689_), .A2(new_n652_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n738_), .A2(new_n740_), .A3(new_n662_), .A4(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(G85gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n657_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n608_), .A2(new_n694_), .A3(new_n652_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(new_n657_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n765_), .B2(new_n770_), .ZN(G1336gat));
  INV_X1    g570(.A(G92gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n764_), .A2(new_n772_), .A3(new_n669_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n769_), .A2(new_n669_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n772_), .B2(new_n774_), .ZN(G1337gat));
  NAND3_X1  g574(.A1(new_n764_), .A2(new_n432_), .A3(new_n556_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n769_), .A2(new_n432_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n567_), .B2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g578(.A(new_n493_), .B(new_n767_), .C1(new_n700_), .C2(new_n707_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(G106gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(G106gat), .ZN(new_n783_));
  XOR2_X1   g582(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n784_));
  NOR3_X1   g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n397_), .B(new_n768_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT113), .B(new_n784_), .C1(new_n786_), .C2(new_n557_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n764_), .A2(new_n557_), .A3(new_n493_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT53), .B1(new_n785_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT113), .B1(new_n786_), .B2(new_n557_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n780_), .A2(new_n781_), .A3(G106gat), .ZN(new_n792_));
  INV_X1    g591(.A(new_n784_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n787_), .A4(new_n788_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n790_), .A2(new_n796_), .ZN(G1339gat));
  OAI21_X1  g596(.A(new_n603_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n591_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n583_), .A2(KEYINPUT55), .A3(new_n590_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(KEYINPUT114), .A2(G230gat), .A3(G233gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n802_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n583_), .A2(KEYINPUT55), .A3(new_n590_), .A4(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n805_), .A2(new_n601_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT56), .B1(new_n803_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n806_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n798_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n518_), .A2(new_n523_), .A3(new_n528_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n534_), .C1(new_n523_), .C2(new_n525_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n604_), .A2(new_n537_), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n689_), .B1(new_n810_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT57), .B(new_n689_), .C1(new_n810_), .C2(new_n814_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n603_), .A2(new_n537_), .A3(new_n812_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n698_), .B(KEYINPUT115), .C1(new_n820_), .C2(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(KEYINPUT58), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n819_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n809_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n807_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT115), .B1(new_n828_), .B2(new_n698_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n817_), .B(new_n818_), .C1(new_n823_), .C2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n663_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n741_), .A2(new_n832_), .A3(new_n539_), .A4(new_n608_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT54), .B1(new_n655_), .B2(new_n694_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n831_), .A2(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n398_), .A2(new_n461_), .A3(new_n464_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n418_), .B1(new_n839_), .B2(new_n539_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n841_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n835_), .B1(new_n830_), .B2(new_n663_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n838_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n844_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT118), .B1(new_n844_), .B2(KEYINPUT117), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n817_), .A2(new_n818_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n698_), .B1(new_n820_), .B2(KEYINPUT58), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n822_), .A3(new_n821_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n652_), .B1(new_n851_), .B2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n838_), .B(new_n850_), .C1(new_n856_), .C2(new_n835_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n849_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n539_), .A2(new_n418_), .ZN(new_n859_));
  AOI22_X1  g658(.A1(new_n842_), .A2(new_n843_), .B1(new_n858_), .B2(new_n859_), .ZN(G1340gat));
  OAI21_X1  g659(.A(new_n416_), .B1(new_n608_), .B2(KEYINPUT60), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n416_), .A2(KEYINPUT60), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n837_), .A2(new_n838_), .A3(new_n861_), .A4(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n608_), .B1(new_n849_), .B2(new_n857_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n416_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT119), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n863_), .B(new_n867_), .C1(new_n864_), .C2(new_n416_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1341gat));
  INV_X1    g668(.A(new_n839_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(new_n413_), .A3(new_n652_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n663_), .B1(new_n849_), .B2(new_n857_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n413_), .ZN(G1342gat));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n411_), .A3(new_n632_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n699_), .B1(new_n849_), .B2(new_n857_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n411_), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n464_), .A2(new_n493_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n669_), .A2(new_n877_), .A3(new_n461_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n837_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n694_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n662_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g683(.A1(new_n880_), .A2(new_n652_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n879_), .B2(new_n699_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n689_), .A2(G162gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n879_), .B2(new_n889_), .ZN(G1347gat));
  NAND2_X1  g689(.A1(new_n669_), .A2(new_n461_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n464_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n837_), .A2(new_n397_), .A3(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(new_n252_), .A3(new_n694_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n892_), .A2(new_n694_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT120), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n837_), .A2(new_n397_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(G169gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(G169gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n895_), .B1(new_n900_), .B2(new_n901_), .ZN(G1348gat));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n903_), .B(new_n251_), .C1(new_n893_), .C2(new_n608_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n894_), .A2(new_n662_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n221_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n903_), .B1(new_n905_), .B2(new_n251_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1349gat));
  NAND2_X1  g707(.A1(new_n894_), .A2(new_n652_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(G183gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n281_), .B1(KEYINPUT122), .B2(G183gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n909_), .B2(new_n912_), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n893_), .B2(new_n699_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n632_), .A2(new_n226_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n893_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n914_), .B(KEYINPUT123), .C1(new_n893_), .C2(new_n915_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1351gat));
  NOR2_X1   g719(.A1(new_n891_), .A2(new_n877_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT124), .B1(new_n845_), .B2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n924_), .B(new_n921_), .C1(new_n856_), .C2(new_n835_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n694_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT125), .B(G197gat), .Z(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1352gat));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n662_), .ZN(new_n930_));
  AOI21_X1  g729(.A(KEYINPUT126), .B1(new_n930_), .B2(G204gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n608_), .B1(new_n923_), .B2(new_n925_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933_));
  INV_X1    g732(.A(G204gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936_));
  AND4_X1   g735(.A1(new_n936_), .A2(new_n926_), .A3(new_n934_), .A4(new_n662_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n932_), .B2(new_n934_), .ZN(new_n938_));
  OAI22_X1  g737(.A1(new_n931_), .A2(new_n935_), .B1(new_n937_), .B2(new_n938_), .ZN(G1353gat));
  OR2_X1    g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  NAND2_X1  g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  AND4_X1   g740(.A1(new_n652_), .A2(new_n926_), .A3(new_n940_), .A4(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n926_), .B2(new_n652_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1354gat));
  INV_X1    g743(.A(new_n926_), .ZN(new_n945_));
  OR3_X1    g744(.A1(new_n945_), .A2(G218gat), .A3(new_n689_), .ZN(new_n946_));
  OAI21_X1  g745(.A(G218gat), .B1(new_n945_), .B2(new_n699_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1355gat));
endmodule


