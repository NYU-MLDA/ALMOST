//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(G169gat), .B1(KEYINPUT84), .B2(KEYINPUT22), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n206_), .B1(KEYINPUT84), .B2(KEYINPUT22), .ZN(new_n207_));
  INV_X1    g006(.A(G169gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT22), .ZN(new_n209_));
  AOI21_X1  g008(.A(G176gat), .B1(new_n209_), .B2(KEYINPUT83), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(KEYINPUT83), .B2(new_n209_), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n204_), .B(new_n205_), .C1(new_n207_), .C2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT25), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT77), .B1(new_n214_), .B2(G183gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT26), .B(G190gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n215_), .B(new_n216_), .C1(new_n217_), .C2(KEYINPUT77), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT79), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR3_X1   g021(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n220_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n208_), .A3(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(KEYINPUT79), .A3(new_n221_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n205_), .A2(KEYINPUT24), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n219_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  AOI211_X1 g031(.A(KEYINPUT80), .B(new_n230_), .C1(new_n224_), .C2(new_n228_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n213_), .B(new_n218_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n224_), .A2(new_n235_), .A3(new_n228_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n203_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n236_), .B2(new_n203_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n234_), .A2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n227_), .A2(KEYINPUT79), .A3(new_n221_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT79), .B1(new_n227_), .B2(new_n221_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n231_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT80), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n230_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n219_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n213_), .B1(new_n248_), .B2(new_n218_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n212_), .B1(new_n241_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT30), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n218_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT81), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(new_n234_), .A3(new_n240_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT30), .A3(new_n212_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(KEYINPUT86), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G227gat), .A2(G233gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT85), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G71gat), .B(G99gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G15gat), .B(G43gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n257_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G127gat), .B(G134gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G113gat), .B(G120gat), .Z(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G113gat), .B(G120gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n268_), .A2(KEYINPUT87), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT87), .B1(new_n268_), .B2(new_n270_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT31), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n264_), .B1(KEYINPUT88), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n252_), .A2(new_n256_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT86), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n263_), .B1(new_n278_), .B2(new_n257_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n274_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT88), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  OR3_X1    g081(.A1(new_n275_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n282_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n285_));
  XOR2_X1   g084(.A(G155gat), .B(G162gat), .Z(new_n286_));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT89), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(KEYINPUT89), .A2(G141gat), .A3(G148gat), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G141gat), .ZN(new_n294_));
  INV_X1    g093(.A(G148gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n288_), .A2(new_n293_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n291_), .A2(new_n299_), .A3(new_n292_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n302_), .B(new_n303_), .C1(new_n299_), .C2(new_n289_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n286_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n268_), .A2(KEYINPUT87), .A3(new_n270_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n268_), .A2(new_n270_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT87), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n298_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n285_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT4), .B1(new_n273_), .B2(new_n306_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n312_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n315_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G1gat), .B(G29gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G85gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT0), .B(G57gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n316_), .A2(new_n319_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(KEYINPUT4), .ZN(new_n326_));
  INV_X1    g125(.A(new_n314_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n315_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n323_), .B1(new_n329_), .B2(new_n318_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n283_), .A2(new_n284_), .A3(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G22gat), .B(G50gat), .Z(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(new_n306_), .B2(KEYINPUT29), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335_));
  INV_X1    g134(.A(new_n333_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n298_), .A2(new_n305_), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G211gat), .B(G218gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT21), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(KEYINPUT91), .ZN(new_n344_));
  OR2_X1    g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n346_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n343_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n341_), .A2(new_n345_), .A3(new_n346_), .A4(new_n344_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT92), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n348_), .A2(new_n351_), .A3(KEYINPUT92), .A4(new_n350_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n306_), .A2(KEYINPUT29), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n335_), .B1(new_n298_), .B2(new_n305_), .ZN(new_n360_));
  OAI211_X1 g159(.A(G228gat), .B(G233gat), .C1(new_n360_), .C2(new_n352_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G78gat), .B(G106gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT94), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(new_n361_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT94), .A3(new_n362_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n340_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n362_), .A2(KEYINPUT93), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n359_), .B(new_n361_), .C1(KEYINPUT93), .C2(new_n362_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n369_), .A2(new_n370_), .B1(KEYINPUT93), .B2(new_n362_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n367_), .B1(new_n371_), .B2(new_n340_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT22), .B(G169gat), .Z(new_n374_));
  OAI211_X1 g173(.A(new_n204_), .B(new_n205_), .C1(G176gat), .C2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n235_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n217_), .A2(new_n216_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n203_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n375_), .B(new_n352_), .C1(new_n246_), .C2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT95), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n246_), .A2(new_n378_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n375_), .A4(new_n352_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT19), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT20), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n380_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n250_), .B2(new_n356_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n356_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n212_), .B(new_n391_), .C1(new_n241_), .C2(new_n249_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n352_), .B1(new_n381_), .B2(new_n375_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(new_n386_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n385_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n390_), .A2(new_n396_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n385_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n401_), .B1(new_n405_), .B2(new_n389_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT27), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n391_), .B1(new_n255_), .B2(new_n212_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n379_), .A2(KEYINPUT20), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n385_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n392_), .A2(new_n404_), .A3(new_n394_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n402_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n405_), .A2(new_n389_), .A3(new_n401_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  NOR4_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .A4(new_n408_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n405_), .A2(new_n389_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n408_), .B1(new_n418_), .B2(new_n402_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n411_), .B1(new_n250_), .B2(new_n356_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n413_), .B1(new_n420_), .B2(new_n404_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n401_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT99), .B1(new_n419_), .B2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n373_), .B(new_n409_), .C1(new_n417_), .C2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n332_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n372_), .A2(new_n331_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n417_), .B2(new_n423_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT100), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n402_), .A2(KEYINPUT32), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n421_), .A2(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n325_), .A2(new_n330_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n390_), .A2(new_n396_), .A3(new_n431_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT98), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT98), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .A4(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n315_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n311_), .A2(new_n312_), .A3(new_n328_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n323_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT97), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(KEYINPUT33), .B(new_n324_), .C1(new_n316_), .C2(new_n319_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n440_), .A2(KEYINPUT97), .A3(new_n323_), .A4(new_n441_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n330_), .A2(KEYINPUT33), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n447_), .A2(new_n403_), .A3(new_n406_), .A4(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n437_), .A2(new_n439_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n373_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n427_), .B(KEYINPUT100), .C1(new_n417_), .C2(new_n423_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n430_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n283_), .A2(new_n284_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n425_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G29gat), .B(G36gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G43gat), .B(G50gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT15), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G8gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT73), .ZN(new_n461_));
  OR2_X1    g260(.A1(G15gat), .A2(G22gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G15gat), .A2(G22gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G1gat), .A2(G8gat), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n462_), .A2(new_n463_), .B1(KEYINPUT14), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n461_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n459_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT75), .ZN(new_n468_));
  INV_X1    g267(.A(new_n466_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n458_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G229gat), .A2(G233gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n466_), .B(new_n458_), .Z(new_n473_));
  INV_X1    g272(.A(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G113gat), .B(G141gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT76), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G169gat), .B(G197gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n480_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n472_), .A2(new_n475_), .A3(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n455_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT65), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT65), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT6), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n496_));
  INV_X1    g295(.A(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G85gat), .ZN(new_n500_));
  INV_X1    g299(.A(G92gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G85gat), .A2(G92gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(KEYINPUT9), .A3(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(KEYINPUT9), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n499_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT66), .B1(new_n495_), .B2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n499_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n487_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n491_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT66), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n508_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n493_), .A2(new_n519_), .A3(new_n494_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n502_), .A2(new_n503_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n524_), .A2(new_n525_), .A3(KEYINPUT68), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT68), .ZN(new_n527_));
  INV_X1    g326(.A(new_n523_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT7), .ZN(new_n529_));
  INV_X1    g328(.A(G99gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n497_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n516_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n509_), .A2(new_n510_), .A3(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n528_), .B1(new_n533_), .B2(new_n521_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n527_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n515_), .B1(new_n526_), .B2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n539_));
  XOR2_X1   g338(.A(G71gat), .B(G78gat), .Z(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n538_), .A2(KEYINPUT11), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n540_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT12), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n537_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT64), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n534_), .A2(new_n535_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n515_), .A2(new_n551_), .A3(new_n544_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT12), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n514_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(new_n544_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n548_), .A2(new_n550_), .A3(new_n552_), .A4(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n550_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n513_), .B(new_n507_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n558_), .A2(new_n545_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n544_), .B1(new_n515_), .B2(new_n551_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n557_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT69), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT71), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n562_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT13), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n562_), .A2(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n562_), .A2(new_n570_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(KEYINPUT13), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT72), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n544_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n469_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT74), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G127gat), .B(G155gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT16), .ZN(new_n584_));
  XOR2_X1   g383(.A(G183gat), .B(G211gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT17), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n582_), .B(new_n588_), .ZN(new_n589_));
  OR3_X1    g388(.A1(new_n581_), .A2(KEYINPUT17), .A3(new_n587_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n537_), .A2(new_n459_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT35), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n554_), .A2(new_n458_), .B1(new_n596_), .B2(new_n595_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n592_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n592_), .B2(new_n599_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(KEYINPUT36), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n605_), .B(KEYINPUT36), .Z(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT37), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(KEYINPUT37), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n485_), .A2(new_n578_), .A3(new_n591_), .A4(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n331_), .A2(KEYINPUT101), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n331_), .A2(KEYINPUT101), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n614_), .A2(G1gat), .A3(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n610_), .A2(KEYINPUT103), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n455_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n481_), .A2(new_n483_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n577_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n591_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n331_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n618_), .A2(new_n619_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n620_), .A2(new_n632_), .A3(new_n633_), .ZN(G1324gat));
  OR2_X1    g433(.A1(new_n417_), .A2(new_n423_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n409_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n626_), .A2(new_n636_), .A3(new_n630_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n637_), .A2(new_n638_), .A3(G8gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n637_), .B2(G8gat), .ZN(new_n640_));
  INV_X1    g439(.A(new_n636_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(G8gat), .ZN(new_n642_));
  OAI22_X1  g441(.A1(new_n639_), .A2(new_n640_), .B1(new_n614_), .B2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g443(.A(G15gat), .B1(new_n631_), .B2(new_n454_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT41), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n614_), .A2(G15gat), .A3(new_n454_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1326gat));
  OAI21_X1  g447(.A(G22gat), .B1(new_n631_), .B2(new_n373_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT42), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n373_), .A2(G22gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(new_n614_), .B2(new_n651_), .ZN(G1327gat));
  INV_X1    g451(.A(new_n577_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(new_n624_), .A3(new_n591_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n485_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n434_), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT43), .B1(new_n455_), .B2(new_n613_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  INV_X1    g458(.A(new_n613_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n454_), .ZN(new_n661_));
  AOI22_X1  g460(.A1(new_n429_), .A2(new_n428_), .B1(new_n450_), .B2(new_n373_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n662_), .B2(new_n452_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n659_), .B(new_n660_), .C1(new_n663_), .C2(new_n425_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n658_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n628_), .A2(new_n591_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(KEYINPUT44), .A3(new_n666_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n617_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(G29gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n657_), .B1(new_n673_), .B2(new_n675_), .ZN(G1328gat));
  NAND3_X1  g475(.A1(new_n669_), .A2(new_n636_), .A3(new_n671_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n641_), .A2(G36gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n655_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n678_), .A2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(KEYINPUT46), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1329gat));
  XOR2_X1   g485(.A(KEYINPUT105), .B(G43gat), .Z(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(new_n655_), .B2(new_n454_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT106), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n669_), .A2(G43gat), .A3(new_n661_), .A4(new_n671_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g491(.A1(new_n670_), .A2(new_n373_), .A3(new_n672_), .ZN(new_n693_));
  INV_X1    g492(.A(G50gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n372_), .A2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT107), .Z(new_n696_));
  OAI22_X1  g495(.A1(new_n693_), .A2(new_n694_), .B1(new_n655_), .B2(new_n696_), .ZN(G1331gat));
  NAND2_X1  g496(.A1(new_n591_), .A2(new_n484_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n578_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n626_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(G57gat), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n331_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n455_), .A2(new_n627_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n660_), .A2(new_n577_), .A3(new_n629_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(KEYINPUT108), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n674_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n702_), .B1(new_n709_), .B2(new_n701_), .ZN(G1332gat));
  OAI21_X1  g509(.A(G64gat), .B1(new_n700_), .B2(new_n641_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT48), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n641_), .A2(G64gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n705_), .B2(new_n713_), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n700_), .B2(new_n454_), .ZN(new_n715_));
  XOR2_X1   g514(.A(KEYINPUT109), .B(KEYINPUT49), .Z(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n454_), .A2(G71gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n705_), .B2(new_n718_), .ZN(G1334gat));
  OR3_X1    g518(.A1(new_n705_), .A2(G78gat), .A3(new_n373_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n626_), .A2(new_n372_), .A3(new_n699_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(G78gat), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n722_), .A2(new_n723_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n720_), .B1(new_n724_), .B2(new_n725_), .ZN(G1335gat));
  NAND3_X1  g525(.A1(new_n653_), .A2(new_n484_), .A3(new_n629_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n658_), .B2(new_n664_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n331_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n578_), .A2(new_n591_), .A3(new_n624_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n703_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n674_), .A2(new_n500_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n730_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT111), .Z(G1336gat));
  OAI21_X1  g534(.A(G92gat), .B1(new_n729_), .B2(new_n641_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n732_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n501_), .A3(new_n636_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1337gat));
  OAI21_X1  g538(.A(G99gat), .B1(new_n729_), .B2(new_n454_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n661_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n740_), .B(KEYINPUT112), .C1(new_n732_), .C2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g543(.A1(new_n737_), .A2(new_n497_), .A3(new_n372_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n373_), .B(new_n727_), .C1(new_n658_), .C2(new_n664_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n497_), .B1(new_n747_), .B2(KEYINPUT113), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT113), .B1(new_n728_), .B2(new_n372_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n746_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n727_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n665_), .A2(KEYINPUT113), .A3(new_n372_), .A4(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G106gat), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n754_), .A2(new_n749_), .A3(KEYINPUT52), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n745_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n745_), .C1(new_n751_), .C2(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1339gat));
  AOI21_X1  g559(.A(new_n698_), .B1(new_n576_), .B2(new_n573_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n613_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(new_n613_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n562_), .A2(new_n568_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n627_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n556_), .A2(KEYINPUT114), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT114), .B1(new_n556_), .B2(new_n769_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT12), .B1(new_n558_), .B2(new_n545_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n559_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n773_), .A2(new_n548_), .A3(KEYINPUT55), .A4(new_n550_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n552_), .B1(new_n560_), .B2(KEYINPUT12), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT68), .B1(new_n524_), .B2(new_n525_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n534_), .A2(new_n527_), .A3(new_n535_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n546_), .B1(new_n778_), .B2(new_n515_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n557_), .B1(new_n775_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n774_), .A2(new_n780_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n770_), .A2(new_n771_), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n768_), .B1(new_n782_), .B2(new_n568_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n781_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n775_), .A2(new_n779_), .A3(new_n557_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(KEYINPUT55), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n556_), .A2(KEYINPUT114), .A3(new_n769_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n567_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n767_), .B1(new_n783_), .B2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n468_), .A2(new_n470_), .A3(new_n474_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n482_), .B1(new_n473_), .B2(new_n471_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n483_), .A2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n571_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n624_), .B1(new_n791_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n795_), .B1(new_n562_), .B2(new_n568_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n567_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n567_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT58), .B(new_n800_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n660_), .A3(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n624_), .B(KEYINPUT57), .C1(new_n791_), .C2(new_n796_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n799_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n765_), .B1(new_n809_), .B2(new_n629_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n454_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n424_), .A2(new_n617_), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n812_), .A3(new_n814_), .ZN(new_n815_));
  NOR4_X1   g614(.A1(new_n810_), .A2(new_n454_), .A3(new_n424_), .A4(new_n617_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G113gat), .B1(new_n818_), .B2(new_n484_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n811_), .A2(new_n812_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n816_), .A2(KEYINPUT115), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(G113gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n627_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n819_), .B1(new_n824_), .B2(new_n826_), .ZN(G1340gat));
  OAI21_X1  g626(.A(G120gat), .B1(new_n818_), .B2(new_n578_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n577_), .A2(KEYINPUT60), .ZN(new_n829_));
  INV_X1    g628(.A(G120gat), .ZN(new_n830_));
  MUX2_X1   g629(.A(KEYINPUT60), .B(new_n829_), .S(new_n830_), .Z(new_n831_));
  NAND3_X1  g630(.A1(new_n822_), .A2(new_n823_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n828_), .A2(KEYINPUT117), .A3(new_n832_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n818_), .A2(new_n838_), .A3(new_n629_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n824_), .B2(new_n629_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT118), .B(new_n838_), .C1(new_n824_), .C2(new_n629_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n839_), .B1(new_n842_), .B2(new_n843_), .ZN(G1342gat));
  XOR2_X1   g643(.A(KEYINPUT119), .B(G134gat), .Z(new_n845_));
  NOR3_X1   g644(.A1(new_n818_), .A2(new_n613_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(G134gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n822_), .A2(new_n823_), .A3(new_n625_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(G1343gat));
  NOR2_X1   g648(.A1(new_n810_), .A2(new_n661_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n636_), .A2(new_n373_), .A3(new_n617_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n484_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n294_), .ZN(G1344gat));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n578_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n295_), .ZN(G1345gat));
  INV_X1    g655(.A(new_n852_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(KEYINPUT120), .A3(new_n591_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n852_), .B2(new_n629_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1346gat));
  OR3_X1    g662(.A1(new_n852_), .A2(G162gat), .A3(new_n624_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G162gat), .B1(new_n852_), .B2(new_n613_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n484_), .A2(new_n374_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n636_), .A2(new_n373_), .A3(new_n617_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n810_), .A2(new_n454_), .A3(new_n868_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n869_), .A2(KEYINPUT123), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(KEYINPUT123), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n867_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n810_), .A2(new_n454_), .A3(new_n484_), .A4(new_n868_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n208_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n873_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n876_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n874_), .B2(new_n208_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n809_), .A2(new_n629_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n765_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n868_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n882_), .A2(new_n661_), .A3(new_n627_), .A4(new_n883_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n884_), .A2(new_n873_), .A3(G169gat), .A4(new_n876_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n879_), .A2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n872_), .B1(new_n877_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT124), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n872_), .B(new_n889_), .C1(new_n877_), .C2(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1348gat));
  INV_X1    g690(.A(new_n869_), .ZN(new_n892_));
  OAI21_X1  g691(.A(G176gat), .B1(new_n892_), .B2(new_n578_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n870_), .A2(new_n871_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n653_), .A2(new_n226_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  AOI21_X1  g695(.A(G183gat), .B1(new_n869_), .B2(new_n591_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n894_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n629_), .A2(new_n217_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n894_), .B2(new_n613_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n625_), .A2(new_n216_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n894_), .B2(new_n902_), .ZN(G1351gat));
  INV_X1    g702(.A(new_n426_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n850_), .A2(new_n904_), .A3(new_n636_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n907_), .A2(G197gat), .A3(new_n627_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G197gat), .B1(new_n907_), .B2(new_n627_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1352gat));
  XNOR2_X1  g709(.A(new_n905_), .B(KEYINPUT125), .ZN(new_n911_));
  OR3_X1    g710(.A1(new_n911_), .A2(G204gat), .A3(new_n578_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G204gat), .B1(new_n911_), .B2(new_n578_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1353gat));
  NAND2_X1  g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n591_), .A2(new_n915_), .ZN(new_n916_));
  XOR2_X1   g715(.A(new_n916_), .B(KEYINPUT126), .Z(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(KEYINPUT127), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n907_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n918_), .A2(KEYINPUT127), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n907_), .B(new_n919_), .C1(KEYINPUT127), .C2(new_n918_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1354gat));
  OAI21_X1  g723(.A(G218gat), .B1(new_n911_), .B2(new_n613_), .ZN(new_n925_));
  INV_X1    g724(.A(G218gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n907_), .A2(new_n926_), .A3(new_n625_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1355gat));
endmodule


