//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT88), .B(G197gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(new_n206_), .B2(G204gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT21), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT89), .B1(new_n205_), .B2(G204gat), .ZN(new_n212_));
  INV_X1    g011(.A(G204gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n212_), .B1(G197gat), .B2(new_n213_), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n205_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT21), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n209_), .A2(KEYINPUT90), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n219_), .B1(new_n209_), .B2(KEYINPUT90), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n207_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT91), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n207_), .A2(new_n218_), .A3(KEYINPUT91), .A4(new_n220_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n217_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G155gat), .B(G162gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT86), .ZN(new_n229_));
  NOR3_X1   g028(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n227_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G141gat), .A2(G148gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(G141gat), .A2(G148gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G155gat), .A2(G162gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(KEYINPUT1), .B2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(KEYINPUT1), .ZN(new_n240_));
  AOI211_X1 g039(.A(new_n235_), .B(new_n236_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT29), .B1(new_n234_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n226_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G228gat), .ZN(new_n244_));
  INV_X1    g043(.A(G233gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n226_), .B(new_n242_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n203_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n234_), .A2(new_n241_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT29), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT28), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n254_), .A3(new_n251_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G22gat), .B(G50gat), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n253_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n249_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n247_), .A2(new_n248_), .A3(new_n203_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT92), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT92), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT87), .ZN(new_n266_));
  OR3_X1    g065(.A1(new_n257_), .A2(new_n258_), .A3(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n267_), .B(new_n268_), .C1(new_n261_), .C2(new_n249_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(G15gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT30), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT31), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G183gat), .ZN(new_n278_));
  INV_X1    g077(.A(G190gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT23), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT84), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(G183gat), .A3(G190gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT85), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(G183gat), .B2(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(KEYINPUT22), .B(G169gat), .Z(new_n290_));
  OAI21_X1  g089(.A(new_n289_), .B1(G176gat), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n286_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n280_), .A2(new_n283_), .A3(KEYINPUT82), .ZN(new_n294_));
  INV_X1    g093(.A(G169gat), .ZN(new_n295_));
  INV_X1    g094(.A(G176gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n299_), .A2(new_n282_), .A3(G183gat), .A4(G190gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n294_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT83), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT25), .B(G183gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT26), .B(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(KEYINPUT80), .A2(new_n306_), .B1(new_n289_), .B2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n294_), .A2(new_n298_), .A3(KEYINPUT83), .A4(new_n300_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n306_), .A2(KEYINPUT80), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n303_), .A2(new_n309_), .A3(new_n310_), .A4(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n293_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G71gat), .B(G99gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G43gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n313_), .B(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G127gat), .B(G134gat), .Z(new_n317_));
  XOR2_X1   g116(.A(G113gat), .B(G120gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n316_), .A2(new_n319_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n277_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n313_), .B(new_n315_), .Z(new_n324_));
  XOR2_X1   g123(.A(new_n317_), .B(new_n318_), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(new_n276_), .A3(new_n320_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n250_), .A2(new_n319_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n325_), .B1(new_n234_), .B2(new_n241_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n250_), .A2(new_n319_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT97), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT97), .B1(new_n330_), .B2(KEYINPUT4), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n329_), .A2(new_n330_), .A3(KEYINPUT4), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n335_), .B1(new_n342_), .B2(new_n334_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT0), .B(G57gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n343_), .B(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n328_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT19), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n353_));
  NAND2_X1  g152(.A1(new_n297_), .A2(new_n287_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n305_), .B(KEYINPUT93), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n304_), .B2(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n294_), .B(new_n300_), .C1(G183gat), .C2(G190gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT95), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n291_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n359_), .A2(new_n285_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n216_), .A2(new_n211_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT20), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n226_), .A2(new_n313_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n352_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n352_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n226_), .A2(new_n313_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G8gat), .B(G36gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n368_), .A2(new_n379_), .A3(new_n373_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT99), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n370_), .A2(new_n372_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n352_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n359_), .A2(new_n285_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n362_), .A2(new_n363_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n369_), .B1(new_n391_), .B2(new_n226_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n365_), .A2(new_n293_), .A3(new_n312_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n371_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n386_), .B1(new_n388_), .B2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n371_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(KEYINPUT99), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n380_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT27), .A3(new_n382_), .ZN(new_n399_));
  AND4_X1   g198(.A1(new_n271_), .A2(new_n350_), .A3(new_n385_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n379_), .A2(KEYINPUT32), .ZN(new_n401_));
  INV_X1    g200(.A(new_n397_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n366_), .A2(new_n367_), .A3(new_n352_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT99), .B1(new_n403_), .B2(new_n396_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n343_), .A2(new_n348_), .ZN(new_n406_));
  AOI211_X1 g205(.A(new_n347_), .B(new_n335_), .C1(new_n342_), .C2(new_n334_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n401_), .ZN(new_n408_));
  OAI22_X1  g207(.A1(new_n406_), .A2(new_n407_), .B1(new_n408_), .B2(new_n374_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n342_), .A2(new_n334_), .ZN(new_n410_));
  OAI211_X1 g209(.A(KEYINPUT33), .B(new_n347_), .C1(new_n410_), .C2(new_n335_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT98), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n333_), .B1(new_n332_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n331_), .A2(KEYINPUT98), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n347_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n342_), .A2(new_n334_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n412_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n411_), .B1(new_n418_), .B2(new_n406_), .ZN(new_n419_));
  OAI22_X1  g218(.A1(new_n405_), .A2(new_n409_), .B1(new_n419_), .B2(new_n383_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n271_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n349_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n399_), .A2(new_n422_), .A3(new_n270_), .A4(new_n385_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n400_), .B1(new_n424_), .B2(new_n328_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT13), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT64), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT64), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT6), .ZN(new_n430_));
  AND2_X1   g229(.A1(G99gat), .A2(G106gat), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT7), .ZN(new_n434_));
  INV_X1    g233(.A(G99gat), .ZN(new_n435_));
  INV_X1    g234(.A(G106gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n432_), .A2(new_n433_), .A3(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G85gat), .B(G92gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT65), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n429_), .A2(KEYINPUT6), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n427_), .A2(KEYINPUT64), .ZN(new_n444_));
  OAI22_X1  g243(.A1(new_n443_), .A2(new_n444_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n438_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT65), .ZN(new_n451_));
  INV_X1    g250(.A(new_n441_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n442_), .A2(KEYINPUT8), .A3(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n436_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT9), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(G85gat), .A3(G92gat), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n457_), .B(new_n459_), .C1(new_n458_), .C2(new_n441_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n445_), .A2(new_n449_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n451_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT8), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G57gat), .B(G64gat), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n466_), .A2(KEYINPUT11), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(KEYINPUT11), .ZN(new_n468_));
  XOR2_X1   g267(.A(G71gat), .B(G78gat), .Z(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n468_), .A2(new_n469_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n454_), .A2(new_n465_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G230gat), .A2(G233gat), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n454_), .B2(new_n465_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI211_X1 g281(.A(new_n472_), .B(new_n482_), .C1(new_n454_), .C2(new_n465_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n475_), .B(new_n476_), .C1(new_n479_), .C2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n473_), .ZN(new_n485_));
  OAI211_X1 g284(.A(G230gat), .B(G233gat), .C1(new_n485_), .C2(new_n477_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G120gat), .B(G148gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT5), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G176gat), .B(G204gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n484_), .A2(new_n486_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n426_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n484_), .A2(new_n486_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n490_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n484_), .A2(new_n486_), .A3(new_n491_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(KEYINPUT13), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G36gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G29gat), .ZN(new_n501_));
  INV_X1    g300(.A(G29gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G36gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G50gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G43gat), .ZN(new_n506_));
  INV_X1    g305(.A(G43gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G50gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n501_), .A2(new_n503_), .A3(new_n506_), .A4(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G1gat), .ZN(new_n513_));
  INV_X1    g312(.A(G8gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G1gat), .A2(G8gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AND2_X1   g316(.A1(G15gat), .A2(G22gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(G15gat), .A2(G22gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT14), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(G1gat), .B2(G8gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n517_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n524_), .A2(new_n521_), .A3(new_n516_), .A4(new_n515_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n512_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n504_), .A2(new_n509_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n501_), .A2(new_n503_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n523_), .B(new_n525_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT75), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT76), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n527_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n531_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT76), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n526_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n535_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT15), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n512_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n523_), .A2(new_n525_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n540_), .B(KEYINPUT77), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n530_), .A3(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G169gat), .B(G197gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  NAND3_X1  g351(.A1(new_n542_), .A2(new_n549_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT78), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n552_), .B1(new_n542_), .B2(new_n549_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n542_), .A2(new_n549_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT78), .ZN(new_n558_));
  INV_X1    g357(.A(new_n552_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT79), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n556_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n557_), .A2(new_n559_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(KEYINPUT78), .A3(new_n553_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT79), .B1(new_n565_), .B2(new_n560_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n425_), .A2(new_n499_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n454_), .A2(new_n465_), .A3(new_n512_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT35), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n454_), .A2(new_n465_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(new_n545_), .ZN(new_n578_));
  AOI211_X1 g377(.A(KEYINPUT68), .B(new_n544_), .C1(new_n454_), .C2(new_n465_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n575_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  AOI211_X1 g379(.A(new_n573_), .B(new_n572_), .C1(new_n569_), .C2(KEYINPUT69), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n572_), .A2(new_n573_), .ZN(new_n583_));
  OAI221_X1 g382(.A(new_n575_), .B1(KEYINPUT69), .B2(new_n583_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n582_), .A2(new_n584_), .A3(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n587_), .B(KEYINPUT36), .Z(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT71), .Z(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n590_), .B1(new_n593_), .B2(KEYINPUT72), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT72), .ZN(new_n595_));
  AOI211_X1 g394(.A(new_n595_), .B(new_n592_), .C1(new_n582_), .C2(new_n584_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT37), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT73), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n582_), .A2(new_n584_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n591_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT37), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n590_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n597_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n598_), .B1(new_n597_), .B2(new_n602_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n472_), .B(new_n546_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G183gat), .B(G211gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT17), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n608_), .A2(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n613_), .A2(KEYINPUT17), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n608_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n605_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n568_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n513_), .A3(new_n349_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n494_), .A2(new_n498_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n556_), .A2(new_n561_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT100), .Z(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(new_n618_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n600_), .A2(new_n590_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n425_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n634_), .B2(new_n422_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n622_), .A2(new_n623_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n624_), .A2(new_n635_), .A3(new_n636_), .ZN(G1324gat));
  AND2_X1   g436(.A1(new_n399_), .A2(new_n385_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n633_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT101), .B1(new_n640_), .B2(G8gat), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n514_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n643_), .B1(new_n620_), .B2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(KEYINPUT101), .A3(G8gat), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n641_), .A2(new_n642_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g448(.A(new_n328_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n273_), .B1(new_n633_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT102), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(KEYINPUT41), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(KEYINPUT41), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n621_), .A2(new_n273_), .A3(new_n650_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(G1326gat));
  INV_X1    g455(.A(G22gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n633_), .B2(new_n270_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT42), .Z(new_n659_));
  NAND3_X1  g458(.A1(new_n621_), .A2(new_n657_), .A3(new_n270_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT103), .ZN(G1327gat));
  INV_X1    g461(.A(new_n618_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n630_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n568_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n666_), .B2(new_n349_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n628_), .A2(new_n663_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n424_), .A2(new_n328_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n400_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT43), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT105), .B1(new_n673_), .B2(new_n605_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n597_), .A2(new_n602_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT73), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n597_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n679_));
  NOR4_X1   g478(.A1(new_n425_), .A2(new_n678_), .A3(new_n679_), .A4(KEYINPUT43), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n674_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n605_), .A2(KEYINPUT104), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n678_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n685_), .B2(new_n425_), .ZN(new_n686_));
  AOI211_X1 g485(.A(new_n668_), .B(new_n670_), .C1(new_n681_), .C2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n681_), .A2(new_n686_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n669_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(KEYINPUT106), .A3(new_n668_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n670_), .B1(new_n681_), .B2(new_n686_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(KEYINPUT44), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n687_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n422_), .A2(new_n502_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n667_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n500_), .B1(new_n694_), .B2(new_n639_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n665_), .A2(G36gat), .A3(new_n638_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT45), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n700_), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n638_), .B(new_n687_), .C1(new_n690_), .C2(new_n693_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT46), .B(new_n702_), .C1(new_n703_), .C2(new_n500_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1329gat));
  XOR2_X1   g504(.A(KEYINPUT107), .B(G43gat), .Z(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n666_), .B2(new_n650_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n328_), .A2(new_n507_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n694_), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n710_), .ZN(new_n712_));
  AOI211_X1 g511(.A(new_n707_), .B(new_n712_), .C1(new_n694_), .C2(new_n708_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1330gat));
  AOI21_X1  g513(.A(G50gat), .B1(new_n666_), .B2(new_n270_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n271_), .A2(new_n505_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n694_), .B2(new_n716_), .ZN(G1331gat));
  NOR3_X1   g516(.A1(new_n425_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(new_n619_), .ZN(new_n719_));
  INV_X1    g518(.A(G57gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n349_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n563_), .A2(new_n566_), .A3(new_n618_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n632_), .A2(new_n499_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G57gat), .B1(new_n723_), .B2(new_n422_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1332gat));
  OAI21_X1  g524(.A(G64gat), .B1(new_n723_), .B2(new_n638_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT48), .ZN(new_n727_));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n719_), .A2(new_n728_), .A3(new_n639_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1333gat));
  OAI21_X1  g529(.A(G71gat), .B1(new_n723_), .B2(new_n328_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT49), .ZN(new_n732_));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n719_), .A2(new_n733_), .A3(new_n650_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1334gat));
  OAI21_X1  g534(.A(G78gat), .B1(new_n723_), .B2(new_n271_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT50), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n271_), .A2(G78gat), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT109), .Z(new_n739_));
  NAND2_X1  g538(.A1(new_n719_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(G1335gat));
  OAI211_X1 g540(.A(new_n499_), .B(new_n618_), .C1(new_n561_), .C2(new_n556_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n681_), .B2(new_n686_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(new_n349_), .ZN(new_n744_));
  INV_X1    g543(.A(G85gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n718_), .A2(new_n664_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n349_), .A2(new_n745_), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n744_), .A2(new_n745_), .B1(new_n746_), .B2(new_n747_), .ZN(G1336gat));
  INV_X1    g547(.A(G92gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n746_), .B2(new_n638_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT110), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n638_), .A2(new_n749_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n743_), .B2(new_n752_), .ZN(G1337gat));
  NAND2_X1  g552(.A1(new_n455_), .A2(new_n456_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n746_), .A2(new_n754_), .A3(new_n328_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n743_), .A2(new_n650_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G99gat), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(G1338gat));
  NAND4_X1  g558(.A1(new_n718_), .A2(new_n436_), .A3(new_n270_), .A4(new_n664_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n743_), .A2(new_n270_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(G106gat), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT52), .B(new_n436_), .C1(new_n743_), .C2(new_n270_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n765_), .B(new_n766_), .Z(G1339gat));
  NOR2_X1   g566(.A1(new_n639_), .A2(new_n270_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n349_), .A3(new_n650_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n484_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n475_), .B1(new_n479_), .B2(new_n483_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(G230gat), .A3(G233gat), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n773_), .B1(new_n484_), .B2(new_n772_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT56), .B(new_n490_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n484_), .A2(new_n772_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT55), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n776_), .A3(new_n774_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n784_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n490_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n781_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n490_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n788_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n786_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n530_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(new_n548_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n552_), .B1(new_n547_), .B2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n535_), .A2(new_n539_), .A3(new_n548_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n553_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n497_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n771_), .B1(new_n792_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n799_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n791_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT58), .B(new_n801_), .C1(new_n804_), .C2(new_n786_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n800_), .A2(new_n605_), .A3(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n798_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n626_), .A2(new_n497_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n787_), .A2(new_n789_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n779_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n807_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  AOI211_X1 g611(.A(KEYINPUT115), .B(new_n808_), .C1(new_n809_), .C2(new_n779_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n630_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT57), .B(new_n630_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n806_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n618_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n625_), .A2(new_n722_), .A3(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n562_), .B1(new_n556_), .B2(new_n561_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n565_), .A2(KEYINPUT79), .A3(new_n560_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n663_), .A3(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT113), .B1(new_n499_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n820_), .B1(new_n678_), .B2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n827_), .B(new_n820_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT118), .B1(new_n819_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n834_), .B(new_n831_), .C1(new_n818_), .C2(new_n618_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n770_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837_), .B2(new_n626_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(KEYINPUT59), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n831_), .B1(new_n818_), .B2(new_n618_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n769_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n839_), .B1(new_n840_), .B2(new_n845_), .ZN(new_n846_));
  AOI211_X1 g645(.A(KEYINPUT120), .B(new_n844_), .C1(new_n836_), .C2(KEYINPUT59), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n567_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n838_), .B1(new_n848_), .B2(new_n850_), .ZN(G1340gat));
  AOI211_X1 g650(.A(new_n625_), .B(new_n844_), .C1(new_n836_), .C2(KEYINPUT59), .ZN(new_n852_));
  INV_X1    g651(.A(G120gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n625_), .B2(KEYINPUT60), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(KEYINPUT60), .B2(new_n853_), .ZN(new_n855_));
  OAI22_X1  g654(.A1(new_n852_), .A2(new_n853_), .B1(new_n836_), .B2(new_n855_), .ZN(G1341gat));
  AOI21_X1  g655(.A(G127gat), .B1(new_n837_), .B2(new_n663_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n663_), .A2(KEYINPUT121), .A3(G127gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(KEYINPUT121), .B2(G127gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n848_), .B2(new_n859_), .ZN(G1342gat));
  AOI21_X1  g659(.A(G134gat), .B1(new_n837_), .B2(new_n631_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n605_), .A2(G134gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n848_), .B2(new_n862_), .ZN(G1343gat));
  NAND2_X1  g662(.A1(new_n819_), .A2(new_n832_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n834_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n841_), .A2(KEYINPUT118), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NOR4_X1   g666(.A1(new_n639_), .A2(new_n422_), .A3(new_n271_), .A4(new_n650_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n626_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT122), .B(G141gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1344gat));
  NAND2_X1  g671(.A1(new_n869_), .A2(new_n499_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G148gat), .ZN(G1345gat));
  OAI211_X1 g673(.A(new_n663_), .B(new_n868_), .C1(new_n833_), .C2(new_n835_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n875_), .A2(KEYINPUT123), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(KEYINPUT123), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1346gat));
  AOI21_X1  g680(.A(G162gat), .B1(new_n869_), .B2(new_n631_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n682_), .A2(new_n684_), .A3(G162gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n869_), .B2(new_n883_), .ZN(G1347gat));
  NOR3_X1   g683(.A1(new_n638_), .A2(new_n349_), .A3(new_n328_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n271_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n841_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n888_), .A2(new_n290_), .A3(new_n561_), .A4(new_n556_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n295_), .B1(new_n887_), .B2(new_n626_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(KEYINPUT62), .B2(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(KEYINPUT62), .B2(new_n890_), .ZN(G1348gat));
  AOI21_X1  g691(.A(new_n270_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n893_), .A2(G176gat), .A3(new_n499_), .A4(new_n885_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n296_), .B1(new_n888_), .B2(new_n625_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n894_), .A2(new_n895_), .A3(KEYINPUT124), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1349gat));
  NOR3_X1   g699(.A1(new_n888_), .A2(new_n618_), .A3(new_n304_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n893_), .A2(new_n663_), .A3(new_n885_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n278_), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n888_), .B2(new_n678_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n887_), .A2(new_n631_), .A3(new_n358_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1351gat));
  NOR4_X1   g705(.A1(new_n638_), .A2(new_n349_), .A3(new_n271_), .A4(new_n650_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n867_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n626_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n499_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G204gat), .ZN(G1353gat));
  OAI21_X1  g712(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n914_));
  NAND2_X1  g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n663_), .A2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n908_), .B2(new_n916_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT126), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n917_), .B(new_n920_), .ZN(G1354gat));
  AOI21_X1  g720(.A(G218gat), .B1(new_n909_), .B2(new_n631_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n605_), .A2(G218gat), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(KEYINPUT127), .Z(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n909_), .B2(new_n924_), .ZN(G1355gat));
endmodule


