//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n962_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT68), .B(KEYINPUT35), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G29gat), .B(G36gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n208_), .A2(new_n209_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n207_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n208_), .A2(new_n209_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(new_n210_), .A3(new_n206_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(KEYINPUT15), .A3(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT65), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT6), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT6), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(G99gat), .A3(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n222_), .A2(new_n223_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT7), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n221_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n225_), .A2(new_n230_), .A3(new_n232_), .A4(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT8), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(KEYINPUT64), .B(G92gat), .Z(new_n244_));
  INV_X1    g043(.A(G85gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(KEYINPUT9), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n244_), .A2(new_n246_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n237_), .A2(KEYINPUT9), .A3(new_n238_), .ZN(new_n248_));
  OR2_X1    g047(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n223_), .A3(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  NOR4_X1   g052(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n234_), .B1(new_n233_), .B2(new_n221_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n227_), .A2(new_n229_), .B1(new_n231_), .B2(KEYINPUT7), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n239_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n253_), .B1(new_n258_), .B2(KEYINPUT8), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n220_), .B1(new_n243_), .B2(new_n259_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n259_), .A2(new_n216_), .A3(new_n243_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI211_X1 g061(.A(new_n204_), .B(new_n205_), .C1(new_n260_), .C2(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n204_), .A2(new_n205_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n204_), .A2(new_n205_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n260_), .A2(new_n264_), .A3(new_n262_), .A4(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G190gat), .B(G218gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G134gat), .B(G162gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT36), .Z(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  NOR4_X1   g073(.A1(new_n263_), .A2(new_n267_), .A3(KEYINPUT36), .A4(new_n271_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT37), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT37), .B1(new_n274_), .B2(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G8gat), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n281_), .A2(KEYINPUT70), .ZN(new_n282_));
  INV_X1    g081(.A(G15gat), .ZN(new_n283_));
  INV_X1    g082(.A(G22gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G15gat), .A2(G22gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G1gat), .A2(G8gat), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n285_), .A2(new_n286_), .B1(KEYINPUT14), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n281_), .A2(KEYINPUT70), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n282_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n282_), .B2(new_n289_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(G231gat), .A2(G233gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n292_), .B(new_n293_), .Z(new_n294_));
  INV_X1    g093(.A(G64gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G57gat), .ZN(new_n296_));
  INV_X1    g095(.A(G57gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G64gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n298_), .A3(KEYINPUT11), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT66), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G57gat), .B(G64gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(KEYINPUT11), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(new_n298_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT11), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(G71gat), .A2(G78gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(G71gat), .A2(G78gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n300_), .A2(new_n303_), .A3(new_n306_), .A4(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(new_n301_), .B2(KEYINPUT11), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n302_), .B1(new_n301_), .B2(KEYINPUT11), .ZN(new_n312_));
  AND4_X1   g111(.A1(new_n302_), .A2(new_n296_), .A3(new_n298_), .A4(KEYINPUT11), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n294_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G127gat), .B(G155gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G183gat), .B(G211gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT72), .B(KEYINPUT17), .Z(new_n321_));
  NOR3_X1   g120(.A1(new_n315_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n314_), .A2(new_n310_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n294_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n314_), .A2(new_n310_), .A3(KEYINPUT67), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT67), .B1(new_n314_), .B2(new_n310_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT73), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n324_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n320_), .B(KEYINPUT17), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n324_), .A2(new_n329_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n325_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n280_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G230gat), .ZN(new_n337_));
  INV_X1    g136(.A(G233gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n259_), .A2(new_n243_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n328_), .B2(new_n340_), .ZN(new_n341_));
  OAI22_X1  g140(.A1(new_n326_), .A2(new_n327_), .B1(new_n259_), .B2(new_n243_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT12), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT12), .B(new_n323_), .C1(new_n259_), .C2(new_n243_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT67), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n300_), .A2(new_n303_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n314_), .A2(new_n310_), .A3(KEYINPUT67), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n241_), .A2(new_n242_), .B1(new_n252_), .B2(new_n247_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n258_), .A2(KEYINPUT8), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .A4(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n342_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n339_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n346_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G120gat), .B(G148gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT5), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G176gat), .B(G204gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n346_), .A2(new_n356_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT13), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n362_), .A2(KEYINPUT13), .A3(new_n364_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n336_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT74), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n373_));
  OR2_X1    g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT2), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381_));
  INV_X1    g180(.A(G141gat), .ZN(new_n382_));
  INV_X1    g181(.A(G148gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n379_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n376_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT1), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n374_), .A2(new_n390_), .A3(new_n375_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n382_), .A2(new_n383_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n391_), .A2(new_n377_), .A3(new_n392_), .A4(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n388_), .A2(new_n389_), .A3(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n395_), .A2(KEYINPUT28), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(KEYINPUT28), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G22gat), .B(G50gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n396_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n388_), .A2(new_n394_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT28), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(new_n389_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n395_), .A2(KEYINPUT28), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n398_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n373_), .B1(new_n400_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n399_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(new_n404_), .A3(new_n398_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(KEYINPUT79), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n388_), .A2(new_n394_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT29), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT21), .ZN(new_n415_));
  INV_X1    g214(.A(G197gat), .ZN(new_n416_));
  INV_X1    g215(.A(G204gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT80), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT80), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G204gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n416_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G197gat), .A2(G204gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n415_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G218gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G211gat), .ZN(new_n425_));
  INV_X1    g224(.A(G211gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(G218gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n418_), .A2(new_n420_), .A3(new_n416_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n415_), .B1(G197gat), .B2(G204gat), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n423_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n418_), .A2(new_n420_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n422_), .B1(new_n433_), .B2(G197gat), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n415_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G228gat), .A2(G233gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n414_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n389_), .B1(new_n388_), .B2(new_n394_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n423_), .A2(new_n431_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n412_), .B1(new_n439_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT82), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n439_), .A2(new_n443_), .A3(new_n412_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT81), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n439_), .A2(new_n443_), .A3(new_n448_), .A4(new_n412_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n410_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n446_), .A2(KEYINPUT83), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n439_), .A2(new_n443_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n411_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(KEYINPUT83), .A3(new_n411_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n400_), .A2(new_n405_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n372_), .B1(new_n451_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n454_), .A2(KEYINPUT82), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n444_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n460_), .A2(new_n462_), .A3(new_n447_), .A4(new_n449_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n406_), .A2(new_n409_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT84), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n459_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G8gat), .B(G36gat), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n470_), .B(KEYINPUT88), .ZN(new_n475_));
  INV_X1    g274(.A(new_n473_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n474_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G226gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT19), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G183gat), .A2(G190gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT23), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n489_));
  INV_X1    g288(.A(G169gat), .ZN(new_n490_));
  INV_X1    g289(.A(G176gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n488_), .B(new_n489_), .C1(new_n492_), .C2(KEYINPUT24), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT24), .B1(new_n490_), .B2(new_n491_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT26), .B(G190gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT75), .ZN(new_n499_));
  INV_X1    g298(.A(G183gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT25), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n500_), .A2(KEYINPUT25), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n498_), .B(new_n501_), .C1(new_n502_), .C2(new_n499_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n488_), .A2(new_n489_), .ZN(new_n504_));
  OR2_X1    g303(.A1(G183gat), .A2(G190gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT22), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n508_));
  OAI21_X1  g307(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n497_), .A2(new_n503_), .B1(new_n506_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT20), .B1(new_n512_), .B2(new_n442_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT25), .B(G183gat), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n493_), .B1(new_n498_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT85), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n495_), .B1(new_n494_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n517_), .B2(new_n494_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n514_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n442_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n513_), .B1(KEYINPUT86), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT86), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n523_), .A3(new_n442_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n485_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n516_), .A2(new_n519_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n437_), .B1(new_n526_), .B2(new_n514_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n512_), .A2(new_n442_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n527_), .A2(KEYINPUT20), .A3(new_n485_), .A4(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n483_), .B1(new_n525_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n521_), .A2(KEYINPUT86), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT20), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n497_), .A2(new_n503_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n514_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n533_), .B1(new_n536_), .B2(new_n437_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n532_), .A2(new_n524_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n485_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n540_), .A2(new_n480_), .A3(new_n482_), .A4(new_n529_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n531_), .A2(KEYINPUT89), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT27), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n529_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT89), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n483_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n483_), .B(KEYINPUT95), .Z(new_n548_));
  INV_X1    g347(.A(new_n521_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n485_), .B1(new_n549_), .B2(new_n513_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n527_), .A2(KEYINPUT20), .A3(new_n539_), .A4(new_n528_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(KEYINPUT27), .B(new_n531_), .C1(new_n548_), .C2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n547_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n469_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G227gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(new_n283_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G43gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G71gat), .B(G99gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n559_), .A2(new_n561_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT76), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT76), .B1(new_n562_), .B2(new_n563_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n512_), .A2(KEYINPUT30), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n512_), .A2(KEYINPUT30), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n567_), .A3(new_n570_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n564_), .B(new_n565_), .C1(new_n569_), .C2(new_n568_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n572_), .A3(KEYINPUT77), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT31), .ZN(new_n574_));
  XOR2_X1   g373(.A(G127gat), .B(G134gat), .Z(new_n575_));
  XOR2_X1   g374(.A(G113gat), .B(G120gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT31), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n571_), .A2(new_n572_), .A3(KEYINPUT77), .A4(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n574_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n413_), .B(new_n577_), .ZN(new_n584_));
  AND2_X1   g383(.A1(G225gat), .A2(G233gat), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n578_), .A2(new_n413_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n401_), .A2(new_n577_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(KEYINPUT4), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT4), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n578_), .A2(new_n590_), .A3(new_n413_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT90), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT90), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n578_), .A2(new_n593_), .A3(new_n590_), .A4(new_n413_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n586_), .B1(new_n595_), .B2(new_n585_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G1gat), .B(G29gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT91), .B(G85gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT0), .B(G57gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT94), .B1(new_n596_), .B2(new_n601_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n596_), .A2(new_n605_), .A3(new_n601_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n583_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n556_), .A2(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n451_), .A2(new_n372_), .A3(new_n458_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT84), .B1(new_n465_), .B2(new_n466_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n547_), .A2(new_n554_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT96), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n555_), .A2(new_n615_), .A3(new_n468_), .A4(new_n607_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT32), .B1(new_n479_), .B2(new_n481_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT92), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n544_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n617_), .ZN(new_n620_));
  AOI21_X1  g419(.A(KEYINPUT93), .B1(new_n552_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT93), .ZN(new_n622_));
  AOI211_X1 g421(.A(new_n622_), .B(new_n617_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n604_), .A2(new_n619_), .A3(new_n606_), .A4(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n542_), .A2(new_n546_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n627_));
  OR3_X1    g426(.A1(new_n596_), .A2(new_n627_), .A3(new_n601_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n584_), .A2(new_n585_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n601_), .B(new_n629_), .C1(new_n595_), .C2(new_n585_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n627_), .B1(new_n596_), .B2(new_n601_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n625_), .B1(new_n626_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n469_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n614_), .A2(new_n616_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n583_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n609_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G229gat), .A2(G233gat), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n292_), .A2(new_n216_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n215_), .B(new_n213_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n640_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n220_), .B2(new_n292_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n641_), .B1(new_n643_), .B2(new_n638_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G113gat), .B(G141gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G169gat), .B(G197gat), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n645_), .B(new_n646_), .Z(new_n647_));
  XNOR2_X1  g446(.A(new_n644_), .B(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n637_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n371_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT97), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n607_), .A2(G1gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n654_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT97), .B1(new_n651_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n637_), .A2(new_n276_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n369_), .A2(new_n334_), .A3(new_n649_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n607_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n655_), .A2(KEYINPUT38), .A3(new_n657_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n660_), .A2(KEYINPUT98), .A3(new_n664_), .A4(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1324gat));
  OR3_X1    g469(.A1(new_n651_), .A2(G8gat), .A3(new_n555_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G8gat), .B1(new_n663_), .B2(new_n555_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(KEYINPUT39), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(KEYINPUT39), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g475(.A(G15gat), .B1(new_n663_), .B2(new_n636_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n678_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n652_), .A2(new_n283_), .A3(new_n583_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(G1326gat));
  OAI21_X1  g481(.A(G22gat), .B1(new_n663_), .B2(new_n469_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT42), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n652_), .A2(new_n284_), .A3(new_n468_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(new_n276_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(new_n335_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n369_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n637_), .A2(new_n649_), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n607_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G29gat), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n280_), .B(KEYINPUT100), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n637_), .B2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n280_), .A2(KEYINPUT43), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT101), .B1(new_n637_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n468_), .A2(new_n547_), .A3(new_n554_), .A4(new_n607_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n700_), .A2(KEYINPUT96), .B1(new_n633_), .B2(new_n469_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n583_), .B1(new_n701_), .B2(new_n616_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n699_), .B(new_n696_), .C1(new_n702_), .C2(new_n609_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n695_), .A2(new_n698_), .A3(new_n703_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n335_), .A2(new_n649_), .A3(new_n369_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n704_), .A2(KEYINPUT44), .A3(new_n705_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n692_), .A2(G29gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n693_), .B1(new_n712_), .B2(new_n713_), .ZN(G1328gat));
  NOR2_X1   g513(.A1(new_n555_), .A2(G36gat), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n691_), .A2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT45), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n704_), .A2(KEYINPUT44), .A3(new_n705_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n707_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n555_), .ZN(new_n720_));
  INV_X1    g519(.A(G36gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n709_), .A2(new_n613_), .A3(new_n710_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G36gat), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n716_), .A2(KEYINPUT45), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n691_), .B2(new_n715_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT46), .B1(new_n728_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n725_), .B1(new_n727_), .B2(new_n732_), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT104), .B(new_n731_), .C1(new_n726_), .C2(G36gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n724_), .B1(new_n733_), .B2(new_n734_), .ZN(G1329gat));
  AOI21_X1  g534(.A(G43gat), .B1(new_n691_), .B2(new_n583_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT105), .Z(new_n737_));
  NAND2_X1  g536(.A1(new_n583_), .A2(G43gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n711_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g539(.A(G50gat), .B1(new_n691_), .B2(new_n468_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n468_), .A2(G50gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n712_), .B2(new_n742_), .ZN(G1331gat));
  NOR3_X1   g542(.A1(new_n689_), .A2(new_n648_), .A3(new_n334_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n661_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n692_), .A2(G57gat), .ZN(new_n747_));
  OR3_X1    g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n637_), .A2(new_n648_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT106), .B1(new_n637_), .B2(new_n648_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n336_), .A2(new_n689_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(new_n607_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n751_), .B1(G57gat), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT108), .ZN(G1332gat));
  NAND3_X1  g560(.A1(new_n661_), .A2(new_n613_), .A3(new_n744_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G64gat), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n763_), .A2(KEYINPUT109), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(KEYINPUT109), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(KEYINPUT48), .A3(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT48), .B1(new_n764_), .B2(new_n765_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n758_), .A2(G64gat), .A3(new_n555_), .ZN(new_n768_));
  OR3_X1    g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(G1333gat));
  OAI21_X1  g568(.A(G71gat), .B1(new_n745_), .B2(new_n636_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT49), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n636_), .A2(G71gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n758_), .B2(new_n772_), .ZN(G1334gat));
  OAI21_X1  g572(.A(G78gat), .B1(new_n745_), .B2(new_n469_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT50), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n469_), .A2(G78gat), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT110), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n758_), .B2(new_n777_), .ZN(G1335gat));
  AND3_X1   g577(.A1(new_n756_), .A2(new_n369_), .A3(new_n688_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n245_), .A3(new_n692_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n369_), .A2(new_n334_), .A3(new_n649_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT111), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n704_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n607_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n780_), .A2(new_n784_), .ZN(G1336gat));
  AOI21_X1  g584(.A(G92gat), .B1(new_n779_), .B2(new_n613_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n244_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n783_), .A2(new_n555_), .A3(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1337gat));
  AND3_X1   g588(.A1(new_n583_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n779_), .A2(new_n790_), .B1(new_n791_), .B2(KEYINPUT51), .ZN(new_n792_));
  OAI21_X1  g591(.A(G99gat), .B1(new_n783_), .B2(new_n636_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n791_), .A2(KEYINPUT51), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n779_), .A2(new_n223_), .A3(new_n468_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n704_), .A2(new_n468_), .A3(new_n782_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g602(.A1(new_n556_), .A2(new_n607_), .A3(new_n636_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n276_), .A2(new_n806_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n643_), .A2(KEYINPUT116), .ZN(new_n808_));
  INV_X1    g607(.A(new_n638_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n643_), .A2(KEYINPUT116), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n639_), .A2(new_n640_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n647_), .B1(new_n812_), .B2(new_n638_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n811_), .A2(new_n813_), .B1(new_n644_), .B2(new_n647_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n365_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT117), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n817_), .A3(new_n365_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n648_), .A2(new_n364_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n350_), .A2(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n345_), .B1(new_n822_), .B2(KEYINPUT12), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n354_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n821_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n341_), .A2(new_n344_), .A3(KEYINPUT55), .A4(new_n345_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n354_), .B(new_n345_), .C1(new_n822_), .C2(KEYINPUT12), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n339_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n825_), .A2(new_n826_), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(KEYINPUT113), .B2(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n829_), .A2(new_n361_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(KEYINPUT113), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n829_), .B2(new_n361_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n829_), .A2(new_n361_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n830_), .B1(new_n837_), .B2(new_n831_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n820_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n819_), .B1(new_n839_), .B2(KEYINPUT115), .ZN(new_n840_));
  INV_X1    g639(.A(new_n820_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n829_), .A2(new_n361_), .A3(new_n832_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n346_), .A2(new_n821_), .B1(new_n827_), .B2(new_n339_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n363_), .B1(new_n843_), .B2(new_n826_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n844_), .B2(new_n834_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT114), .B1(new_n844_), .B2(KEYINPUT56), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT115), .B(new_n841_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n807_), .B1(new_n840_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n837_), .B2(new_n831_), .ZN(new_n851_));
  AOI211_X1 g650(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n829_), .C2(new_n361_), .ZN(new_n852_));
  OAI22_X1  g651(.A1(new_n851_), .A2(new_n852_), .B1(new_n831_), .B2(new_n837_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n814_), .A2(new_n364_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(KEYINPUT58), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n280_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n853_), .B(new_n854_), .C1(new_n856_), .C2(KEYINPUT58), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n849_), .A2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n841_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n847_), .A3(new_n819_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n866_), .B2(new_n687_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT120), .B1(new_n862_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n280_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n869_), .A2(new_n860_), .B1(new_n866_), .B2(new_n807_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n687_), .B1(new_n840_), .B2(new_n848_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n806_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n868_), .A2(new_n874_), .A3(new_n334_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n280_), .A2(new_n649_), .A3(new_n689_), .A4(new_n335_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT54), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n805_), .B1(new_n875_), .B2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G113gat), .B1(new_n878_), .B2(new_n648_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n863_), .A2(new_n864_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n276_), .B1(new_n880_), .B2(new_n847_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n849_), .B(new_n861_), .C1(new_n881_), .C2(KEYINPUT57), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n877_), .B1(new_n883_), .B2(new_n335_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n804_), .ZN(new_n886_));
  OAI211_X1 g685(.A(KEYINPUT121), .B(new_n886_), .C1(new_n878_), .C2(new_n885_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n877_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n335_), .B1(new_n882_), .B2(KEYINPUT120), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n874_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT59), .B1(new_n891_), .B2(new_n805_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT121), .B1(new_n892_), .B2(new_n886_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n888_), .A2(new_n893_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n648_), .A2(G113gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n879_), .B1(new_n894_), .B2(new_n895_), .ZN(G1340gat));
  INV_X1    g695(.A(G120gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n689_), .B2(KEYINPUT60), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n878_), .B(new_n898_), .C1(KEYINPUT60), .C2(new_n897_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n892_), .A2(new_n369_), .A3(new_n886_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n901_), .B2(new_n897_), .ZN(G1341gat));
  AOI21_X1  g701(.A(G127gat), .B1(new_n878_), .B2(new_n335_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n335_), .A2(G127gat), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n894_), .B2(new_n905_), .ZN(G1342gat));
  AOI21_X1  g705(.A(G134gat), .B1(new_n878_), .B2(new_n276_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n859_), .A2(G134gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n894_), .B2(new_n908_), .ZN(G1343gat));
  NAND2_X1  g708(.A1(new_n875_), .A2(new_n877_), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n469_), .A2(new_n583_), .A3(new_n613_), .A4(new_n607_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n649_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT122), .B(G141gat), .Z(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1344gat));
  NOR2_X1   g714(.A1(new_n912_), .A2(new_n689_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n383_), .ZN(G1345gat));
  NOR2_X1   g716(.A1(new_n912_), .A2(new_n334_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT61), .B(G155gat), .Z(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1346gat));
  AND2_X1   g719(.A1(new_n910_), .A2(new_n911_), .ZN(new_n921_));
  AOI21_X1  g720(.A(G162gat), .B1(new_n921_), .B2(new_n276_), .ZN(new_n922_));
  INV_X1    g721(.A(G162gat), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n912_), .A2(new_n923_), .A3(new_n694_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT123), .B1(new_n922_), .B2(new_n924_), .ZN(new_n925_));
  OR3_X1    g724(.A1(new_n912_), .A2(new_n923_), .A3(new_n694_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n923_), .B1(new_n912_), .B2(new_n687_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n929_), .ZN(G1347gat));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n608_), .A2(new_n555_), .A3(new_n468_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n884_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n648_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n931_), .B1(new_n935_), .B2(G169gat), .ZN(new_n936_));
  AOI211_X1 g735(.A(KEYINPUT62), .B(new_n490_), .C1(new_n934_), .C2(new_n648_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT22), .B(G169gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n648_), .A2(new_n938_), .ZN(new_n939_));
  XOR2_X1   g738(.A(new_n939_), .B(KEYINPUT124), .Z(new_n940_));
  OAI22_X1  g739(.A1(new_n936_), .A2(new_n937_), .B1(new_n933_), .B2(new_n940_), .ZN(G1348gat));
  AND2_X1   g740(.A1(new_n910_), .A2(new_n932_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n689_), .A2(new_n491_), .ZN(new_n943_));
  AND3_X1   g742(.A1(new_n942_), .A2(KEYINPUT125), .A3(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(KEYINPUT125), .B1(new_n942_), .B2(new_n943_), .ZN(new_n945_));
  AOI21_X1  g744(.A(G176gat), .B1(new_n934_), .B2(new_n369_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n944_), .A2(new_n945_), .A3(new_n946_), .ZN(G1349gat));
  AOI21_X1  g746(.A(G183gat), .B1(new_n942_), .B2(new_n335_), .ZN(new_n948_));
  OR2_X1    g747(.A1(new_n334_), .A2(new_n515_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n949_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n884_), .A2(new_n932_), .A3(new_n950_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(KEYINPUT126), .ZN(new_n952_));
  OAI21_X1  g751(.A(KEYINPUT127), .B1(new_n948_), .B2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n910_), .A2(new_n932_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n500_), .B1(new_n954_), .B2(new_n334_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n951_), .A2(KEYINPUT126), .ZN(new_n957_));
  OR2_X1    g756(.A1(new_n951_), .A2(KEYINPUT126), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n955_), .A2(new_n956_), .A3(new_n957_), .A4(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n953_), .A2(new_n959_), .ZN(G1350gat));
  OAI21_X1  g759(.A(G190gat), .B1(new_n933_), .B2(new_n280_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n276_), .A2(new_n498_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n933_), .B2(new_n962_), .ZN(G1351gat));
  NOR4_X1   g762(.A1(new_n891_), .A2(new_n555_), .A3(new_n583_), .A4(new_n612_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(new_n648_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g765(.A(G204gat), .B1(new_n964_), .B2(new_n369_), .ZN(new_n967_));
  AND2_X1   g766(.A1(new_n964_), .A2(new_n369_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n967_), .B1(new_n433_), .B2(new_n968_), .ZN(G1353gat));
  OR2_X1    g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n970_), .B1(new_n964_), .B2(new_n335_), .ZN(new_n971_));
  AND2_X1   g770(.A1(new_n964_), .A2(new_n335_), .ZN(new_n972_));
  XOR2_X1   g771(.A(KEYINPUT63), .B(G211gat), .Z(new_n973_));
  AOI21_X1  g772(.A(new_n971_), .B1(new_n972_), .B2(new_n973_), .ZN(G1354gat));
  NAND3_X1  g773(.A1(new_n964_), .A2(new_n424_), .A3(new_n276_), .ZN(new_n975_));
  AND2_X1   g774(.A1(new_n964_), .A2(new_n859_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n975_), .B1(new_n976_), .B2(new_n424_), .ZN(G1355gat));
endmodule


