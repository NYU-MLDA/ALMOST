//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_;
  XNOR2_X1  g000(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G155gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G183gat), .B(G211gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT76), .B(G127gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT78), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT73), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213_));
  INV_X1    g012(.A(G1gat), .ZN(new_n214_));
  INV_X1    g013(.A(G8gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n211_), .A2(KEYINPUT73), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n211_), .A2(KEYINPUT73), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n219_), .A2(new_n216_), .A3(new_n213_), .A4(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G231gat), .A2(G233gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT74), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n222_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G57gat), .ZN(new_n226_));
  INV_X1    g025(.A(G64gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G57gat), .A2(G64gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G71gat), .B(G78gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n228_), .A2(new_n234_), .A3(new_n229_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n230_), .A2(new_n232_), .A3(KEYINPUT11), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n225_), .B(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n210_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n241_));
  XNOR2_X1  g040(.A(new_n207_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G232gat), .A2(G233gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n246_), .B(KEYINPUT34), .Z(new_n247_));
  INV_X1    g046(.A(G99gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT10), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G99gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G106gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT64), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G106gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n252_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G85gat), .A2(G92gat), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n259_), .A2(KEYINPUT9), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G99gat), .A2(G106gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT6), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(G85gat), .A2(G92gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(KEYINPUT9), .A3(new_n259_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n258_), .A2(new_n260_), .A3(new_n265_), .A4(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT7), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n270_), .A2(new_n263_), .A3(new_n264_), .A4(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT8), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n266_), .A2(new_n259_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n268_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT67), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n279_), .B(new_n268_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n280_));
  INV_X1    g079(.A(G50gat), .ZN(new_n281_));
  OR2_X1    g080(.A1(G29gat), .A2(G36gat), .ZN(new_n282_));
  INV_X1    g081(.A(G43gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G29gat), .A2(G36gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n283_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n281_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n282_), .A2(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G43gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(G50gat), .A3(new_n285_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(KEYINPUT15), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT15), .ZN(new_n293_));
  NOR3_X1   g092(.A1(new_n286_), .A2(new_n281_), .A3(new_n287_), .ZN(new_n294_));
  AOI21_X1  g093(.A(G50gat), .B1(new_n290_), .B2(new_n285_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n278_), .A2(new_n280_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n288_), .A2(new_n291_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n277_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n247_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n292_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n272_), .A2(new_n274_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT8), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n279_), .B1(new_n305_), .B2(new_n268_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n280_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n301_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n299_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT68), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n247_), .B(KEYINPUT35), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n300_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n308_), .A2(new_n310_), .A3(new_n309_), .A4(new_n312_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT69), .B(G190gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G218gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G134gat), .B(G162gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n320_), .B(KEYINPUT36), .Z(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n320_), .A2(KEYINPUT36), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n314_), .A2(new_n315_), .A3(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT37), .ZN(new_n328_));
  INV_X1    g127(.A(new_n321_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n330_), .B2(KEYINPUT70), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n326_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n327_), .B1(new_n326_), .B2(new_n331_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n330_), .A2(KEYINPUT72), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(KEYINPUT72), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n335_), .A2(new_n328_), .A3(new_n336_), .A4(new_n325_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n245_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(KEYINPUT80), .Z(new_n339_));
  AOI21_X1  g138(.A(new_n238_), .B1(new_n305_), .B2(new_n268_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n238_), .B(new_n268_), .C1(new_n276_), .C2(new_n275_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n305_), .A2(KEYINPUT65), .A3(new_n268_), .A4(new_n238_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n340_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT66), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G230gat), .A2(G233gat), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT12), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n238_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n277_), .A2(new_n237_), .A3(new_n236_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n351_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n341_), .A2(new_n347_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n350_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G120gat), .B(G148gat), .ZN(new_n359_));
  INV_X1    g158(.A(G204gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT5), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G176gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n357_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n363_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT13), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n222_), .A2(new_n298_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n222_), .A2(new_n298_), .ZN(new_n372_));
  OAI211_X1 g171(.A(G229gat), .B(G233gat), .C1(new_n371_), .C2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n301_), .A2(new_n222_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n298_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n221_), .A3(new_n218_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G229gat), .A2(G233gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G113gat), .B(G141gat), .ZN(new_n379_));
  INV_X1    g178(.A(G169gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G197gat), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n373_), .A2(new_n378_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n373_), .B2(new_n378_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n370_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G127gat), .B(G134gat), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n389_), .A2(G113gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(G113gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G120gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(G120gat), .A3(new_n391_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT3), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT2), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  AND2_X1   g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT95), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT1), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n397_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n402_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(new_n406_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n396_), .A2(new_n411_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n401_), .A2(new_n404_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n413_), .A2(new_n394_), .A3(new_n406_), .A4(new_n395_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(KEYINPUT4), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n405_), .A2(new_n410_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n396_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n388_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n388_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n420_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT0), .B(G57gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G85gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(G1gat), .B(G29gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n422_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G176gat), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n432_), .B(KEYINPUT24), .C1(new_n380_), .C2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT25), .ZN(new_n435_));
  INV_X1    g234(.A(G183gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n440_));
  NAND2_X1  g239(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT26), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT26), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n439_), .A2(new_n440_), .A3(new_n442_), .A4(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n437_), .A2(new_n438_), .B1(KEYINPUT26), .B2(new_n441_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n440_), .B1(new_n447_), .B2(new_n444_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n434_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT84), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G183gat), .A2(G190gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(KEYINPUT23), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(KEYINPUT23), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT23), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(G183gat), .A3(G190gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n456_), .A3(KEYINPUT85), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n453_), .B(new_n457_), .C1(new_n432_), .C2(KEYINPUT24), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n460_));
  AND2_X1   g259(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n442_), .B(new_n444_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT82), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n445_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n434_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n450_), .A2(new_n459_), .A3(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n380_), .A2(new_n433_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G169gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(new_n433_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n454_), .A2(new_n456_), .ZN(new_n471_));
  INV_X1    g270(.A(G190gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n436_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  OR2_X1    g274(.A1(G211gat), .A2(G218gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G211gat), .A2(G218gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT90), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(new_n480_), .A3(new_n477_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G197gat), .B(G204gat), .Z(new_n482_));
  AOI22_X1  g281(.A1(new_n479_), .A2(new_n481_), .B1(new_n482_), .B2(KEYINPUT21), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(new_n360_), .B2(G197gat), .ZN(new_n485_));
  INV_X1    g284(.A(G197gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n485_), .A2(new_n487_), .B1(G197gat), .B2(new_n360_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT21), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n479_), .A2(new_n481_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n488_), .A2(new_n489_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n483_), .A2(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n467_), .A2(new_n475_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n431_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n429_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n468_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n497_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT26), .B(G190gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n439_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n498_), .A2(new_n471_), .A3(new_n499_), .A4(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n470_), .A2(KEYINPUT92), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n457_), .A2(new_n473_), .A3(new_n453_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT93), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n470_), .A2(KEYINPUT92), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT93), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n457_), .A2(new_n507_), .A3(new_n473_), .A4(new_n453_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n503_), .A2(new_n505_), .A3(new_n506_), .A4(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n502_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n483_), .A2(new_n490_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n491_), .A2(new_n492_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n494_), .A2(KEYINPUT20), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G226gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT19), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n464_), .A2(new_n465_), .A3(new_n434_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n465_), .B1(new_n464_), .B2(new_n434_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n458_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n475_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n513_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n517_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n502_), .A2(new_n493_), .A3(new_n509_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n523_), .A2(KEYINPUT20), .A3(new_n524_), .A4(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT18), .B(G64gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(G92gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G8gat), .B(G36gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  NAND3_X1  g329(.A1(new_n518_), .A2(new_n526_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n493_), .B1(new_n467_), .B2(new_n475_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n525_), .A2(KEYINPUT20), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n517_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n494_), .A2(KEYINPUT20), .A3(new_n524_), .A4(new_n514_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n530_), .B(KEYINPUT97), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n531_), .B(KEYINPUT27), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n518_), .A2(new_n530_), .A3(new_n526_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n530_), .B1(new_n518_), .B2(new_n526_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n428_), .B(new_n538_), .C1(new_n541_), .C2(KEYINPUT27), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT29), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n413_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT28), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G228gat), .A2(G233gat), .ZN(new_n547_));
  INV_X1    g346(.A(G22gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n546_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n513_), .B1(new_n544_), .B2(new_n413_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(new_n281_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G78gat), .B(G106gat), .Z(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n553_), .A2(new_n554_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n551_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n555_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n550_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n396_), .B(KEYINPUT31), .Z(new_n561_));
  XNOR2_X1  g360(.A(G15gat), .B(G43gat), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n467_), .A2(new_n563_), .A3(new_n475_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n467_), .B2(new_n475_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n562_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G71gat), .B(G99gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G227gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT86), .B(KEYINPUT87), .Z(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT30), .B1(new_n521_), .B2(new_n522_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n562_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n467_), .A2(new_n563_), .A3(new_n475_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n566_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n571_), .B1(new_n566_), .B2(new_n575_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT88), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n571_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n564_), .A2(new_n565_), .A3(new_n562_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n573_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n580_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n566_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT88), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n561_), .B1(new_n579_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n584_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n561_), .B1(new_n587_), .B2(new_n578_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n560_), .B1(new_n586_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n561_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n578_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n583_), .A2(KEYINPUT88), .A3(new_n584_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n557_), .A2(new_n559_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n594_), .A2(new_n588_), .A3(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n543_), .B1(new_n590_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n592_), .A2(new_n593_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n588_), .B1(new_n598_), .B2(new_n561_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT94), .B1(new_n539_), .B2(new_n540_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n518_), .A2(new_n526_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n530_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n531_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n426_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(KEYINPUT33), .B(new_n426_), .C1(new_n419_), .C2(new_n421_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n415_), .A2(new_n388_), .A3(new_n418_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n426_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n412_), .A2(new_n420_), .A3(new_n414_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n608_), .A2(new_n609_), .A3(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n600_), .A2(new_n605_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT96), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n518_), .A2(new_n526_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n536_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n530_), .A2(KEYINPUT32), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n518_), .A2(new_n526_), .A3(KEYINPUT96), .A4(new_n619_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n427_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n615_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n599_), .A2(new_n624_), .A3(new_n595_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n597_), .A2(new_n625_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n339_), .A2(new_n387_), .A3(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n214_), .A3(new_n427_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT99), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n335_), .A2(new_n336_), .A3(new_n325_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n626_), .A2(new_n632_), .A3(new_n244_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n387_), .B(KEYINPUT98), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G1gat), .B1(new_n636_), .B2(new_n428_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n631_), .B(new_n637_), .C1(new_n629_), .C2(new_n628_), .ZN(G1324gat));
  OAI21_X1  g437(.A(new_n538_), .B1(new_n541_), .B2(KEYINPUT27), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT100), .B1(new_n636_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n634_), .A2(new_n642_), .A3(new_n635_), .A4(new_n639_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n641_), .A2(G8gat), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT39), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n641_), .A2(new_n646_), .A3(G8gat), .A4(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n627_), .A2(new_n215_), .A3(new_n639_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(KEYINPUT40), .A3(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n636_), .B2(new_n599_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT41), .Z(new_n656_));
  INV_X1    g455(.A(G15gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n599_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n627_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT101), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n656_), .A2(new_n660_), .ZN(G1326gat));
  OAI21_X1  g460(.A(G22gat), .B1(new_n636_), .B2(new_n595_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT42), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n627_), .A2(new_n548_), .A3(new_n560_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1327gat));
  NAND2_X1  g464(.A1(new_n326_), .A2(new_n331_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT71), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n326_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n337_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n586_), .A2(new_n589_), .A3(new_n560_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n595_), .B1(new_n594_), .B2(new_n588_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n542_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n599_), .A2(new_n624_), .A3(new_n595_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n675_), .A2(KEYINPUT102), .A3(KEYINPUT43), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT43), .B1(new_n675_), .B2(KEYINPUT102), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n245_), .B(new_n635_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n669_), .B1(new_n597_), .B2(new_n625_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n675_), .A2(KEYINPUT102), .A3(KEYINPUT43), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n686_), .A2(KEYINPUT44), .A3(new_n245_), .A4(new_n635_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n680_), .A2(new_n427_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n632_), .B1(new_n597_), .B2(new_n625_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n690_), .A2(new_n387_), .A3(new_n245_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n428_), .A2(G29gat), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT103), .Z(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(new_n694_), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n680_), .A2(new_n639_), .A3(new_n687_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698_));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n691_), .A2(new_n698_), .A3(new_n699_), .A4(new_n639_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n690_), .A2(new_n699_), .A3(new_n387_), .A4(new_n245_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT104), .B1(new_n701_), .B2(new_n640_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n700_), .A2(KEYINPUT45), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT45), .B1(new_n700_), .B2(new_n702_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n697_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT46), .B1(new_n706_), .B2(KEYINPUT105), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n708_), .B(new_n709_), .C1(new_n697_), .C2(new_n705_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1329gat));
  XNOR2_X1  g510(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n599_), .A2(new_n283_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n680_), .A2(new_n687_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n680_), .A2(KEYINPUT106), .A3(new_n687_), .A4(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G43gat), .B1(new_n691_), .B2(new_n658_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n712_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n712_), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n722_), .B(new_n719_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1330gat));
  AND4_X1   g523(.A1(G50gat), .A2(new_n680_), .A3(new_n560_), .A4(new_n687_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G50gat), .B1(new_n691_), .B2(new_n560_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1331gat));
  NOR2_X1   g526(.A1(new_n370_), .A2(new_n386_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n634_), .A2(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n729_), .A2(new_n226_), .A3(new_n428_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n339_), .A2(new_n626_), .A3(new_n728_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n427_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n730_), .B1(new_n226_), .B2(new_n733_), .ZN(G1332gat));
  OAI21_X1  g533(.A(G64gat), .B1(new_n729_), .B2(new_n640_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT48), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(new_n227_), .A3(new_n639_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1333gat));
  OAI21_X1  g537(.A(G71gat), .B1(new_n729_), .B2(new_n599_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT108), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT49), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n741_), .ZN(new_n743_));
  OR3_X1    g542(.A1(new_n731_), .A2(G71gat), .A3(new_n599_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n729_), .B2(new_n595_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT50), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n595_), .A2(G78gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n731_), .B2(new_n748_), .ZN(G1335gat));
  AND3_X1   g548(.A1(new_n690_), .A2(new_n245_), .A3(new_n728_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n427_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n244_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n728_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(new_n428_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n751_), .B1(new_n754_), .B2(G85gat), .ZN(G1336gat));
  INV_X1    g554(.A(G92gat), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n753_), .A2(new_n756_), .A3(new_n640_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G92gat), .B1(new_n750_), .B2(new_n639_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1337gat));
  NAND3_X1  g558(.A1(new_n750_), .A2(new_n252_), .A3(new_n658_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT110), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n752_), .A2(new_n658_), .A3(new_n728_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n762_), .A2(KEYINPUT109), .A3(G99gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT109), .B1(new_n762_), .B2(G99gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  AND2_X1   g564(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(G1338gat));
  XNOR2_X1  g566(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n768_));
  OAI21_X1  g567(.A(G106gat), .B1(new_n753_), .B2(new_n595_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT52), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(G106gat), .C1(new_n753_), .C2(new_n595_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n750_), .A2(new_n257_), .A3(new_n560_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n768_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n768_), .ZN(new_n777_));
  AOI211_X1 g576(.A(new_n777_), .B(new_n774_), .C1(new_n770_), .C2(new_n772_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1339gat));
  XNOR2_X1  g578(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n338_), .A2(new_n385_), .A3(new_n370_), .A4(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n370_), .A2(new_n669_), .A3(new_n385_), .A4(new_n244_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n780_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n385_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n343_), .A2(new_n344_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n353_), .A2(new_n787_), .A3(new_n355_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n347_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n357_), .A2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n353_), .A2(KEYINPUT55), .A3(new_n355_), .A4(new_n356_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n363_), .ZN(new_n795_));
  XOR2_X1   g594(.A(KEYINPUT114), .B(KEYINPUT56), .Z(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(new_n794_), .B2(new_n363_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n786_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n377_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n374_), .A2(new_n376_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n377_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n382_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(new_n383_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n369_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n786_), .B(KEYINPUT115), .C1(new_n795_), .C2(new_n797_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n800_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT57), .B1(new_n808_), .B2(new_n632_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(KEYINPUT57), .A3(new_n632_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n363_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n368_), .B(new_n805_), .C1(new_n795_), .C2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n794_), .A2(new_n363_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n363_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(KEYINPUT58), .A3(new_n368_), .A4(new_n805_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n815_), .A2(new_n821_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n822_), .A2(new_n669_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n810_), .A2(new_n811_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n785_), .B1(new_n245_), .B2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n639_), .A2(new_n428_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n590_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828_), .B2(new_n386_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n808_), .A2(KEYINPUT57), .A3(new_n632_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n822_), .A2(new_n669_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n831_), .A2(new_n809_), .A3(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n830_), .B1(new_n833_), .B2(new_n244_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n785_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n824_), .A2(KEYINPUT116), .A3(new_n245_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n827_), .A2(KEYINPUT59), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT59), .B1(new_n825_), .B2(new_n827_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n386_), .A2(G113gat), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT118), .Z(new_n846_));
  AOI21_X1  g645(.A(new_n829_), .B1(new_n844_), .B2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(new_n370_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n839_), .A2(new_n848_), .A3(new_n841_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G120gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n393_), .B1(new_n370_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n828_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n393_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1341gat));
  AOI21_X1  g652(.A(G127gat), .B1(new_n828_), .B2(new_n244_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n244_), .A2(G127gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n844_), .B2(new_n855_), .ZN(G1342gat));
  XOR2_X1   g655(.A(KEYINPUT119), .B(G134gat), .Z(new_n857_));
  NOR2_X1   g656(.A1(new_n669_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n842_), .A2(new_n843_), .A3(new_n859_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n825_), .A2(new_n632_), .A3(new_n827_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(G134gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT120), .B1(new_n860_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n843_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n858_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867_));
  INV_X1    g666(.A(new_n862_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n863_), .A2(new_n869_), .ZN(G1343gat));
  NOR2_X1   g669(.A1(new_n825_), .A2(new_n671_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n826_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n386_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n848_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g676(.A1(new_n872_), .A2(new_n245_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT121), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n878_), .B(new_n880_), .ZN(G1346gat));
  NOR2_X1   g680(.A1(new_n872_), .A2(new_n632_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n670_), .A2(G162gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT122), .ZN(new_n884_));
  OAI22_X1  g683(.A1(new_n882_), .A2(G162gat), .B1(new_n872_), .B2(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT123), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n640_), .A2(new_n427_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n590_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n837_), .A2(new_n386_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G169gat), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n891_), .A2(KEYINPUT124), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(KEYINPUT124), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(KEYINPUT62), .A3(new_n893_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n837_), .A2(new_n889_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n386_), .A3(new_n469_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n891_), .A2(KEYINPUT124), .A3(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n894_), .A2(new_n896_), .A3(new_n898_), .ZN(G1348gat));
  NOR2_X1   g698(.A1(new_n825_), .A2(new_n888_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(G176gat), .A3(new_n848_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n895_), .A2(new_n848_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n903_), .B(KEYINPUT126), .C1(G176gat), .C2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n901_), .B(KEYINPUT125), .ZN(new_n907_));
  AOI21_X1  g706(.A(G176gat), .B1(new_n895_), .B2(new_n848_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n909_), .ZN(G1349gat));
  AOI21_X1  g709(.A(G183gat), .B1(new_n900_), .B2(new_n244_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n245_), .A2(new_n439_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n895_), .B2(new_n912_), .ZN(G1350gat));
  INV_X1    g712(.A(new_n632_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n895_), .A2(new_n500_), .A3(new_n914_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n895_), .A2(new_n670_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n472_), .ZN(G1351gat));
  NAND2_X1  g716(.A1(new_n871_), .A2(new_n887_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n385_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(new_n486_), .ZN(G1352gat));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n370_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n360_), .ZN(G1353gat));
  INV_X1    g721(.A(new_n918_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n244_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  AND2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n927_), .B1(new_n924_), .B2(new_n925_), .ZN(G1354gat));
  NOR2_X1   g727(.A1(new_n918_), .A2(new_n632_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n670_), .A2(G218gat), .ZN(new_n930_));
  OAI22_X1  g729(.A1(new_n929_), .A2(G218gat), .B1(new_n918_), .B2(new_n930_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


