//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT80), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G141gat), .ZN(new_n208_));
  INV_X1    g007(.A(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT81), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n216_), .B(new_n217_), .C1(new_n218_), .C2(new_n211_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n203_), .B(new_n204_), .C1(new_n214_), .C2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n212_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT82), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G127gat), .B(G134gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n224_), .B(new_n225_), .Z(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n221_), .A2(new_n226_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G225gat), .A2(G233gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G1gat), .B(G29gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G85gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT0), .B(G57gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n232_), .B(new_n233_), .Z(new_n234_));
  AND3_X1   g033(.A1(new_n227_), .A2(KEYINPUT4), .A3(new_n228_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n223_), .A2(new_n236_), .A3(new_n226_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n229_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n230_), .B(new_n234_), .C1(new_n235_), .C2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT93), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT33), .ZN(new_n243_));
  XOR2_X1   g042(.A(G8gat), .B(G36gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(G64gat), .B(G92gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT20), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G183gat), .A2(G190gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT23), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(G183gat), .B2(G190gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT89), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n254_), .A2(KEYINPUT89), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n253_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT22), .B(G169gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT90), .ZN(new_n259_));
  INV_X1    g058(.A(G176gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n262_), .A2(KEYINPUT24), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n252_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G190gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT25), .B(G183gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n262_), .A2(KEYINPUT24), .A3(new_n254_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n257_), .A2(new_n261_), .B1(new_n265_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G197gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT84), .B1(new_n272_), .B2(G204gat), .ZN(new_n273_));
  INV_X1    g072(.A(G204gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n273_), .B1(G197gat), .B2(new_n274_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n272_), .A2(KEYINPUT84), .A3(G204gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT21), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G211gat), .B(G218gat), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n272_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT85), .B1(new_n272_), .B2(G204gat), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n279_), .B(new_n280_), .C1(G197gat), .C2(new_n274_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n277_), .B(new_n278_), .C1(KEYINPUT21), .C2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT21), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n250_), .B1(new_n271_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT88), .ZN(new_n289_));
  XOR2_X1   g088(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G183gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT25), .B1(new_n293_), .B2(KEYINPUT74), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n293_), .A2(KEYINPUT25), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n266_), .B(new_n294_), .C1(new_n295_), .C2(KEYINPUT74), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n269_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n264_), .B1(new_n297_), .B2(KEYINPUT75), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(KEYINPUT75), .B2(new_n297_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n258_), .A2(new_n260_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n300_), .B(KEYINPUT76), .Z(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n254_), .A3(new_n253_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n287_), .B(new_n292_), .C1(new_n303_), .C2(new_n286_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n286_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n257_), .A2(new_n261_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n265_), .A2(new_n270_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n282_), .A2(new_n285_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n250_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n292_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n249_), .B1(new_n305_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT92), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n299_), .A2(new_n302_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(new_n310_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT20), .B1(new_n271_), .B2(new_n286_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n291_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(new_n304_), .A3(new_n248_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n313_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n305_), .A2(new_n312_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(KEYINPUT92), .A3(new_n248_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n234_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n227_), .A2(new_n228_), .A3(new_n238_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n237_), .A2(new_n229_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n324_), .B(new_n325_), .C1(new_n235_), .C2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT33), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n240_), .A2(new_n241_), .A3(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n243_), .A2(new_n323_), .A3(new_n327_), .A4(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n230_), .B1(new_n235_), .B2(new_n239_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n324_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(KEYINPUT94), .A3(new_n240_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT94), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n334_), .A3(new_n324_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n248_), .A2(KEYINPUT32), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n287_), .B1(new_n303_), .B2(new_n286_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n291_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n306_), .A2(new_n292_), .A3(new_n311_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n321_), .B2(new_n336_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n333_), .A2(new_n335_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n330_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G71gat), .B(G99gat), .ZN(new_n344_));
  INV_X1    g143(.A(G43gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT30), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(new_n226_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT77), .B(G15gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n303_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT79), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n315_), .A2(new_n352_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n349_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(new_n348_), .A3(new_n359_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT83), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n367_), .A2(G228gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(G228gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n366_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n286_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n221_), .B(KEYINPUT82), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n212_), .B2(new_n220_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n370_), .B1(new_n286_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G78gat), .B(G106gat), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n223_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT28), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n381_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT28), .B1(new_n223_), .B2(KEYINPUT29), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n372_), .A2(new_n383_), .A3(new_n373_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n381_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n379_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n374_), .A2(new_n377_), .A3(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n380_), .A2(new_n385_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n380_), .A2(new_n391_), .B1(new_n385_), .B2(new_n389_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n365_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n343_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n380_), .A2(new_n391_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n389_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n388_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n365_), .A2(new_n392_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n362_), .A2(new_n364_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n402_), .A2(new_n404_), .B1(new_n335_), .B2(new_n333_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n320_), .A2(new_n322_), .A3(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n338_), .A2(new_n339_), .ZN(new_n408_));
  OAI211_X1 g207(.A(KEYINPUT27), .B(new_n319_), .C1(new_n408_), .C2(new_n248_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n405_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n397_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G232gat), .A2(G233gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G29gat), .B(G36gat), .Z(new_n416_));
  XOR2_X1   g215(.A(G43gat), .B(G50gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT7), .ZN(new_n421_));
  INV_X1    g220(.A(G99gat), .ZN(new_n422_));
  INV_X1    g221(.A(G106gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G99gat), .A2(G106gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT6), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(G99gat), .A3(G106gat), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n429_), .A2(new_n431_), .A3(KEYINPUT67), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT67), .B1(new_n429_), .B2(new_n431_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n427_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(G85gat), .A2(G92gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G85gat), .A2(G92gat), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n437_), .A2(KEYINPUT8), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n435_), .A2(new_n436_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n429_), .A2(new_n431_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n439_), .B1(new_n440_), .B2(new_n426_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n434_), .A2(new_n438_), .B1(new_n441_), .B2(KEYINPUT8), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n422_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n423_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT64), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n444_), .A2(KEYINPUT64), .A3(new_n423_), .A4(new_n445_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n448_), .B(new_n449_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n450_));
  OR2_X1    g249(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G92gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n455_));
  INV_X1    g254(.A(G92gat), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n456_), .A2(KEYINPUT9), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n454_), .A2(new_n455_), .B1(new_n437_), .B2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n450_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n442_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n420_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n429_), .A2(new_n431_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT67), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n429_), .A2(new_n431_), .A3(KEYINPUT67), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n426_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n438_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n437_), .B1(new_n427_), .B2(new_n462_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT8), .ZN(new_n469_));
  OAI22_X1  g268(.A1(new_n466_), .A2(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n437_), .A2(new_n457_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n456_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n455_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n464_), .A2(new_n465_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n449_), .A4(new_n448_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n477_), .A2(new_n418_), .ZN(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT72), .B(new_n415_), .C1(new_n461_), .C2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G190gat), .B(G218gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G134gat), .B(G162gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT36), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n461_), .A2(new_n478_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n479_), .B(new_n483_), .C1(new_n484_), .C2(KEYINPUT35), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n415_), .B1(new_n484_), .B2(KEYINPUT72), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n482_), .A2(KEYINPUT36), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT98), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT98), .ZN(new_n492_));
  INV_X1    g291(.A(new_n490_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n488_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n412_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT73), .B(G1gat), .ZN(new_n498_));
  INV_X1    g297(.A(G8gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT14), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n497_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G1gat), .B(G8gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n497_), .B(new_n503_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n420_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n507_), .B2(new_n418_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n418_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n418_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n509_), .A2(new_n512_), .B1(new_n516_), .B2(new_n511_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G113gat), .B(G141gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(G169gat), .B(G197gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n517_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G71gat), .B(G78gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(KEYINPUT11), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n526_));
  INV_X1    g325(.A(new_n524_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n525_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n507_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G127gat), .B(G155gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT16), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G183gat), .B(G211gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n537_), .A2(new_n538_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n533_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n533_), .A2(new_n539_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G230gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n460_), .B2(new_n530_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n530_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n442_), .B2(new_n459_), .ZN(new_n549_));
  XOR2_X1   g348(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(KEYINPUT12), .B(new_n525_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n442_), .B2(new_n459_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT68), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n477_), .A2(new_n556_), .A3(new_n553_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n547_), .A2(new_n551_), .A3(new_n555_), .A4(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n470_), .A2(new_n476_), .A3(new_n530_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n549_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n546_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G120gat), .B(G148gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT5), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n558_), .A2(new_n561_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n565_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n568_), .B1(new_n571_), .B2(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR4_X1   g373(.A1(new_n496_), .A2(new_n522_), .A3(new_n544_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n333_), .A2(new_n335_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(G1gat), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n343_), .A2(new_n396_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(new_n522_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n489_), .A2(KEYINPUT37), .A3(new_n490_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n493_), .B2(new_n488_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(new_n544_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n581_), .A2(new_n586_), .A3(new_n573_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT96), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(KEYINPUT96), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n591_), .A2(new_n498_), .A3(new_n577_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n591_), .A2(KEYINPUT38), .A3(new_n498_), .A4(new_n577_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT97), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT97), .ZN(new_n595_));
  OAI221_X1 g394(.A(new_n579_), .B1(KEYINPUT38), .B2(new_n592_), .C1(new_n594_), .C2(new_n595_), .ZN(G1324gat));
  XNOR2_X1  g395(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n597_));
  INV_X1    g396(.A(new_n410_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n575_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT99), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(G8gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n599_), .B2(G8gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT39), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n603_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n601_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n598_), .A2(new_n499_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n590_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n597_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n597_), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n610_), .B(new_n613_), .C1(new_n604_), .C2(new_n607_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n612_), .A2(new_n614_), .ZN(G1325gat));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n575_), .B2(new_n403_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT41), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n591_), .A2(new_n616_), .A3(new_n403_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1326gat));
  INV_X1    g419(.A(G22gat), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n393_), .A2(new_n394_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT101), .Z(new_n623_));
  AOI21_X1  g422(.A(new_n621_), .B1(new_n575_), .B2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT42), .Z(new_n625_));
  NAND3_X1  g424(.A1(new_n591_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1327gat));
  NAND2_X1  g426(.A1(new_n491_), .A2(new_n494_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n544_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(new_n574_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n581_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT104), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n581_), .A2(new_n633_), .A3(new_n630_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(G29gat), .B1(new_n635_), .B2(new_n577_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n402_), .A2(new_n404_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n638_), .A2(new_n410_), .A3(new_n576_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n395_), .B1(new_n330_), .B2(new_n342_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n637_), .B(new_n585_), .C1(new_n639_), .C2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n412_), .A2(KEYINPUT102), .A3(new_n637_), .A4(new_n585_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n585_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT43), .B1(new_n580_), .B2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n574_), .A2(new_n522_), .A3(new_n543_), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT44), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(KEYINPUT44), .A3(new_n648_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT103), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n647_), .A2(new_n652_), .A3(KEYINPUT44), .A4(new_n648_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n649_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n577_), .A2(G29gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n636_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  INV_X1    g455(.A(G36gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n635_), .A2(new_n657_), .A3(new_n598_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n658_), .B(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n654_), .A2(new_n598_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n661_), .B(KEYINPUT46), .C1(new_n662_), .C2(new_n657_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT46), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n658_), .B(new_n659_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n657_), .B1(new_n654_), .B2(new_n598_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(G1329gat));
  NAND2_X1  g467(.A1(new_n651_), .A2(new_n653_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670_));
  INV_X1    g469(.A(new_n649_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n365_), .A2(new_n345_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .A4(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT47), .ZN(new_n674_));
  INV_X1    g473(.A(new_n672_), .ZN(new_n675_));
  AOI211_X1 g474(.A(new_n649_), .B(new_n675_), .C1(new_n651_), .C2(new_n653_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n632_), .A2(new_n403_), .A3(new_n634_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n670_), .B1(new_n677_), .B2(new_n345_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n673_), .B(new_n674_), .C1(new_n676_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n669_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n678_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n674_), .B1(new_n683_), .B2(new_n673_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1330gat));
  AOI21_X1  g484(.A(G50gat), .B1(new_n635_), .B2(new_n623_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n622_), .A2(G50gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n654_), .B2(new_n687_), .ZN(G1331gat));
  NOR2_X1   g487(.A1(new_n580_), .A2(new_n521_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n585_), .A2(new_n573_), .A3(new_n544_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n691_), .A2(G57gat), .A3(new_n576_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n574_), .A2(new_n522_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n496_), .A2(new_n544_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n577_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n692_), .B1(G57gat), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT107), .ZN(G1332gat));
  INV_X1    g496(.A(G64gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n694_), .B2(new_n598_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT48), .Z(new_n700_));
  INV_X1    g499(.A(new_n691_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n698_), .A3(new_n598_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1333gat));
  INV_X1    g502(.A(G71gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n694_), .B2(new_n403_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT49), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n701_), .A2(new_n704_), .A3(new_n403_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1334gat));
  INV_X1    g507(.A(G78gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n694_), .B2(new_n623_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT50), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n701_), .A2(new_n709_), .A3(new_n623_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1335gat));
  NOR4_X1   g512(.A1(new_n580_), .A2(new_n521_), .A3(new_n573_), .A4(new_n629_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n577_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n693_), .A2(new_n543_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n647_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n576_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n715_), .B1(new_n717_), .B2(new_n718_), .ZN(G1336gat));
  NAND3_X1  g518(.A1(new_n714_), .A2(new_n456_), .A3(new_n598_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n717_), .A2(new_n598_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n456_), .ZN(G1337gat));
  NAND2_X1  g521(.A1(new_n717_), .A2(new_n403_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G99gat), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n714_), .A2(new_n403_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n727_), .A2(KEYINPUT109), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(KEYINPUT109), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n724_), .A2(new_n725_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT51), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n729_), .A3(new_n731_), .ZN(G1338gat));
  NAND3_X1  g531(.A1(new_n714_), .A2(new_n423_), .A3(new_n622_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n717_), .A2(new_n622_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(G106gat), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT52), .B(new_n423_), .C1(new_n717_), .C2(new_n622_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g538(.A1(new_n558_), .A2(KEYINPUT55), .ZN(new_n740_));
  AOI22_X1  g539(.A1(KEYINPUT68), .A2(new_n554_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n557_), .A4(new_n547_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n551_), .A2(new_n555_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n546_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n565_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(KEYINPUT110), .A3(new_n749_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n740_), .A2(new_n743_), .B1(new_n546_), .B2(new_n745_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n751_), .B2(new_n565_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753_));
  INV_X1    g552(.A(new_n749_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n751_), .B2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n750_), .A2(new_n752_), .A3(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n522_), .A2(new_n566_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n520_), .B1(new_n516_), .B2(new_n510_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n509_), .A2(new_n513_), .A3(new_n511_), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n517_), .A2(new_n520_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT111), .B(new_n761_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n758_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n495_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT57), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n766_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT112), .B1(new_n772_), .B2(new_n628_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n771_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n747_), .A2(new_n775_), .A3(new_n749_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT113), .B1(new_n751_), .B2(new_n754_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n752_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n566_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(new_n761_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT114), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT58), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(KEYINPUT114), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n585_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n774_), .A2(new_n786_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n787_), .A2(KEYINPUT117), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n772_), .A2(new_n628_), .A3(new_n771_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n787_), .B2(KEYINPUT117), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n543_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n586_), .A2(new_n522_), .A3(new_n573_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n792_), .A2(KEYINPUT54), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(KEYINPUT54), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n791_), .A2(new_n796_), .ZN(new_n797_));
  OR3_X1    g596(.A1(new_n598_), .A2(new_n576_), .A3(new_n404_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT116), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n800_));
  INV_X1    g599(.A(new_n789_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n774_), .A2(new_n786_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n774_), .A2(new_n786_), .A3(KEYINPUT115), .A4(new_n801_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n544_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n795_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n799_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n797_), .A2(new_n800_), .B1(new_n809_), .B2(KEYINPUT59), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n521_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G113gat), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n522_), .A2(G113gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n809_), .B2(new_n813_), .ZN(G1340gat));
  AND2_X1   g613(.A1(new_n810_), .A2(new_n574_), .ZN(new_n815_));
  XOR2_X1   g614(.A(KEYINPUT118), .B(G120gat), .Z(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(KEYINPUT60), .B2(new_n816_), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n815_), .A2(new_n816_), .B1(new_n809_), .B2(new_n818_), .ZN(G1341gat));
  NAND2_X1  g618(.A1(new_n810_), .A2(new_n543_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(G127gat), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n544_), .A2(G127gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n809_), .B2(new_n822_), .ZN(G1342gat));
  OAI21_X1  g622(.A(new_n800_), .B1(new_n791_), .B2(new_n796_), .ZN(new_n824_));
  INV_X1    g623(.A(G134gat), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n645_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n799_), .B1(new_n806_), .B2(new_n795_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n824_), .B(new_n826_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n830_), .B(G134gat), .C1(new_n828_), .C2(new_n628_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n807_), .A2(new_n628_), .A3(new_n808_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT119), .B1(new_n832_), .B2(new_n825_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n829_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n829_), .B(KEYINPUT120), .C1(new_n831_), .C2(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1343gat));
  INV_X1    g637(.A(new_n402_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n807_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n598_), .A2(new_n576_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n521_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n574_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT121), .B(G148gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1345gat));
  NAND2_X1  g647(.A1(new_n843_), .A2(new_n543_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT61), .B(G155gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1346gat));
  AOI21_X1  g650(.A(new_n402_), .B1(new_n806_), .B2(new_n795_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n585_), .A2(G162gat), .ZN(new_n853_));
  XOR2_X1   g652(.A(new_n853_), .B(KEYINPUT122), .Z(new_n854_));
  AND3_X1   g653(.A1(new_n852_), .A2(new_n841_), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n840_), .A2(new_n495_), .A3(new_n842_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(G162gat), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n856_), .B(KEYINPUT123), .C1(G162gat), .C2(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1347gat));
  NOR2_X1   g661(.A1(new_n410_), .A2(new_n577_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n403_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n623_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n521_), .B(new_n865_), .C1(new_n791_), .C2(new_n796_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G169gat), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(KEYINPUT62), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n797_), .A2(new_n865_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n521_), .A3(new_n259_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n871_), .B(new_n874_), .C1(KEYINPUT62), .C2(new_n869_), .ZN(G1348gat));
  AOI21_X1  g674(.A(G176gat), .B1(new_n873_), .B2(new_n574_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n622_), .B1(new_n806_), .B2(new_n795_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n864_), .A2(new_n260_), .A3(new_n573_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(G1349gat));
  NOR2_X1   g678(.A1(new_n544_), .A2(new_n267_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT125), .B1(new_n873_), .B2(new_n880_), .ZN(new_n881_));
  AND4_X1   g680(.A1(KEYINPUT125), .A2(new_n797_), .A3(new_n865_), .A4(new_n880_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n864_), .A2(new_n544_), .ZN(new_n883_));
  AOI21_X1  g682(.A(G183gat), .B1(new_n877_), .B2(new_n883_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n881_), .A2(new_n882_), .A3(new_n884_), .ZN(G1350gat));
  OAI21_X1  g684(.A(G190gat), .B1(new_n872_), .B2(new_n645_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n628_), .A2(new_n266_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n872_), .B2(new_n887_), .ZN(G1351gat));
  NAND2_X1  g687(.A1(new_n852_), .A2(new_n863_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT126), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n852_), .A2(new_n891_), .A3(new_n863_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G197gat), .B1(new_n893_), .B2(new_n521_), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n272_), .B(new_n522_), .C1(new_n890_), .C2(new_n892_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1352gat));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n574_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G204gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n893_), .A2(new_n274_), .A3(new_n574_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1353gat));
  XOR2_X1   g699(.A(KEYINPUT63), .B(G211gat), .Z(new_n901_));
  INV_X1    g700(.A(new_n892_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n891_), .B1(new_n852_), .B2(new_n863_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n543_), .B(new_n901_), .C1(new_n902_), .C2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n544_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n905_));
  OR2_X1    g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(G1354gat));
  NAND2_X1  g707(.A1(new_n893_), .A2(new_n628_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT127), .B(G218gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n645_), .A2(new_n910_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n909_), .A2(new_n910_), .B1(new_n893_), .B2(new_n911_), .ZN(G1355gat));
endmodule


