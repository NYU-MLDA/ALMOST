//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n973_, new_n974_, new_n976_, new_n977_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n984_, new_n985_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n992_, new_n993_;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G92gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G85gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT9), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n206_), .A2(new_n210_), .A3(new_n215_), .A4(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n207_), .A2(new_n208_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AOI211_X1 g024(.A(KEYINPUT8), .B(new_n221_), .C1(new_n225_), .C2(new_n215_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n217_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n213_), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n222_), .B(new_n230_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n227_), .B1(new_n233_), .B2(new_n209_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n220_), .B1(new_n226_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G71gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G78gat), .ZN(new_n237_));
  INV_X1    g036(.A(G78gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G71gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(KEYINPUT11), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n243_), .B1(new_n241_), .B2(KEYINPUT11), .ZN(new_n244_));
  INV_X1    g043(.A(G64gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G57gat), .ZN(new_n246_));
  INV_X1    g045(.A(G57gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G64gat), .ZN(new_n248_));
  AND4_X1   g047(.A1(new_n243_), .A2(new_n246_), .A3(new_n248_), .A4(KEYINPUT11), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n242_), .B1(new_n244_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT11), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT65), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(new_n248_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n246_), .A2(new_n248_), .A3(new_n243_), .A4(KEYINPUT11), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n252_), .A2(new_n255_), .A3(new_n240_), .A4(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n250_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n202_), .B1(new_n235_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n219_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n215_), .B1(new_n221_), .B2(new_n204_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n231_), .A2(new_n232_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n230_), .A2(new_n222_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n209_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT8), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n233_), .A2(new_n227_), .A3(new_n209_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n262_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n250_), .A2(new_n257_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(KEYINPUT66), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n235_), .A2(new_n258_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n259_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G230gat), .A2(G233gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n274_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n268_), .A2(KEYINPUT12), .A3(new_n269_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(new_n235_), .B2(new_n258_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n276_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G120gat), .B(G148gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT5), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G176gat), .B(G204gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n285_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n275_), .A2(new_n280_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT13), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n290_), .A2(KEYINPUT67), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(KEYINPUT67), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(KEYINPUT13), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n293_), .A2(KEYINPUT68), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(KEYINPUT68), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n291_), .A2(new_n292_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT69), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G226gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G211gat), .B(G218gat), .Z(new_n302_));
  INV_X1    g101(.A(KEYINPUT21), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G197gat), .B(G204gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(KEYINPUT86), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT86), .ZN(new_n307_));
  INV_X1    g106(.A(G197gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(G204gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(KEYINPUT21), .A3(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n304_), .A2(new_n303_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n305_), .A2(new_n310_), .B1(new_n302_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT22), .B(G169gat), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT92), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(KEYINPUT92), .A3(new_n316_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(G183gat), .A3(G190gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G183gat), .ZN(new_n324_));
  INV_X1    g123(.A(G190gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT23), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(KEYINPUT79), .B(KEYINPUT23), .C1(new_n324_), .C2(new_n325_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n323_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n319_), .B(new_n320_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT26), .B(G190gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT25), .B(G183gat), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n336_), .A2(new_n337_), .B1(new_n326_), .B2(new_n322_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n316_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT91), .B1(new_n333_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n334_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n333_), .A2(KEYINPUT91), .A3(new_n339_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n335_), .B(new_n338_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n312_), .B1(new_n332_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n326_), .A2(new_n322_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT78), .B(G183gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(G190gat), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(G169gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(KEYINPUT80), .A2(KEYINPUT22), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(new_n314_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n351_), .B1(new_n334_), .B2(new_n350_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G183gat), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n336_), .B(new_n355_), .C1(new_n347_), .C2(new_n354_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n341_), .A2(KEYINPUT24), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n341_), .A2(KEYINPUT24), .A3(new_n316_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n353_), .B1(new_n359_), .B2(new_n330_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n305_), .A2(new_n310_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n311_), .A2(new_n302_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT20), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n301_), .B1(new_n345_), .B2(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G8gat), .B(G36gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT18), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n332_), .A2(new_n312_), .A3(new_n344_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n300_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n365_), .A2(new_n369_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n364_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n332_), .A2(new_n344_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n363_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n300_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n371_), .A2(new_n372_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n301_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n369_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n375_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n365_), .A2(new_n373_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n369_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT27), .B1(new_n387_), .B2(new_n374_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G228gat), .ZN(new_n390_));
  INV_X1    g189(.A(G233gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT85), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(G233gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(new_n238_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n396_), .A2(G106gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(G106gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(G141gat), .A2(G148gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT3), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G141gat), .A2(G148gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT2), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(KEYINPUT1), .B2(new_n405_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(KEYINPUT1), .B2(new_n405_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n400_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n412_), .A2(new_n402_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n312_), .B1(new_n415_), .B2(KEYINPUT29), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n399_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n404_), .A2(new_n408_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT29), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI22_X1  g220(.A1(new_n421_), .A2(new_n312_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n418_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n417_), .A2(KEYINPUT87), .A3(new_n422_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G22gat), .B(G50gat), .Z(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT28), .B1(new_n415_), .B2(KEYINPUT29), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n419_), .A2(new_n430_), .A3(new_n420_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n428_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n429_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n427_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n428_), .A2(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT83), .ZN(new_n437_));
  INV_X1    g236(.A(new_n427_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n432_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n425_), .A2(new_n426_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n425_), .A2(new_n435_), .A3(new_n439_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT88), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n425_), .A2(new_n426_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n435_), .A2(new_n439_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n425_), .A2(new_n435_), .A3(new_n439_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n443_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n389_), .B1(new_n442_), .B2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G71gat), .B(G99gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n330_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n452_), .A2(new_n356_), .A3(new_n357_), .A4(new_n358_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(KEYINPUT30), .A3(new_n353_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT30), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n360_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G15gat), .B(G43gat), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G227gat), .A2(G233gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n461_), .B(KEYINPUT81), .Z(new_n462_));
  AOI21_X1  g261(.A(new_n458_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n460_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n462_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT30), .B1(new_n453_), .B2(new_n353_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n360_), .A2(new_n455_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n457_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n465_), .B1(new_n468_), .B2(new_n459_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n451_), .B1(new_n464_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n462_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n465_), .A3(new_n459_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n450_), .A3(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(KEYINPUT82), .A3(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G127gat), .B(G134gat), .Z(new_n475_));
  XOR2_X1   g274(.A(G113gat), .B(G120gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n477_), .B(KEYINPUT31), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G29gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(G85gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT0), .B(G57gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  NAND2_X1  g283(.A1(G225gat), .A2(G233gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n419_), .A2(new_n477_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n477_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n415_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n419_), .A2(new_n477_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(KEYINPUT4), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n490_), .A2(new_n491_), .A3(new_n485_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n484_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n488_), .A2(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n484_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT94), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n494_), .A2(new_n484_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(new_n493_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n495_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n470_), .A2(KEYINPUT82), .A3(new_n473_), .A4(new_n478_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n480_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n449_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n369_), .A2(KEYINPUT32), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n385_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n379_), .A2(new_n381_), .A3(KEYINPUT32), .A4(new_n369_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT95), .B1(new_n509_), .B2(new_n502_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT93), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n369_), .B1(new_n365_), .B2(new_n373_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n511_), .B1(new_n375_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n484_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n485_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n490_), .A2(new_n491_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n492_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT33), .B1(new_n496_), .B2(new_n497_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT33), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n499_), .A2(new_n521_), .A3(new_n493_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n519_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n387_), .A2(KEYINPUT93), .A3(new_n374_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n513_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n496_), .A2(KEYINPUT94), .A3(new_n497_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n500_), .B1(new_n499_), .B2(new_n493_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n493_), .A2(new_n494_), .ZN(new_n528_));
  OAI22_X1  g327(.A1(new_n526_), .A2(new_n527_), .B1(new_n484_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT95), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n507_), .A2(new_n508_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n510_), .A2(new_n525_), .A3(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT88), .B1(new_n440_), .B2(new_n441_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n446_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n389_), .A2(new_n534_), .A3(new_n535_), .A4(new_n502_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n480_), .A2(new_n503_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n505_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G29gat), .B(G36gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G15gat), .B(G22gat), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G1gat), .B(G8gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT76), .B(G1gat), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n550_), .A2(G8gat), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n548_), .B(new_n549_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n549_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n552_), .B1(new_n550_), .B2(G8gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n554_), .B1(new_n555_), .B2(new_n547_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n542_), .B(new_n543_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT15), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n546_), .A2(new_n553_), .A3(new_n556_), .A4(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n553_), .A2(new_n556_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n544_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n553_), .A2(new_n557_), .A3(new_n556_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n557_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n564_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G169gat), .B(G197gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n569_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n541_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT34), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n582_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT72), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n544_), .B2(new_n268_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n584_), .B1(new_n587_), .B2(KEYINPUT71), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n546_), .A2(new_n558_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n587_), .B1(new_n589_), .B2(new_n268_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  OAI221_X1 g390(.A(new_n587_), .B1(KEYINPUT71), .B2(new_n584_), .C1(new_n589_), .C2(new_n268_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G190gat), .B(G218gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT74), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n593_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n596_), .B(KEYINPUT36), .Z(new_n601_));
  NOR2_X1   g400(.A1(new_n593_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n578_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n593_), .A2(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n593_), .A2(new_n599_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n577_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n560_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(new_n269_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT77), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT16), .ZN(new_n615_));
  XOR2_X1   g414(.A(G183gat), .B(G211gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT17), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n613_), .B(new_n619_), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n611_), .A2(KEYINPUT17), .A3(new_n618_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n608_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n297_), .A2(new_n576_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT96), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n502_), .A2(new_n550_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n628_), .A2(KEYINPUT38), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(KEYINPUT38), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n604_), .A2(new_n605_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n631_), .B1(new_n541_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n540_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n636_));
  OAI211_X1 g435(.A(KEYINPUT97), .B(new_n632_), .C1(new_n636_), .C2(new_n505_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n296_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n574_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n623_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n502_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n629_), .A2(new_n630_), .A3(new_n644_), .ZN(G1324gat));
  INV_X1    g444(.A(G8gat), .ZN(new_n646_));
  INV_X1    g445(.A(new_n389_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n626_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n638_), .A2(new_n647_), .A3(new_n641_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n638_), .A2(KEYINPUT98), .A3(new_n647_), .A4(new_n641_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  OAI21_X1  g453(.A(G8gat), .B1(new_n654_), .B2(KEYINPUT99), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI22_X1  g455(.A1(new_n653_), .A2(new_n656_), .B1(KEYINPUT99), .B2(new_n654_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(KEYINPUT99), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n658_), .B(new_n655_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n648_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT40), .B(new_n648_), .C1(new_n657_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  INV_X1    g463(.A(G15gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n626_), .A2(new_n665_), .A3(new_n635_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G15gat), .B1(new_n643_), .B2(new_n540_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  INV_X1    g471(.A(new_n536_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n626_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G22gat), .B1(new_n643_), .B2(new_n536_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(new_n676_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(G1327gat));
  NOR2_X1   g478(.A1(new_n622_), .A2(new_n632_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n296_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n576_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n529_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n541_), .B2(new_n607_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n687_), .B(new_n608_), .C1(new_n636_), .C2(new_n505_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n639_), .A2(new_n574_), .A3(new_n623_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  AOI211_X1 g492(.A(new_n693_), .B(new_n690_), .C1(new_n686_), .C2(new_n688_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n529_), .A2(G29gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n685_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(KEYINPUT102), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n692_), .A2(new_n694_), .A3(new_n389_), .ZN(new_n701_));
  INV_X1    g500(.A(G36gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT101), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n689_), .A2(new_n691_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n693_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n689_), .A2(KEYINPUT44), .A3(new_n691_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n647_), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(G36gat), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n703_), .A2(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n389_), .A2(G36gat), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n683_), .A2(KEYINPUT45), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT45), .B1(new_n683_), .B2(new_n712_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(KEYINPUT46), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n700_), .B1(new_n710_), .B2(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n699_), .B(new_n717_), .C1(new_n703_), .C2(new_n709_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  NAND3_X1  g520(.A1(new_n695_), .A2(G43gat), .A3(new_n635_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n683_), .A2(new_n540_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(G43gat), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g524(.A(G50gat), .B1(new_n684_), .B2(new_n673_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n673_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n695_), .B2(new_n727_), .ZN(G1331gat));
  NAND2_X1  g527(.A1(new_n622_), .A2(new_n575_), .ZN(new_n729_));
  AOI211_X1 g528(.A(new_n729_), .B(new_n297_), .C1(new_n637_), .C2(new_n634_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G57gat), .B1(new_n731_), .B2(new_n502_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n541_), .A2(new_n574_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n296_), .A3(new_n624_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n247_), .A3(new_n529_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n732_), .A2(new_n736_), .ZN(G1332gat));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n245_), .A3(new_n647_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G64gat), .B1(new_n731_), .B2(new_n389_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(KEYINPUT48), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(KEYINPUT48), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n738_), .B1(new_n740_), .B2(new_n741_), .ZN(G1333gat));
  NAND3_X1  g541(.A1(new_n735_), .A2(new_n236_), .A3(new_n635_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G71gat), .B1(new_n731_), .B2(new_n540_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(KEYINPUT49), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(KEYINPUT49), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n743_), .B1(new_n745_), .B2(new_n746_), .ZN(G1334gat));
  NAND3_X1  g546(.A1(new_n735_), .A2(new_n238_), .A3(new_n673_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G78gat), .B1(new_n731_), .B2(new_n536_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT50), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(KEYINPUT50), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(G1335gat));
  NOR3_X1   g551(.A1(new_n639_), .A2(new_n574_), .A3(new_n622_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n689_), .A2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754_), .B2(new_n502_), .ZN(new_n755_));
  NOR4_X1   g554(.A1(new_n297_), .A2(new_n541_), .A3(new_n574_), .A4(new_n681_), .ZN(new_n756_));
  INV_X1    g555(.A(G85gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n529_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(G1336gat));
  AOI21_X1  g558(.A(G92gat), .B1(new_n756_), .B2(new_n647_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT103), .ZN(new_n761_));
  INV_X1    g560(.A(new_n754_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n389_), .A2(new_n203_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT104), .Z(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n762_), .B2(new_n764_), .ZN(G1337gat));
  AND3_X1   g564(.A1(new_n635_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n756_), .A2(new_n766_), .B1(KEYINPUT105), .B2(KEYINPUT51), .ZN(new_n767_));
  OAI21_X1  g566(.A(G99gat), .B1(new_n754_), .B2(new_n540_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n769_), .B(new_n770_), .Z(G1338gat));
  NAND3_X1  g570(.A1(new_n756_), .A2(new_n217_), .A3(new_n673_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n689_), .A2(new_n673_), .A3(new_n753_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(G106gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G106gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT107), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n772_), .B(new_n779_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT106), .B(KEYINPUT53), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n778_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1339gat));
  NAND3_X1  g583(.A1(new_n607_), .A2(new_n575_), .A3(new_n622_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(KEYINPUT108), .B(KEYINPUT54), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n639_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n787_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n296_), .B2(new_n785_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n259_), .B(new_n270_), .C1(new_n277_), .C2(new_n279_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n273_), .B1(new_n235_), .B2(new_n258_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT12), .B1(new_n268_), .B2(new_n269_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n235_), .A2(new_n258_), .A3(new_n278_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n793_), .A2(new_n274_), .B1(new_n797_), .B2(KEYINPUT55), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n797_), .A2(new_n799_), .A3(KEYINPUT55), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT110), .B1(new_n280_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n285_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n285_), .A2(KEYINPUT56), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n799_), .B1(new_n797_), .B2(KEYINPUT55), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n280_), .A2(KEYINPUT110), .A3(new_n801_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n807_), .B1(new_n814_), .B2(new_n798_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT111), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n806_), .A2(new_n811_), .A3(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n574_), .A2(KEYINPUT109), .A3(new_n288_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT109), .B1(new_n574_), .B2(new_n288_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n559_), .A2(new_n561_), .A3(new_n564_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n564_), .B1(new_n561_), .B2(new_n565_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n572_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n562_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(KEYINPUT112), .A3(new_n573_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n822_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n569_), .A2(new_n573_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n289_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT114), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n830_), .A2(new_n289_), .A3(new_n835_), .A4(new_n832_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n817_), .A2(new_n820_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n792_), .B1(new_n837_), .B2(new_n633_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n632_), .A2(KEYINPUT57), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT115), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n830_), .A2(new_n288_), .A3(new_n832_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n803_), .B2(new_n285_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n815_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n841_), .B(KEYINPUT58), .C1(new_n815_), .C2(new_n842_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n608_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n287_), .B1(new_n814_), .B2(new_n798_), .ZN(new_n848_));
  OAI22_X1  g647(.A1(KEYINPUT111), .A2(new_n815_), .B1(new_n848_), .B2(KEYINPUT56), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n809_), .A2(new_n810_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n820_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n834_), .A2(new_n836_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854_));
  INV_X1    g653(.A(new_n839_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n838_), .A2(new_n840_), .A3(new_n847_), .A4(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n791_), .B1(new_n857_), .B2(new_n623_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n449_), .A2(new_n540_), .A3(new_n502_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861_), .B2(new_n574_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT116), .ZN(new_n863_));
  INV_X1    g662(.A(new_n791_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n840_), .A2(new_n856_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n633_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n847_), .B1(new_n866_), .B2(KEYINPUT57), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n623_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT117), .B1(new_n857_), .B2(new_n623_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n864_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n860_), .A2(KEYINPUT59), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n868_), .A2(new_n864_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n859_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n872_), .A2(new_n873_), .B1(KEYINPUT59), .B2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(G113gat), .A3(new_n574_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n863_), .A2(new_n877_), .ZN(G1340gat));
  XNOR2_X1  g677(.A(KEYINPUT118), .B(G120gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n297_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n876_), .B2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n639_), .B2(KEYINPUT60), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(KEYINPUT60), .B2(new_n879_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n875_), .A2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT119), .B1(new_n881_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n879_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n875_), .A2(KEYINPUT59), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n854_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n888_));
  AOI211_X1 g687(.A(KEYINPUT115), .B(new_n839_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n574_), .A2(new_n288_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT109), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n574_), .A2(KEYINPUT109), .A3(new_n288_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT111), .B1(new_n803_), .B2(new_n808_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n842_), .A2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n897_), .B2(new_n816_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n834_), .A2(new_n836_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n632_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n607_), .B1(new_n844_), .B2(new_n843_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n900_), .A2(new_n792_), .B1(new_n846_), .B2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n622_), .B1(new_n890_), .B2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT117), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n868_), .A2(new_n869_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n791_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n873_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n887_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n886_), .B1(new_n908_), .B2(new_n297_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n910_));
  INV_X1    g709(.A(new_n884_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n885_), .A2(new_n912_), .ZN(G1341gat));
  OAI21_X1  g712(.A(G127gat), .B1(new_n908_), .B2(new_n623_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n623_), .A2(G127gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n875_), .B2(new_n915_), .ZN(G1342gat));
  AOI21_X1  g715(.A(G134gat), .B1(new_n861_), .B2(new_n633_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n608_), .A2(G134gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT120), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n876_), .B2(new_n919_), .ZN(G1343gat));
  NOR3_X1   g719(.A1(new_n536_), .A2(new_n647_), .A3(new_n502_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n858_), .A2(new_n635_), .A3(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n574_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n880_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G148gat), .ZN(G1345gat));
  OAI211_X1 g726(.A(new_n540_), .B(new_n921_), .C1(new_n903_), .C2(new_n791_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT121), .B1(new_n928_), .B2(new_n623_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n858_), .A2(new_n635_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n930_), .A2(new_n931_), .A3(new_n622_), .A4(new_n921_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n933_));
  AND3_X1   g732(.A1(new_n929_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n929_), .B2(new_n932_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT61), .B(G155gat), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n934_), .A2(new_n935_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n931_), .B1(new_n923_), .B2(new_n622_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n928_), .A2(KEYINPUT121), .A3(new_n623_), .ZN(new_n940_));
  OAI21_X1  g739(.A(KEYINPUT122), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n929_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n936_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n938_), .A2(new_n943_), .ZN(G1346gat));
  NAND3_X1  g743(.A1(new_n923_), .A2(G162gat), .A3(new_n608_), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n874_), .A2(new_n540_), .A3(new_n633_), .A4(new_n921_), .ZN(new_n946_));
  INV_X1    g745(.A(G162gat), .ZN(new_n947_));
  AND3_X1   g746(.A1(new_n946_), .A2(KEYINPUT123), .A3(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(KEYINPUT123), .B1(new_n946_), .B2(new_n947_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n945_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(KEYINPUT124), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n952_), .B(new_n945_), .C1(new_n948_), .C2(new_n949_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1347gat));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n673_), .A2(new_n504_), .A3(new_n389_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n906_), .A2(new_n575_), .A3(new_n957_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n955_), .B1(new_n958_), .B2(new_n349_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n872_), .A2(new_n574_), .A3(new_n956_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n960_), .A2(KEYINPUT125), .A3(G169gat), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n959_), .A2(KEYINPUT62), .A3(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(KEYINPUT125), .B1(new_n960_), .B2(G169gat), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n963_), .A2(new_n964_), .B1(new_n313_), .B2(new_n958_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n962_), .A2(new_n965_), .ZN(G1348gat));
  NOR2_X1   g765(.A1(new_n858_), .A2(new_n957_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n967_), .A2(G176gat), .A3(new_n880_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(KEYINPUT126), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n906_), .A2(new_n957_), .ZN(new_n970_));
  AOI21_X1  g769(.A(G176gat), .B1(new_n970_), .B2(new_n296_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n969_), .A2(new_n971_), .ZN(G1349gat));
  AOI21_X1  g771(.A(new_n347_), .B1(new_n967_), .B2(new_n622_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n623_), .A2(new_n337_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n973_), .B1(new_n970_), .B2(new_n974_), .ZN(G1350gat));
  NAND3_X1  g774(.A1(new_n970_), .A2(new_n336_), .A3(new_n633_), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n906_), .A2(new_n607_), .A3(new_n957_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n977_), .B2(new_n325_), .ZN(G1351gat));
  NOR3_X1   g777(.A1(new_n536_), .A2(new_n389_), .A3(new_n529_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n930_), .A2(new_n979_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n980_), .A2(new_n575_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(KEYINPUT127), .B(G197gat), .ZN(new_n982_));
  XNOR2_X1  g781(.A(new_n981_), .B(new_n982_), .ZN(G1352gat));
  INV_X1    g782(.A(new_n980_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n984_), .A2(new_n880_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n985_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g785(.A1(new_n980_), .A2(new_n623_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n988_));
  AND2_X1   g787(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n987_), .B1(new_n988_), .B2(new_n989_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n990_), .B1(new_n987_), .B2(new_n988_), .ZN(G1354gat));
  OR3_X1    g790(.A1(new_n980_), .A2(G218gat), .A3(new_n632_), .ZN(new_n992_));
  OAI21_X1  g791(.A(G218gat), .B1(new_n980_), .B2(new_n607_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n992_), .A2(new_n993_), .ZN(G1355gat));
endmodule


