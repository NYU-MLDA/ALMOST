//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT67), .B(KEYINPUT6), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n209_), .A2(KEYINPUT67), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(KEYINPUT67), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n206_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n204_), .A2(new_n208_), .A3(new_n212_), .ZN(new_n213_));
  AND2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(G85gat), .B2(G92gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G92gat), .Z(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G85gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT9), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n216_), .B1(new_n219_), .B2(KEYINPUT66), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221_));
  INV_X1    g020(.A(new_n218_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(G92gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n221_), .B1(new_n224_), .B2(KEYINPUT9), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n213_), .B1(new_n220_), .B2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n212_), .A2(new_n208_), .A3(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G85gat), .A2(G92gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n214_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n235_), .A2(KEYINPUT8), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n231_), .A2(new_n238_), .A3(new_n233_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(KEYINPUT8), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n226_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G29gat), .B(G36gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G43gat), .B(G50gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n231_), .A2(new_n238_), .A3(new_n233_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n238_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n241_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n220_), .A2(new_n225_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n213_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n245_), .B(KEYINPUT15), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n246_), .B(new_n255_), .C1(KEYINPUT35), .C2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(KEYINPUT35), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G190gat), .B(G218gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G134gat), .B(G162gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT36), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n261_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n264_), .B(KEYINPUT36), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n266_), .A2(new_n269_), .A3(KEYINPUT37), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n267_), .B(KEYINPUT74), .Z(new_n271_));
  NOR2_X1   g070(.A1(new_n261_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT37), .B1(new_n266_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G57gat), .B(G64gat), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n275_), .A2(KEYINPUT11), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(KEYINPUT11), .ZN(new_n277_));
  XOR2_X1   g076(.A(G71gat), .B(G78gat), .Z(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n277_), .A2(new_n278_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G231gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G1gat), .B(G8gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G15gat), .ZN(new_n287_));
  INV_X1    g086(.A(G22gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G15gat), .A2(G22gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G1gat), .A2(G8gat), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n289_), .A2(new_n290_), .B1(KEYINPUT14), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n286_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n283_), .B(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G127gat), .B(G155gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT16), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G183gat), .B(G211gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT17), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n298_), .A2(new_n299_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n294_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n294_), .A2(new_n300_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n274_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n308_), .A2(new_n311_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G155gat), .B(G162gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n309_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(new_n306_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n319_), .B(new_n320_), .C1(new_n315_), .C2(KEYINPUT1), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G113gat), .B(G120gat), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n323_), .A2(new_n324_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n323_), .B(new_n324_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(new_n321_), .A3(new_n317_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n330_), .A3(KEYINPUT4), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n322_), .A2(new_n327_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n331_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n328_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT91), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n328_), .A2(new_n330_), .A3(KEYINPUT91), .A4(new_n332_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G29gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G85gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(KEYINPUT0), .B(G57gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n336_), .A2(new_n339_), .A3(new_n345_), .A4(new_n340_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G183gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT25), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G183gat), .ZN(new_n353_));
  INV_X1    g152(.A(G190gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT26), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT26), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G190gat), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n351_), .A2(new_n353_), .A3(new_n355_), .A4(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(KEYINPUT24), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(G183gat), .B2(G190gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(G183gat), .A3(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT78), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n369_), .A2(new_n365_), .A3(G183gat), .A4(G190gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n366_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n366_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n367_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G169gat), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n364_), .A2(new_n372_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT30), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n327_), .A2(KEYINPUT31), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n327_), .A2(KEYINPUT31), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n383_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n383_), .A2(new_n387_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n381_), .A2(new_n382_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(G71gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(G99gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(G15gat), .B(G43gat), .Z(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT79), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n394_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n390_), .A2(new_n397_), .ZN(new_n398_));
  OR3_X1    g197(.A1(new_n388_), .A2(new_n389_), .A3(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n349_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT19), .ZN(new_n403_));
  INV_X1    g202(.A(G197gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT82), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G197gat), .ZN(new_n407_));
  INV_X1    g206(.A(G204gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT21), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(G197gat), .B2(G204gat), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n409_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n410_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G218gat), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n416_), .A2(G211gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(G211gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G197gat), .A2(G204gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT82), .B(G197gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(new_n408_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n420_), .B1(new_n424_), .B2(new_n411_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT21), .B1(new_n417_), .B2(new_n418_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n405_), .A2(new_n407_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n421_), .B1(new_n427_), .B2(G204gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n428_), .B2(KEYINPUT84), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n430_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n415_), .A2(new_n425_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT20), .B1(new_n432_), .B2(new_n380_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n409_), .A2(new_n412_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT83), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n408_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n411_), .B1(new_n436_), .B2(new_n421_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n409_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n435_), .A2(new_n437_), .A3(new_n419_), .A4(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(KEYINPUT84), .B(new_n422_), .C1(new_n423_), .C2(new_n408_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n426_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n431_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n379_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n358_), .A2(KEYINPUT87), .A3(new_n361_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n363_), .B1(new_n373_), .B2(new_n367_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT87), .B1(new_n358_), .B2(new_n361_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n444_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n403_), .B1(new_n433_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT95), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n453_), .B(new_n403_), .C1(new_n433_), .C2(new_n450_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT89), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n444_), .A2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(KEYINPUT89), .B(new_n379_), .C1(new_n371_), .C2(new_n375_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n459_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n362_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(KEYINPUT88), .A3(new_n445_), .A4(new_n446_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n443_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n403_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n432_), .B2(new_n380_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n452_), .A2(new_n454_), .A3(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G8gat), .B(G36gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(G64gat), .B(G92gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT27), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n465_), .A2(new_n468_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n456_), .A2(new_n457_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n479_), .A2(new_n432_), .A3(new_n460_), .A4(new_n463_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n377_), .A2(new_n379_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n363_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n358_), .A2(new_n361_), .A3(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n371_), .B2(new_n483_), .ZN(new_n484_));
  AOI211_X1 g283(.A(new_n467_), .B(new_n403_), .C1(new_n443_), .C2(new_n484_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n478_), .A2(new_n403_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n475_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n477_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n466_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n467_), .B1(new_n443_), .B2(new_n484_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n480_), .A2(new_n466_), .A3(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n475_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n485_), .A2(new_n480_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT20), .B1(new_n443_), .B2(new_n484_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n479_), .A2(new_n460_), .A3(new_n463_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n494_), .B1(new_n443_), .B2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n493_), .B(new_n487_), .C1(new_n496_), .C2(new_n466_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n497_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n476_), .A2(new_n488_), .B1(new_n498_), .B2(new_n477_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n322_), .A2(KEYINPUT29), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G22gat), .B(G50gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT28), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n500_), .B(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G228gat), .A2(G233gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI221_X4 g304(.A(new_n505_), .B1(new_n322_), .B2(KEYINPUT29), .C1(new_n439_), .C2(new_n442_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n322_), .A2(KEYINPUT29), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n504_), .B1(new_n443_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n506_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n503_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT86), .ZN(new_n514_));
  INV_X1    g313(.A(new_n507_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n505_), .B1(new_n432_), .B2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n443_), .A2(new_n504_), .A3(new_n507_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n509_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n513_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n514_), .B1(new_n513_), .B2(new_n519_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n512_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n518_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT86), .B1(new_n510_), .B2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n500_), .B(new_n502_), .Z(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n519_), .B2(KEYINPUT85), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n513_), .A2(new_n519_), .A3(new_n514_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n524_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n401_), .A2(new_n499_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT96), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n488_), .A2(new_n476_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n498_), .A2(new_n477_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n349_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n522_), .A2(new_n535_), .A3(new_n528_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n531_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n522_), .A2(new_n535_), .A3(new_n528_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n499_), .A2(new_n538_), .A3(KEYINPUT96), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n487_), .A2(KEYINPUT32), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n470_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n493_), .B1(new_n496_), .B2(new_n466_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n349_), .B1(new_n543_), .B2(new_n541_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n348_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT92), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n328_), .A2(new_n330_), .A3(new_n333_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n346_), .A2(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT93), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n331_), .A2(new_n332_), .A3(new_n335_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n331_), .A2(KEYINPUT94), .A3(new_n332_), .A4(new_n335_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(KEYINPUT93), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n551_), .A2(new_n554_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n348_), .A2(new_n545_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n348_), .A2(KEYINPUT92), .A3(new_n545_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n548_), .A2(new_n557_), .A3(new_n558_), .A4(new_n559_), .ZN(new_n560_));
  OAI22_X1  g359(.A1(new_n542_), .A2(new_n544_), .B1(new_n560_), .B2(new_n498_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n529_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n537_), .A2(new_n539_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n399_), .A2(new_n400_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n530_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n281_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT12), .B1(new_n567_), .B2(KEYINPUT70), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n569_), .B(new_n570_), .C1(new_n242_), .C2(new_n281_), .ZN(new_n571_));
  AND2_X1   g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n242_), .B2(new_n281_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n568_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT71), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n281_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT69), .B1(new_n253_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT69), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n242_), .A2(new_n579_), .A3(new_n281_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n572_), .B1(new_n581_), .B2(new_n567_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n568_), .A2(new_n571_), .A3(KEYINPUT71), .A4(new_n573_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n576_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT5), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n576_), .A2(new_n582_), .A3(new_n583_), .A4(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT13), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(KEYINPUT72), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(KEYINPUT72), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n592_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n592_), .A2(new_n595_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n293_), .B(new_n245_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n293_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n254_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n293_), .A2(new_n245_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n603_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n601_), .B1(new_n610_), .B2(KEYINPUT76), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(KEYINPUT76), .B2(new_n610_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n605_), .A2(new_n609_), .A3(new_n601_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT77), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n605_), .A2(KEYINPUT77), .A3(new_n609_), .A4(new_n601_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n612_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR4_X1   g418(.A1(new_n305_), .A2(new_n566_), .A3(new_n598_), .A4(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(G1gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n349_), .B(KEYINPUT97), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n620_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT38), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n563_), .A2(new_n565_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n530_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n266_), .A2(new_n269_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n628_), .A2(KEYINPUT98), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT98), .B1(new_n628_), .B2(new_n630_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n598_), .A2(new_n619_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n304_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n633_), .A2(new_n535_), .A3(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n625_), .B1(new_n621_), .B2(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(G8gat), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n633_), .A2(new_n635_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(new_n534_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n620_), .A2(new_n638_), .A3(new_n534_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(KEYINPUT40), .A3(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1325gat));
  NAND2_X1  g447(.A1(new_n639_), .A2(new_n564_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(G15gat), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n633_), .A2(new_n565_), .A3(new_n635_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT99), .B1(new_n652_), .B2(new_n287_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(KEYINPUT41), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n620_), .A2(new_n287_), .A3(new_n564_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(new_n651_), .B2(new_n653_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1326gat));
  INV_X1    g457(.A(new_n529_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n288_), .B1(new_n639_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT42), .Z(new_n661_));
  NAND3_X1  g460(.A1(new_n620_), .A2(new_n288_), .A3(new_n659_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1327gat));
  NOR2_X1   g462(.A1(new_n566_), .A2(new_n619_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n304_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n629_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n598_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n349_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT100), .B1(new_n566_), .B2(new_n274_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n634_), .A2(new_n665_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n270_), .A2(new_n273_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n499_), .A2(new_n538_), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n677_), .A2(new_n531_), .B1(new_n529_), .B2(new_n561_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n564_), .B1(new_n678_), .B2(new_n539_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n679_), .B2(new_n530_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n675_), .B1(new_n680_), .B2(KEYINPUT100), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n675_), .B1(new_n566_), .B2(new_n274_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n672_), .B(new_n674_), .C1(new_n681_), .C2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n671_), .A2(KEYINPUT101), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n683_), .A3(new_n682_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n689_), .A2(KEYINPUT44), .A3(new_n672_), .A4(new_n674_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n623_), .A2(G29gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n670_), .B1(new_n692_), .B2(new_n693_), .ZN(G1328gat));
  NAND3_X1  g493(.A1(new_n687_), .A2(new_n534_), .A3(new_n690_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G36gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n499_), .A2(G36gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n664_), .A2(new_n667_), .A3(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT45), .Z(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n696_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT102), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n699_), .B1(new_n695_), .B2(G36gat), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(KEYINPUT46), .ZN(new_n706_));
  AND4_X1   g505(.A1(KEYINPUT103), .A2(new_n696_), .A3(KEYINPUT46), .A4(new_n700_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT103), .B1(new_n704_), .B2(KEYINPUT46), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n703_), .A2(new_n706_), .B1(new_n707_), .B2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(G43gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n565_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n692_), .A2(KEYINPUT104), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n668_), .B2(new_n565_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n714_));
  INV_X1    g513(.A(new_n711_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n691_), .B2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n712_), .A2(new_n713_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT47), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n712_), .A2(new_n719_), .A3(new_n716_), .A4(new_n713_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1330gat));
  NAND3_X1  g520(.A1(new_n692_), .A2(G50gat), .A3(new_n659_), .ZN(new_n722_));
  INV_X1    g521(.A(G50gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n723_), .B1(new_n668_), .B2(new_n529_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT105), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n722_), .A2(new_n727_), .A3(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1331gat));
  OR2_X1    g528(.A1(new_n596_), .A2(new_n597_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n305_), .A2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT106), .Z(new_n732_));
  NOR2_X1   g531(.A1(new_n566_), .A2(new_n618_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n623_), .ZN(new_n735_));
  INV_X1    g534(.A(G57gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n598_), .A2(new_n619_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(new_n665_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n739_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT107), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n742_), .B(new_n739_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n741_), .A2(G57gat), .A3(new_n349_), .A4(new_n743_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n744_), .A2(KEYINPUT108), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(KEYINPUT108), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n737_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT109), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n737_), .A2(new_n745_), .A3(new_n749_), .A4(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1332gat));
  INV_X1    g550(.A(G64gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n734_), .A2(new_n752_), .A3(new_n534_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n741_), .A2(new_n534_), .A3(new_n743_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n755_), .A3(G64gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G64gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(G1333gat));
  NAND3_X1  g557(.A1(new_n734_), .A2(new_n392_), .A3(new_n564_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n741_), .A2(new_n564_), .A3(new_n743_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(G71gat), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G71gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1334gat));
  INV_X1    g563(.A(G78gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n734_), .A2(new_n765_), .A3(new_n659_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n741_), .A2(new_n659_), .A3(new_n743_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n767_), .A2(new_n768_), .A3(G78gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n767_), .B2(G78gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT111), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n766_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n738_), .A2(new_n304_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n689_), .A2(new_n672_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n349_), .A2(new_n218_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n730_), .A2(new_n666_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n733_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(new_n622_), .ZN(new_n781_));
  OAI22_X1  g580(.A1(new_n777_), .A2(new_n778_), .B1(G85gat), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT112), .ZN(G1336gat));
  NOR3_X1   g582(.A1(new_n777_), .A2(new_n223_), .A3(new_n499_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n780_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G92gat), .B1(new_n785_), .B2(new_n534_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n777_), .B2(new_n565_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n202_), .A3(new_n564_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(KEYINPUT113), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n790_), .B(new_n792_), .ZN(G1338gat));
  NAND3_X1  g592(.A1(new_n785_), .A2(new_n203_), .A3(new_n659_), .ZN(new_n794_));
  OAI21_X1  g593(.A(G106gat), .B1(new_n777_), .B2(new_n529_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n795_), .A2(KEYINPUT52), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(G106gat), .C1(new_n777_), .C2(new_n529_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n794_), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n794_), .B(new_n801_), .C1(new_n796_), .C2(new_n799_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1339gat));
  NOR2_X1   g604(.A1(new_n534_), .A2(new_n659_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n564_), .A3(new_n623_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT57), .B1(new_n266_), .B2(new_n269_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n618_), .A2(new_n591_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n574_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n568_), .A2(new_n571_), .A3(new_n578_), .A4(new_n580_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n811_), .A2(KEYINPUT55), .B1(new_n812_), .B2(new_n572_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n576_), .A2(new_n814_), .A3(new_n583_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n588_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(KEYINPUT56), .A3(new_n588_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n810_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n607_), .A2(new_n608_), .A3(new_n604_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n601_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n615_), .A2(new_n616_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n592_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n809_), .B1(new_n821_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT117), .ZN(new_n828_));
  INV_X1    g627(.A(new_n810_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT56), .B1(new_n816_), .B2(new_n588_), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n818_), .B(new_n590_), .C1(new_n813_), .C2(new_n815_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n829_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n825_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n809_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n824_), .A2(new_n591_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n836_), .A2(KEYINPUT116), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(KEYINPUT116), .ZN(new_n838_));
  OAI221_X1 g637(.A(KEYINPUT58), .B1(new_n830_), .B2(new_n831_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n839_));
  OAI22_X1  g638(.A1(new_n837_), .A2(new_n838_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n274_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n828_), .A2(new_n835_), .B1(new_n839_), .B2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n629_), .B1(new_n832_), .B2(new_n825_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT115), .B1(new_n844_), .B2(KEYINPUT57), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n821_), .A2(new_n826_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n846_), .B(new_n847_), .C1(new_n848_), .C2(new_n629_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n843_), .A2(KEYINPUT118), .A3(new_n845_), .A4(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n845_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n840_), .A2(new_n841_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n839_), .A3(new_n676_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n834_), .B1(new_n833_), .B2(new_n809_), .ZN(new_n855_));
  AOI211_X1 g654(.A(KEYINPUT117), .B(new_n808_), .C1(new_n832_), .C2(new_n825_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n851_), .B1(new_n852_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n850_), .A2(new_n858_), .A3(new_n665_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n730_), .A2(new_n304_), .A3(new_n619_), .A4(new_n274_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n807_), .B1(new_n859_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n847_), .B1(new_n848_), .B2(new_n629_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n304_), .B1(new_n843_), .B2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n862_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n807_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n865_), .ZN(new_n870_));
  OAI22_X1  g669(.A1(new_n864_), .A2(new_n865_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G113gat), .B1(new_n871_), .B2(new_n619_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n828_), .A2(new_n835_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n873_), .A2(new_n854_), .A3(new_n845_), .A4(new_n849_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n304_), .B1(new_n874_), .B2(new_n851_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n862_), .B1(new_n875_), .B2(new_n850_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT119), .B1(new_n876_), .B2(new_n807_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n864_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n619_), .A2(G113gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n877_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n872_), .A2(new_n881_), .ZN(G1340gat));
  OAI21_X1  g681(.A(G120gat), .B1(new_n871_), .B2(new_n730_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n884_));
  AOI21_X1  g683(.A(G120gat), .B1(new_n598_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n884_), .B2(G120gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n877_), .A2(new_n879_), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n887_), .ZN(G1341gat));
  OAI21_X1  g687(.A(G127gat), .B1(new_n871_), .B2(new_n665_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n665_), .A2(G127gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n877_), .A2(new_n879_), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1342gat));
  OAI21_X1  g691(.A(G134gat), .B1(new_n871_), .B2(new_n274_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n630_), .A2(G134gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n877_), .A2(new_n879_), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1343gat));
  NAND3_X1  g695(.A1(new_n565_), .A2(new_n659_), .A3(new_n623_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n534_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n859_), .B2(new_n863_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n618_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n598_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n876_), .A2(KEYINPUT120), .A3(new_n665_), .A4(new_n899_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n900_), .B2(new_n304_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n859_), .A2(new_n863_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n304_), .A3(new_n898_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT120), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n900_), .A2(new_n908_), .A3(new_n304_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n914_), .A3(new_n905_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n910_), .A2(new_n915_), .ZN(G1346gat));
  AOI21_X1  g715(.A(G162gat), .B1(new_n900_), .B2(new_n629_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n676_), .A2(G162gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT121), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n900_), .B2(new_n919_), .ZN(G1347gat));
  NAND3_X1  g719(.A1(new_n564_), .A2(new_n534_), .A3(new_n622_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT122), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n619_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n659_), .B1(new_n924_), .B2(KEYINPUT123), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(KEYINPUT123), .B2(new_n924_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G169gat), .B1(new_n868_), .B2(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT62), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n923_), .A2(new_n659_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n868_), .B2(new_n931_), .ZN(new_n932_));
  OAI211_X1 g731(.A(KEYINPUT124), .B(new_n930_), .C1(new_n867_), .C2(new_n862_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n935_));
  AND2_X1   g734(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n618_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n928_), .B1(new_n934_), .B2(new_n937_), .ZN(G1348gat));
  INV_X1    g737(.A(G176gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n939_), .B1(new_n934_), .B2(new_n730_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n730_), .A2(new_n939_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n911_), .A2(new_n930_), .A3(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(KEYINPUT125), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n876_), .A2(new_n931_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n944_), .A2(new_n945_), .A3(new_n941_), .ZN(new_n946_));
  AND3_X1   g745(.A1(new_n940_), .A2(new_n943_), .A3(new_n946_), .ZN(G1349gat));
  AOI21_X1  g746(.A(G183gat), .B1(new_n944_), .B2(new_n304_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n934_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n665_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n948_), .B1(new_n949_), .B2(new_n950_), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n934_), .B2(new_n274_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n629_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n934_), .B2(new_n953_), .ZN(G1351gat));
  NOR3_X1   g753(.A1(new_n564_), .A2(new_n499_), .A3(new_n536_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n911_), .A2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(G197gat), .B1(new_n957_), .B2(new_n618_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n956_), .A2(new_n404_), .A3(new_n619_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1352gat));
  NAND3_X1  g759(.A1(new_n957_), .A2(new_n408_), .A3(new_n598_), .ZN(new_n961_));
  OAI21_X1  g760(.A(G204gat), .B1(new_n956_), .B2(new_n730_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1353gat));
  XNOR2_X1  g762(.A(KEYINPUT63), .B(G211gat), .ZN(new_n964_));
  NOR3_X1   g763(.A1(new_n956_), .A2(new_n665_), .A3(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n957_), .A2(new_n304_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(G1354gat));
  NOR3_X1   g767(.A1(new_n956_), .A2(new_n416_), .A3(new_n274_), .ZN(new_n969_));
  INV_X1    g768(.A(new_n955_), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n876_), .A2(new_n630_), .A3(new_n970_), .ZN(new_n971_));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n972_));
  AOI21_X1  g771(.A(G218gat), .B1(new_n971_), .B2(new_n972_), .ZN(new_n973_));
  OAI21_X1  g772(.A(KEYINPUT126), .B1(new_n956_), .B2(new_n630_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n969_), .B1(new_n973_), .B2(new_n974_), .ZN(G1355gat));
endmodule


