//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n215_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT65), .B1(new_n217_), .B2(KEYINPUT9), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n219_), .A3(new_n214_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n216_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n210_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT66), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G57gat), .B(G64gat), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n226_));
  XOR2_X1   g025(.A(G71gat), .B(G78gat), .Z(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n226_), .A2(new_n227_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n209_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT69), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT70), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT67), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT7), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT7), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(new_n237_), .B2(KEYINPUT67), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n233_), .A2(new_n245_), .A3(new_n234_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n236_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n213_), .A2(new_n215_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n231_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  AOI211_X1 g049(.A(KEYINPUT8), .B(new_n248_), .C1(new_n244_), .C2(new_n209_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n223_), .B(new_n230_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n244_), .A2(new_n209_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(new_n231_), .A3(new_n249_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n243_), .B1(new_n235_), .B2(KEYINPUT70), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n248_), .B1(new_n256_), .B2(new_n246_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n257_), .B2(new_n231_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n230_), .B1(new_n258_), .B2(new_n223_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT12), .B1(new_n253_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT64), .Z(new_n262_));
  OAI21_X1  g061(.A(new_n223_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n230_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT12), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n260_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n253_), .A2(new_n259_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n267_), .B(new_n268_), .C1(new_n262_), .C2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT12), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n264_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(new_n252_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n262_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n273_), .A2(new_n274_), .A3(new_n265_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n269_), .A2(new_n262_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G120gat), .B(G148gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT5), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G176gat), .B(G204gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n281_), .B(KEYINPUT72), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n270_), .A2(new_n277_), .A3(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n275_), .A2(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n281_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT13), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n285_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT73), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT37), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G232gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT34), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT35), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n297_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G29gat), .B(G36gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G43gat), .B(G50gat), .Z(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G43gat), .B(G50gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n299_), .B1(new_n263_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT15), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n303_), .A2(KEYINPUT15), .A3(new_n305_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(new_n258_), .B2(new_n223_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n298_), .B1(new_n308_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n263_), .A2(new_n312_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n258_), .A2(new_n223_), .A3(new_n306_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n298_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .A4(new_n299_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n293_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G190gat), .B(G218gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(G134gat), .B(G162gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT36), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n324_), .A2(KEYINPUT36), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n320_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  AOI221_X4 g128(.A(new_n293_), .B1(new_n329_), .B2(new_n325_), .C1(new_n315_), .C2(new_n319_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n292_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n320_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n326_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(new_n329_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n330_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT37), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G231gat), .A2(G233gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n230_), .B(new_n338_), .Z(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT75), .B(G1gat), .ZN(new_n340_));
  INV_X1    g139(.A(G8gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT14), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G15gat), .B(G22gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G8gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n339_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G127gat), .B(G155gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G183gat), .B(G211gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT17), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n350_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n355_), .B(KEYINPUT17), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n357_), .B1(new_n350_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n337_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n291_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT86), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(KEYINPUT86), .A2(G169gat), .A3(G176gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT24), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT23), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(G183gat), .A3(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n369_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(KEYINPUT24), .B2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n370_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT84), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT26), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(G190gat), .ZN(new_n381_));
  INV_X1    g180(.A(G190gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(KEYINPUT26), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT85), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n379_), .A2(new_n381_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT83), .B(G183gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT25), .ZN(new_n387_));
  INV_X1    g186(.A(new_n383_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT85), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n382_), .A2(KEYINPUT26), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT25), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n390_), .A2(KEYINPUT84), .B1(new_n391_), .B2(G183gat), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .A4(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT88), .ZN(new_n394_));
  AND2_X1   g193(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n395_));
  NOR2_X1   g194(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n394_), .B(G169gat), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(G169gat), .B1(new_n395_), .B2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT88), .ZN(new_n399_));
  INV_X1    g198(.A(G169gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(G176gat), .B1(new_n400_), .B2(KEYINPUT22), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n386_), .A2(new_n382_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n367_), .B1(new_n403_), .B2(new_n375_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n378_), .A2(new_n393_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G71gat), .B(G99gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(G15gat), .B(G43gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  XNOR2_X1  g207(.A(new_n405_), .B(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G127gat), .B(G134gat), .Z(new_n410_));
  XOR2_X1   g209(.A(G113gat), .B(G120gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n409_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n415_), .B(KEYINPUT89), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT30), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT31), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n414_), .B(new_n418_), .Z(new_n419_));
  NAND2_X1  g218(.A1(G228gat), .A2(G233gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G78gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G106gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G22gat), .B(G50gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G155gat), .A2(G162gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT90), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT1), .ZN(new_n429_));
  NAND3_X1  g228(.A1(KEYINPUT90), .A2(G155gat), .A3(G162gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT91), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT91), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n428_), .A2(new_n433_), .A3(new_n429_), .A4(new_n430_), .ZN(new_n434_));
  OR2_X1    g233(.A1(G155gat), .A2(G162gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n430_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT90), .B1(G155gat), .B2(G162gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT1), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n432_), .A2(new_n434_), .A3(new_n435_), .A4(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G141gat), .A2(G148gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G141gat), .A2(G148gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n442_), .B(KEYINPUT3), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n440_), .B(KEYINPUT2), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT28), .B1(new_n450_), .B2(KEYINPUT29), .ZN(new_n451_));
  INV_X1    g250(.A(G204gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G197gat), .ZN(new_n453_));
  INV_X1    g252(.A(G197gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G204gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT21), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT93), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G211gat), .B(G218gat), .Z(new_n460_));
  NAND2_X1  g259(.A1(new_n453_), .A2(KEYINPUT92), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT92), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(new_n452_), .A3(G197gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n463_), .A3(new_n455_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n460_), .B1(new_n464_), .B2(KEYINPUT21), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n459_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n453_), .A2(new_n455_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n460_), .A2(KEYINPUT21), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n448_), .B1(new_n439_), .B2(new_n443_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT29), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT28), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n473_), .A3(new_n471_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n451_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n451_), .B2(new_n474_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n425_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n477_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(new_n475_), .A3(new_n424_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n419_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G8gat), .B(G36gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G64gat), .B(G92gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n367_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(KEYINPUT24), .A3(new_n376_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n377_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n393_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n402_), .A2(new_n404_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n469_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT25), .B(G183gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(new_n363_), .A3(new_n376_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT95), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT95), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n375_), .B1(new_n497_), .B2(new_n376_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT22), .B(G169gat), .ZN(new_n506_));
  INV_X1    g305(.A(G176gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n488_), .A2(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(G183gat), .A2(G190gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n375_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT96), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n375_), .A2(KEYINPUT96), .A3(new_n510_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n509_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n468_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n459_), .B2(new_n465_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n505_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G226gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT19), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AND4_X1   g321(.A1(KEYINPUT20), .A2(new_n494_), .A3(new_n519_), .A4(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n496_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n501_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n524_), .A2(new_n525_), .A3(new_n503_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n469_), .B1(new_n526_), .B2(new_n515_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT20), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n405_), .B2(new_n518_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n522_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n487_), .B1(new_n523_), .B2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT20), .B1(new_n493_), .B2(new_n469_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n518_), .B1(new_n505_), .B2(new_n516_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n521_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n487_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n494_), .A2(new_n519_), .A3(KEYINPUT20), .A4(new_n522_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(KEYINPUT98), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT27), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT98), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n534_), .A2(new_n540_), .A3(new_n535_), .A4(new_n536_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n527_), .A2(new_n529_), .A3(new_n522_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n494_), .A2(new_n519_), .A3(KEYINPUT20), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n543_), .B1(new_n544_), .B2(new_n522_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n487_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(KEYINPUT27), .A3(new_n537_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n482_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G225gat), .A2(G233gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n450_), .A2(new_n413_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT99), .B1(new_n470_), .B2(new_n412_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT99), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n470_), .A2(new_n556_), .A3(new_n412_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n552_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n444_), .A2(new_n449_), .A3(new_n412_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n556_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n470_), .A2(new_n412_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT4), .B1(new_n563_), .B2(new_n557_), .ZN(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT100), .B(KEYINPUT4), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n552_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n559_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G1gat), .B(G29gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G57gat), .B(G85gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n555_), .A2(new_n558_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n567_), .B1(new_n577_), .B2(KEYINPUT4), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n576_), .B1(new_n578_), .B2(new_n559_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n550_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n481_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n535_), .A2(KEYINPUT32), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n523_), .B2(new_n530_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n545_), .B2(new_n583_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n564_), .A2(new_n568_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n559_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n574_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n578_), .A2(new_n559_), .A3(new_n576_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n585_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT104), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT104), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n580_), .A2(new_n592_), .A3(new_n585_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n574_), .B1(new_n577_), .B2(new_n552_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n566_), .A2(new_n551_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT102), .B1(new_n564_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT4), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT102), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n596_), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT103), .B(new_n595_), .C1(new_n598_), .C2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n569_), .B2(new_n574_), .ZN(new_n605_));
  NOR4_X1   g404(.A1(new_n578_), .A2(KEYINPUT33), .A3(new_n559_), .A4(new_n576_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n603_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n538_), .A2(new_n541_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n577_), .A2(new_n552_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n576_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n564_), .A2(KEYINPUT102), .A3(new_n597_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n601_), .B1(new_n600_), .B2(new_n596_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n608_), .B1(new_n613_), .B2(KEYINPUT103), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n607_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n582_), .B1(new_n594_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT105), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n575_), .A2(new_n579_), .A3(new_n481_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n548_), .B2(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n575_), .A2(new_n579_), .A3(new_n481_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n620_), .A2(KEYINPUT105), .A3(new_n542_), .A4(new_n547_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n581_), .B1(new_n623_), .B2(new_n419_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n310_), .A2(new_n347_), .A3(new_n348_), .A4(new_n311_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n347_), .A2(new_n348_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT77), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n306_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n303_), .A2(KEYINPUT77), .A3(new_n305_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT78), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n628_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n631_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT77), .B1(new_n303_), .B2(new_n305_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT78), .B1(new_n637_), .B2(new_n349_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n627_), .B(KEYINPUT79), .C1(new_n634_), .C2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n637_), .A2(new_n349_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n633_), .B1(new_n628_), .B2(new_n632_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n637_), .A2(new_n349_), .A3(KEYINPUT78), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n640_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n626_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n625_), .A2(new_n626_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(KEYINPUT79), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT80), .B1(new_n644_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT79), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n634_), .A2(new_n638_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(new_n645_), .ZN(new_n651_));
  OAI22_X1  g450(.A1(new_n634_), .A2(new_n638_), .B1(new_n637_), .B2(new_n349_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n626_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT80), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n651_), .A2(new_n654_), .A3(new_n655_), .A4(new_n639_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G113gat), .B(G141gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G169gat), .B(G197gat), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n657_), .B(new_n658_), .Z(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n648_), .A2(new_n656_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT81), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n651_), .A2(new_n654_), .A3(new_n639_), .A4(new_n659_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT82), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n652_), .A2(new_n653_), .B1(new_n646_), .B2(KEYINPUT79), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(KEYINPUT82), .A3(new_n651_), .A4(new_n659_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT81), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n648_), .A2(new_n656_), .A3(new_n670_), .A4(new_n660_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n663_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n624_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n362_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n580_), .A2(KEYINPUT106), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n580_), .A2(KEYINPUT106), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n676_), .A2(new_n340_), .A3(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT38), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n328_), .A2(new_n330_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n624_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n285_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT13), .B1(new_n283_), .B2(new_n285_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n673_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n360_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n685_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n688_), .A2(KEYINPUT107), .A3(new_n689_), .A4(new_n360_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n580_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G1gat), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n681_), .A2(new_n696_), .ZN(G1324gat));
  NAND3_X1  g496(.A1(new_n676_), .A2(new_n341_), .A3(new_n548_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n684_), .A2(new_n692_), .A3(new_n693_), .A4(new_n548_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT39), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(G8gat), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n700_), .B1(new_n699_), .B2(G8gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n698_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT108), .B(KEYINPUT40), .Z(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1325gat));
  OAI21_X1  g505(.A(G15gat), .B1(new_n694_), .B2(new_n419_), .ZN(new_n707_));
  XOR2_X1   g506(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT110), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  OR3_X1    g509(.A1(new_n675_), .A2(G15gat), .A3(new_n419_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n709_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(G1326gat));
  NAND4_X1  g512(.A1(new_n684_), .A2(new_n692_), .A3(new_n693_), .A4(new_n481_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(G22gat), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n714_), .B2(G22gat), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n582_), .A2(G22gat), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n717_), .A2(new_n718_), .B1(new_n675_), .B2(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT112), .Z(G1327gat));
  NOR2_X1   g520(.A1(new_n682_), .A2(new_n360_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n688_), .A2(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n674_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G29gat), .B1(new_n724_), .B2(new_n580_), .ZN(new_n725_));
  XOR2_X1   g524(.A(KEYINPUT113), .B(KEYINPUT43), .Z(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n331_), .A2(new_n336_), .A3(KEYINPUT114), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT114), .B1(new_n331_), .B2(new_n336_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n727_), .B1(new_n624_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n337_), .A2(KEYINPUT43), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n624_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n419_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n616_), .B2(new_n622_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT115), .B(new_n733_), .C1(new_n737_), .C2(new_n581_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n731_), .A2(new_n735_), .A3(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n690_), .A2(new_n360_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(KEYINPUT44), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT44), .B1(new_n739_), .B2(new_n740_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n679_), .A2(G29gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n725_), .B1(new_n743_), .B2(new_n744_), .ZN(G1328gat));
  INV_X1    g544(.A(G36gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n724_), .A2(new_n746_), .A3(new_n548_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT45), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n724_), .A2(new_n749_), .A3(new_n746_), .A4(new_n548_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n741_), .A2(new_n742_), .A3(new_n549_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n746_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n751_), .B(KEYINPUT46), .C1(new_n752_), .C2(new_n746_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1329gat));
  NAND2_X1  g556(.A1(new_n736_), .A2(G43gat), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n741_), .A2(new_n742_), .A3(new_n758_), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT116), .B(G43gat), .Z(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n724_), .B2(new_n736_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n759_), .A2(KEYINPUT47), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT47), .B1(new_n759_), .B2(new_n761_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1330gat));
  AOI21_X1  g563(.A(G50gat), .B1(new_n724_), .B2(new_n481_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n481_), .A2(G50gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n743_), .B2(new_n766_), .ZN(G1331gat));
  NOR2_X1   g566(.A1(new_n624_), .A2(new_n689_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n688_), .A2(new_n361_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G57gat), .B1(new_n770_), .B2(new_n679_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT117), .Z(new_n772_));
  INV_X1    g571(.A(new_n291_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n662_), .A2(new_n669_), .A3(new_n671_), .A4(new_n360_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n684_), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT118), .B(G57gat), .Z(new_n777_));
  NOR3_X1   g576(.A1(new_n776_), .A2(new_n695_), .A3(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n772_), .A2(new_n778_), .ZN(G1332gat));
  INV_X1    g578(.A(new_n770_), .ZN(new_n780_));
  OR3_X1    g579(.A1(new_n780_), .A2(G64gat), .A3(new_n549_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n775_), .A2(new_n548_), .A3(new_n684_), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n783_));
  AND3_X1   g582(.A1(new_n782_), .A2(G64gat), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n782_), .B2(G64gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1333gat));
  OAI21_X1  g585(.A(G71gat), .B1(new_n776_), .B2(new_n419_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT49), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n419_), .A2(G71gat), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT120), .Z(new_n790_));
  OAI21_X1  g589(.A(new_n788_), .B1(new_n780_), .B2(new_n790_), .ZN(G1334gat));
  OR3_X1    g590(.A1(new_n780_), .A2(G78gat), .A3(new_n582_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G78gat), .B1(new_n776_), .B2(new_n582_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(KEYINPUT50), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(KEYINPUT50), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n792_), .B1(new_n794_), .B2(new_n795_), .ZN(G1335gat));
  AND2_X1   g595(.A1(new_n291_), .A2(new_n722_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n768_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(new_n211_), .A3(new_n679_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n290_), .A2(new_n673_), .A3(new_n691_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n739_), .A2(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(new_n580_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n804_), .B2(new_n211_), .ZN(G1336gat));
  NAND3_X1  g604(.A1(new_n799_), .A2(new_n212_), .A3(new_n548_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n803_), .A2(new_n548_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n212_), .ZN(G1337gat));
  NAND4_X1  g607(.A1(new_n797_), .A2(new_n202_), .A3(new_n736_), .A4(new_n768_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT121), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n803_), .A2(new_n736_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G99gat), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT51), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n810_), .A2(new_n815_), .A3(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1338gat));
  NAND3_X1  g616(.A1(new_n799_), .A2(new_n203_), .A3(new_n481_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n739_), .A2(new_n481_), .A3(new_n802_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n819_), .A2(new_n820_), .A3(G106gat), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n819_), .B2(G106gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT53), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n818_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1339gat));
  INV_X1    g626(.A(new_n679_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n550_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n672_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n662_), .A4(new_n360_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n774_), .A2(KEYINPUT122), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n337_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT123), .B1(new_n834_), .B2(new_n290_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n774_), .B(new_n831_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n688_), .A2(new_n836_), .A3(new_n837_), .A4(new_n337_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n835_), .A2(new_n838_), .A3(KEYINPUT54), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n285_), .B1(new_n663_), .B2(new_n672_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n267_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n274_), .B1(new_n273_), .B2(new_n265_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n260_), .A2(new_n266_), .A3(KEYINPUT55), .A4(new_n262_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT56), .B1(new_n849_), .B2(new_n282_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n275_), .A2(KEYINPUT55), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n847_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT56), .B(new_n282_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n844_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n625_), .A2(new_n653_), .ZN(new_n856_));
  OAI221_X1 g655(.A(new_n660_), .B1(new_n650_), .B2(new_n856_), .C1(new_n653_), .C2(new_n643_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n669_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n682_), .B1(new_n855_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n858_), .B1(new_n284_), .B2(new_n281_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n854_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n850_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n337_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n862_), .B(KEYINPUT58), .C1(new_n863_), .C2(new_n850_), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n860_), .A2(new_n861_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT57), .B(new_n682_), .C1(new_n855_), .C2(new_n859_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n360_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n829_), .B1(new_n843_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(G113gat), .B1(new_n872_), .B2(new_n689_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n871_), .A2(KEYINPUT59), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(KEYINPUT59), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n871_), .A2(KEYINPUT124), .A3(KEYINPUT59), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n874_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n689_), .A2(G113gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n873_), .B1(new_n879_), .B2(new_n880_), .ZN(G1340gat));
  INV_X1    g680(.A(G120gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n688_), .B2(KEYINPUT60), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n872_), .B(new_n883_), .C1(KEYINPUT60), .C2(new_n882_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n291_), .B1(new_n871_), .B2(KEYINPUT59), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n886_), .B2(new_n882_), .ZN(G1341gat));
  OAI211_X1 g686(.A(new_n360_), .B(new_n829_), .C1(new_n843_), .C2(new_n870_), .ZN(new_n888_));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n888_), .A2(KEYINPUT125), .A3(new_n889_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n691_), .A2(new_n889_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n879_), .B2(new_n895_), .ZN(G1342gat));
  AOI21_X1  g695(.A(G134gat), .B1(new_n872_), .B2(new_n683_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n337_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n898_), .A2(G134gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n879_), .B2(new_n899_), .ZN(G1343gat));
  OR2_X1    g699(.A1(new_n843_), .A2(new_n870_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n828_), .A2(new_n736_), .A3(new_n582_), .A4(new_n548_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n689_), .A3(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g703(.A1(new_n901_), .A2(new_n291_), .A3(new_n902_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g705(.A1(new_n901_), .A2(new_n360_), .A3(new_n902_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT61), .B(G155gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1346gat));
  NAND2_X1  g708(.A1(new_n901_), .A2(new_n902_), .ZN(new_n910_));
  INV_X1    g709(.A(G162gat), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n910_), .A2(new_n911_), .A3(new_n730_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n901_), .A2(new_n683_), .A3(new_n902_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n911_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT126), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n913_), .A2(new_n916_), .A3(new_n911_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n912_), .B1(new_n915_), .B2(new_n917_), .ZN(G1347gat));
  NAND3_X1  g717(.A1(new_n828_), .A2(new_n482_), .A3(new_n548_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n901_), .A2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G169gat), .B1(new_n921_), .B2(new_n673_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  OAI211_X1 g723(.A(KEYINPUT62), .B(G169gat), .C1(new_n921_), .C2(new_n673_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n843_), .A2(new_n870_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n919_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n927_), .A2(new_n689_), .A3(new_n506_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n924_), .A2(new_n925_), .A3(new_n928_), .ZN(G1348gat));
  OAI21_X1  g728(.A(G176gat), .B1(new_n921_), .B2(new_n773_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n927_), .A2(new_n507_), .A3(new_n290_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1349gat));
  NAND2_X1  g731(.A1(new_n927_), .A2(new_n360_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n495_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n386_), .B2(new_n933_), .ZN(G1350gat));
  AOI21_X1  g734(.A(new_n382_), .B1(new_n927_), .B2(new_n898_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n682_), .A2(new_n383_), .A3(new_n381_), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n901_), .A2(new_n920_), .A3(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(KEYINPUT127), .B1(new_n936_), .B2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n901_), .A2(new_n898_), .A3(new_n920_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(G190gat), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n927_), .A2(new_n937_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n939_), .A2(new_n944_), .ZN(G1351gat));
  NOR4_X1   g744(.A1(new_n549_), .A2(new_n736_), .A3(new_n580_), .A4(new_n582_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n901_), .A2(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n673_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n454_), .ZN(G1352gat));
  NOR2_X1   g748(.A1(new_n947_), .A2(new_n773_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(new_n452_), .ZN(G1353gat));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n947_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n953_), .B1(new_n954_), .B2(new_n360_), .ZN(new_n955_));
  AND2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  NOR4_X1   g755(.A1(new_n947_), .A2(new_n691_), .A3(new_n952_), .A4(new_n956_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n955_), .A2(new_n957_), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n947_), .B2(new_n337_), .ZN(new_n959_));
  OR2_X1    g758(.A1(new_n682_), .A2(G218gat), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n947_), .B2(new_n960_), .ZN(G1355gat));
endmodule


