//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n987_, new_n988_, new_n990_, new_n991_,
    new_n992_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1010_, new_n1011_, new_n1012_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  AND2_X1   g003(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n205_));
  AND2_X1   g004(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n207_));
  NOR3_X1   g006(.A1(new_n206_), .A2(new_n207_), .A3(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT9), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT9), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n217_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n218_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n214_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G36gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G29gat), .ZN(new_n226_));
  INV_X1    g025(.A(G29gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G36gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G50gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G43gat), .ZN(new_n231_));
  INV_X1    g030(.A(G43gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G50gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n229_), .A2(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n226_), .A2(new_n228_), .A3(new_n231_), .A4(new_n233_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238_));
  INV_X1    g037(.A(G99gat), .ZN(new_n239_));
  INV_X1    g038(.A(G106gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n241_), .A2(new_n211_), .A3(new_n212_), .A4(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n215_), .A2(new_n216_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT8), .ZN(new_n246_));
  INV_X1    g045(.A(G85gat), .ZN(new_n247_));
  INV_X1    g046(.A(G92gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT65), .A3(new_n219_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n245_), .A2(new_n246_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n246_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(new_n244_), .A3(new_n243_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n224_), .A2(new_n237_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n252_), .A2(new_n244_), .A3(new_n243_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n244_), .B2(new_n243_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n259_), .A2(KEYINPUT69), .A3(new_n237_), .A4(new_n224_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT15), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT15), .B1(new_n235_), .B2(new_n236_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n251_), .A2(new_n253_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n206_), .A2(new_n207_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n211_), .B(new_n212_), .C1(new_n266_), .C2(G106gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n223_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n217_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n264_), .B1(new_n265_), .B2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n256_), .A2(new_n260_), .A3(new_n261_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G232gat), .A2(G233gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT34), .Z(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n224_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n255_), .A2(new_n254_), .B1(new_n276_), .B2(new_n264_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n274_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n277_), .A2(new_n261_), .A3(new_n260_), .A4(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n275_), .A2(KEYINPUT35), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT35), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n281_), .A3(new_n260_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n282_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n205_), .B1(new_n280_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(new_n280_), .B2(new_n283_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  OAI221_X1 g088(.A(new_n285_), .B1(new_n287_), .B2(new_n205_), .C1(new_n280_), .C2(new_n283_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT102), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G134gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G127gat), .ZN(new_n296_));
  INV_X1    g095(.A(G127gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G134gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G120gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G113gat), .ZN(new_n301_));
  INV_X1    g100(.A(G113gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G120gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G113gat), .B(G120gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT3), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT2), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n312_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n315_), .A2(KEYINPUT1), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n315_), .B1(new_n316_), .B2(KEYINPUT1), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n324_), .B2(KEYINPUT85), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(G155gat), .B2(G162gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT85), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n315_), .ZN(new_n329_));
  AOI211_X1 g128(.A(KEYINPUT86), .B(new_n322_), .C1(new_n325_), .C2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n324_), .A2(KEYINPUT85), .ZN(new_n332_));
  INV_X1    g131(.A(new_n323_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n329_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n322_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n331_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n309_), .B(new_n318_), .C1(new_n330_), .C2(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n327_), .A2(new_n328_), .A3(new_n315_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n328_), .B1(new_n327_), .B2(new_n315_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n323_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT86), .B1(new_n341_), .B2(new_n322_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n334_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n338_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT82), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n299_), .A2(new_n304_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(KEYINPUT82), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT83), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n306_), .A2(new_n307_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT82), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n308_), .A2(new_n345_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n349_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n337_), .B(KEYINPUT4), .C1(new_n344_), .C2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n349_), .A2(new_n354_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n318_), .B1(new_n330_), .B2(new_n336_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT94), .Z(new_n362_));
  NAND3_X1  g161(.A1(new_n356_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n337_), .B(new_n361_), .C1(new_n344_), .C2(new_n355_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT96), .ZN(new_n366_));
  XOR2_X1   g165(.A(G1gat), .B(G29gat), .Z(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n366_), .B(new_n367_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n369_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n363_), .A2(new_n364_), .A3(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT98), .B(KEYINPUT33), .Z(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT99), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n370_), .A2(new_n373_), .A3(KEYINPUT33), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n363_), .A2(new_n364_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT97), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT97), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n363_), .A2(new_n381_), .A3(new_n384_), .A4(new_n364_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G8gat), .B(G36gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G169gat), .ZN(new_n393_));
  INV_X1    g192(.A(G176gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(KEYINPUT91), .A2(KEYINPUT24), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(KEYINPUT91), .A2(KEYINPUT24), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n395_), .B(new_n396_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(G190gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT26), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT26), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(G190gat), .ZN(new_n404_));
  AND2_X1   g203(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n405_));
  NOR2_X1   g204(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n402_), .B(new_n404_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n399_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G169gat), .A2(G176gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n397_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n400_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT81), .B1(new_n412_), .B2(KEYINPUT23), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(KEYINPUT23), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT23), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(G183gat), .A3(G190gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n413_), .B1(new_n417_), .B2(KEYINPUT81), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n393_), .A2(KEYINPUT22), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT22), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G169gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n421_), .A3(new_n394_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n396_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(G183gat), .A2(G190gat), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n425_));
  OAI22_X1  g224(.A1(new_n411_), .A2(new_n418_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(G197gat), .A2(G204gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G197gat), .A2(G204gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT21), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(KEYINPUT21), .A3(new_n428_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G211gat), .B(G218gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n432_), .A2(new_n433_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT20), .B1(new_n426_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n418_), .ZN(new_n439_));
  AND2_X1   g238(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(G190gat), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n423_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n395_), .A2(KEYINPUT24), .A3(new_n396_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT24), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n409_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n417_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(KEYINPUT79), .A2(KEYINPUT26), .ZN(new_n450_));
  NOR2_X1   g249(.A1(KEYINPUT79), .A2(KEYINPUT26), .ZN(new_n451_));
  OAI21_X1  g250(.A(G190gat), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT80), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n454_), .B(G190gat), .C1(new_n450_), .C2(new_n451_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT25), .B1(new_n440_), .B2(new_n441_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n406_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n457_), .A2(new_n458_), .B1(KEYINPUT26), .B2(new_n401_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n449_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n436_), .B1(new_n445_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G226gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT19), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n438_), .A2(new_n461_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n456_), .A2(new_n459_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n449_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n436_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n396_), .B(new_n422_), .C1(new_n418_), .C2(new_n443_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT20), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n426_), .B2(new_n436_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n464_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT92), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n465_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AOI211_X1 g275(.A(KEYINPUT92), .B(new_n464_), .C1(new_n471_), .C2(new_n473_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n392_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n356_), .A2(new_n361_), .A3(new_n360_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n337_), .B(new_n362_), .C1(new_n344_), .C2(new_n355_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n374_), .A3(new_n480_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n445_), .A2(new_n460_), .A3(new_n436_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n426_), .A2(new_n436_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT20), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n463_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT92), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n474_), .A2(new_n475_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(new_n391_), .A3(new_n487_), .A4(new_n465_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n478_), .A2(new_n481_), .A3(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n376_), .A2(KEYINPUT99), .A3(new_n377_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n380_), .A2(new_n386_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n471_), .A2(new_n464_), .A3(new_n473_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n468_), .A2(new_n470_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n437_), .B1(new_n493_), .B2(new_n436_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n494_), .B2(new_n464_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n391_), .A2(KEYINPUT32), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n486_), .A2(new_n487_), .A3(new_n465_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n376_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n375_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n500_));
  OAI221_X1 g299(.A(new_n497_), .B1(new_n498_), .B2(new_n496_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n491_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n436_), .B1(new_n344_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G228gat), .A2(G233gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT89), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n469_), .B1(new_n358_), .B2(KEYINPUT29), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n506_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G78gat), .B(G106gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n508_), .A2(new_n510_), .A3(KEYINPUT90), .A4(new_n511_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n511_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n509_), .A2(new_n506_), .ZN(new_n517_));
  AOI211_X1 g316(.A(new_n469_), .B(new_n507_), .C1(new_n358_), .C2(KEYINPUT29), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n503_), .B(new_n318_), .C1(new_n330_), .C2(new_n336_), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n342_), .A2(new_n343_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n521_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n523_), .A2(new_n503_), .A3(new_n318_), .A4(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G22gat), .B(G50gat), .Z(new_n526_));
  AND3_X1   g325(.A1(new_n522_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n514_), .A2(new_n515_), .A3(new_n519_), .A4(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT88), .B1(new_n527_), .B2(new_n528_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n522_), .A2(new_n525_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n526_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n522_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n517_), .A2(new_n518_), .A3(new_n516_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n511_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n531_), .B(new_n537_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G71gat), .B(G99gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(new_n232_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT31), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G227gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(G15gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT30), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n493_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n468_), .A2(new_n470_), .A3(new_n548_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n355_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n355_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n544_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n552_), .A3(new_n543_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n530_), .A2(new_n540_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n502_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n499_), .A2(new_n500_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n478_), .A2(new_n488_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT27), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n495_), .A2(KEYINPUT100), .A3(new_n392_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT100), .B1(new_n495_), .B2(new_n392_), .ZN(new_n568_));
  OAI211_X1 g367(.A(KEYINPUT27), .B(new_n488_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n530_), .A2(new_n540_), .A3(new_n558_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n558_), .B1(new_n530_), .B2(new_n540_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n563_), .B(new_n570_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n562_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n294_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT103), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT101), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT68), .ZN(new_n578_));
  XOR2_X1   g377(.A(G57gat), .B(G64gat), .Z(new_n579_));
  INV_X1    g378(.A(KEYINPUT11), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT66), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT66), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(KEYINPUT11), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .A4(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n583_), .B1(new_n584_), .B2(KEYINPUT11), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n584_), .A2(new_n585_), .A3(KEYINPUT11), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n585_), .B1(new_n584_), .B2(KEYINPUT11), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n276_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n578_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n587_), .A2(new_n591_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n259_), .A2(new_n597_), .A3(new_n224_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(KEYINPUT68), .A3(new_n594_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n592_), .A2(new_n276_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT12), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT12), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n592_), .A2(new_n276_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n598_), .A2(KEYINPUT67), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT67), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n259_), .A2(new_n597_), .A3(new_n607_), .A4(new_n224_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n608_), .A3(new_n601_), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n600_), .A2(new_n605_), .B1(new_n595_), .B2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT5), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n610_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n610_), .A2(new_n615_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT13), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n616_), .A2(KEYINPUT13), .A3(new_n617_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G15gat), .B(G22gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G1gat), .A2(G8gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT14), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(G1gat), .ZN(new_n628_));
  INV_X1    g427(.A(G8gat), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n625_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n624_), .A2(new_n625_), .A3(new_n630_), .A4(new_n626_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n264_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n237_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G229gat), .A2(G233gat), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n635_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G113gat), .B(G141gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G169gat), .B(G197gat), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n642_), .B(new_n643_), .Z(new_n644_));
  AND2_X1   g443(.A1(new_n235_), .A2(new_n236_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n634_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n636_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT74), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n646_), .A2(KEYINPUT74), .A3(new_n636_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT75), .B1(new_n651_), .B2(new_n639_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n646_), .A2(KEYINPUT74), .A3(new_n636_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT74), .B1(new_n646_), .B2(new_n636_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT75), .B(new_n639_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n641_), .B(new_n644_), .C1(new_n652_), .C2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT76), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n639_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT75), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n640_), .B1(new_n661_), .B2(new_n655_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT76), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n663_), .A3(new_n644_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n658_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(new_n655_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n644_), .B1(new_n666_), .B2(new_n641_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT77), .B1(new_n665_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT77), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n670_), .B(new_n667_), .C1(new_n658_), .C2(new_n664_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n577_), .B1(new_n623_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n634_), .B(KEYINPUT73), .ZN(new_n674_));
  NAND2_X1  g473(.A1(G231gat), .A2(G233gat), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(new_n592_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT17), .ZN(new_n678_));
  XOR2_X1   g477(.A(G127gat), .B(G155gat), .Z(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT16), .ZN(new_n680_));
  XNOR2_X1  g479(.A(G183gat), .B(G211gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  OR3_X1    g481(.A1(new_n677_), .A2(new_n678_), .A3(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(KEYINPUT17), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n677_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n672_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n622_), .A3(KEYINPUT101), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n673_), .A2(new_n687_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n576_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G1gat), .B1(new_n691_), .B2(new_n563_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n563_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n530_), .A2(new_n540_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n559_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n530_), .A2(new_n540_), .A3(new_n558_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n693_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n560_), .B1(new_n491_), .B2(new_n501_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(new_n672_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n289_), .A2(new_n290_), .A3(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n687_), .A2(new_n621_), .A3(new_n620_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n700_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n563_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n628_), .A3(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT38), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n692_), .A2(new_n709_), .ZN(G1324gat));
  INV_X1    g509(.A(KEYINPUT40), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n691_), .A2(new_n570_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n629_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT104), .B(G8gat), .C1(new_n691_), .C2(new_n570_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(KEYINPUT39), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n570_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n706_), .A2(new_n629_), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n714_), .B2(KEYINPUT39), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n711_), .B1(new_n717_), .B2(new_n720_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n714_), .A2(KEYINPUT39), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n722_), .A2(KEYINPUT40), .A3(new_n716_), .A4(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1325gat));
  OAI21_X1  g523(.A(G15gat), .B1(new_n691_), .B2(new_n559_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT41), .Z(new_n726_));
  NAND3_X1  g525(.A1(new_n706_), .A2(new_n546_), .A3(new_n558_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1326gat));
  INV_X1    g527(.A(new_n694_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G22gat), .B1(new_n691_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT42), .ZN(new_n731_));
  INV_X1    g530(.A(G22gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n706_), .A2(new_n732_), .A3(new_n694_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1327gat));
  AND3_X1   g533(.A1(new_n622_), .A2(new_n291_), .A3(new_n686_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n700_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G29gat), .B1(new_n737_), .B2(new_n707_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739_));
  INV_X1    g538(.A(new_n701_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n291_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n289_), .A2(new_n290_), .A3(new_n701_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n562_), .A2(new_n573_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n739_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n741_), .A2(new_n742_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n574_), .A2(new_n739_), .A3(new_n744_), .A4(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OAI22_X1  g547(.A1(new_n697_), .A2(new_n698_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(KEYINPUT43), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(KEYINPUT43), .ZN(new_n752_));
  OAI22_X1  g551(.A1(new_n745_), .A2(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n673_), .A2(new_n686_), .A3(new_n689_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n227_), .B(new_n563_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n753_), .A2(KEYINPUT44), .A3(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT107), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT105), .B1(new_n743_), .B2(new_n744_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n749_), .A2(new_n750_), .A3(KEYINPUT43), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT106), .B1(new_n749_), .B2(KEYINPUT43), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n747_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n754_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(KEYINPUT44), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n760_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n738_), .B1(new_n758_), .B2(new_n769_), .ZN(G1328gat));
  XOR2_X1   g569(.A(new_n570_), .B(KEYINPUT109), .Z(new_n771_));
  NOR3_X1   g570(.A1(new_n736_), .A2(G36gat), .A3(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT110), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT45), .Z(new_n774_));
  OAI21_X1  g573(.A(new_n718_), .B1(new_n766_), .B2(KEYINPUT44), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n760_), .B2(new_n768_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n225_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n570_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n767_), .B1(new_n766_), .B2(KEYINPUT44), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n761_), .A2(new_n762_), .B1(new_n764_), .B2(new_n747_), .ZN(new_n781_));
  NOR4_X1   g580(.A1(new_n781_), .A2(KEYINPUT107), .A3(new_n754_), .A4(new_n757_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n779_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT108), .B1(new_n783_), .B2(G36gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n774_), .B1(new_n778_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT46), .B(new_n774_), .C1(new_n778_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1329gat));
  AOI21_X1  g588(.A(G43gat), .B1(new_n737_), .B2(new_n558_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n232_), .B(new_n559_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n769_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g592(.A(G50gat), .B1(new_n737_), .B2(new_n694_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n230_), .B(new_n729_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n769_), .ZN(G1331gat));
  NOR2_X1   g595(.A1(new_n622_), .A2(new_n686_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n576_), .A2(new_n672_), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(G57gat), .A3(new_n707_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n799_), .A2(KEYINPUT112), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(KEYINPUT112), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n699_), .A2(new_n688_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT111), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n803_), .A2(new_n704_), .A3(new_n797_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G57gat), .B1(new_n804_), .B2(new_n707_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n800_), .A2(new_n801_), .A3(new_n805_), .ZN(G1332gat));
  INV_X1    g605(.A(G64gat), .ZN(new_n807_));
  INV_X1    g606(.A(new_n771_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT48), .Z(new_n810_));
  NAND3_X1  g609(.A1(new_n804_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1333gat));
  INV_X1    g611(.A(G71gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n798_), .B2(new_n558_), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n814_), .B(KEYINPUT49), .Z(new_n815_));
  NAND3_X1  g614(.A1(new_n804_), .A2(new_n813_), .A3(new_n558_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1334gat));
  INV_X1    g616(.A(G78gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n798_), .B2(new_n694_), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n819_), .B(KEYINPUT50), .Z(new_n820_));
  NAND3_X1  g619(.A1(new_n804_), .A2(new_n818_), .A3(new_n694_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1335gat));
  NOR2_X1   g621(.A1(new_n622_), .A2(new_n687_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n753_), .A2(new_n672_), .A3(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT113), .ZN(new_n825_));
  OAI21_X1  g624(.A(G85gat), .B1(new_n825_), .B2(new_n563_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n803_), .A2(new_n291_), .A3(new_n823_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n247_), .A3(new_n707_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1336gat));
  OAI21_X1  g628(.A(G92gat), .B1(new_n825_), .B2(new_n771_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n248_), .A3(new_n718_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1337gat));
  INV_X1    g631(.A(new_n266_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n827_), .A2(new_n558_), .A3(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n825_), .A2(new_n559_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n239_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT51), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n834_), .C1(new_n835_), .C2(new_n239_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1338gat));
  NAND3_X1  g639(.A1(new_n827_), .A2(new_n240_), .A3(new_n694_), .ZN(new_n841_));
  OAI21_X1  g640(.A(G106gat), .B1(new_n824_), .B2(new_n729_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(KEYINPUT52), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(KEYINPUT52), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g645(.A1(new_n705_), .A2(new_n704_), .A3(new_n672_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(KEYINPUT54), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n847_), .A2(KEYINPUT114), .A3(KEYINPUT54), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n847_), .A2(KEYINPUT115), .A3(KEYINPUT54), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT115), .B1(new_n847_), .B2(KEYINPUT54), .ZN(new_n853_));
  OAI22_X1  g652(.A1(new_n850_), .A2(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n604_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n603_), .B1(new_n592_), .B2(new_n276_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n606_), .B(new_n608_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n857_), .A2(new_n858_), .A3(new_n595_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n857_), .B2(new_n595_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861_));
  INV_X1    g660(.A(new_n599_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT68), .B1(new_n598_), .B2(new_n594_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n605_), .B(KEYINPUT55), .C1(new_n862_), .C2(new_n863_), .ZN(new_n864_));
  OAI22_X1  g663(.A1(new_n859_), .A2(new_n860_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n600_), .A2(new_n605_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n861_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n614_), .B1(new_n865_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT56), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n651_), .A2(new_n638_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n644_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n636_), .A2(new_n639_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n873_), .B(new_n874_), .C1(new_n635_), .C2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n665_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n617_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n880_), .B(new_n614_), .C1(new_n865_), .C2(new_n870_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n872_), .A2(new_n879_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(KEYINPUT119), .A3(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(KEYINPUT119), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n872_), .A2(new_n879_), .A3(new_n885_), .A4(new_n881_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(new_n746_), .A3(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n657_), .A2(KEYINPUT76), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n663_), .B1(new_n662_), .B2(new_n644_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n668_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n670_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n665_), .A2(KEYINPUT77), .A3(new_n668_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n878_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n857_), .A2(new_n595_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT116), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n857_), .A2(new_n858_), .A3(new_n595_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n864_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n895_), .A2(new_n896_), .B1(new_n897_), .B2(KEYINPUT117), .ZN(new_n898_));
  AOI21_X1  g697(.A(KEYINPUT55), .B1(new_n600_), .B2(new_n605_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n615_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n880_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n871_), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n893_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n877_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n291_), .B1(new_n905_), .B2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n887_), .B1(new_n908_), .B2(KEYINPUT57), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n910_));
  AOI211_X1 g709(.A(new_n910_), .B(new_n291_), .C1(new_n905_), .C2(new_n907_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n686_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n854_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n718_), .A2(new_n563_), .A3(new_n696_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n915_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT120), .B1(new_n909_), .B2(new_n911_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n617_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n919_));
  AOI21_X1  g718(.A(KEYINPUT56), .B1(new_n871_), .B2(KEYINPUT118), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n906_), .B1(new_n921_), .B2(new_n904_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n910_), .B1(new_n922_), .B2(new_n291_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n908_), .A2(KEYINPUT57), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .A4(new_n887_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n918_), .A2(new_n686_), .A3(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n917_), .B1(new_n927_), .B2(new_n854_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n916_), .B1(new_n928_), .B2(new_n914_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n916_), .B(KEYINPUT121), .C1(new_n928_), .C2(new_n914_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n931_), .A2(new_n688_), .A3(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G113gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n928_), .A2(new_n302_), .A3(new_n688_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1340gat));
  OAI21_X1  g735(.A(G120gat), .B1(new_n929_), .B2(new_n622_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n300_), .B1(new_n622_), .B2(KEYINPUT60), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n928_), .B(new_n938_), .C1(KEYINPUT60), .C2(new_n300_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(G1341gat));
  AOI21_X1  g739(.A(G127gat), .B1(new_n928_), .B2(new_n687_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n941_), .B(new_n942_), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n931_), .A2(G127gat), .A3(new_n687_), .A4(new_n932_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1342gat));
  NAND3_X1  g744(.A1(new_n931_), .A2(new_n746_), .A3(new_n932_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(G134gat), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n928_), .A2(new_n295_), .A3(new_n293_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1343gat));
  AOI21_X1  g748(.A(new_n695_), .B1(new_n927_), .B2(new_n854_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n950_), .A2(new_n707_), .A3(new_n771_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n951_), .A2(new_n672_), .ZN(new_n952_));
  XOR2_X1   g751(.A(KEYINPUT123), .B(G141gat), .Z(new_n953_));
  XNOR2_X1  g752(.A(new_n952_), .B(new_n953_), .ZN(G1344gat));
  INV_X1    g753(.A(new_n951_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n623_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g756(.A1(new_n955_), .A2(new_n687_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(KEYINPUT61), .B(G155gat), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n958_), .B(new_n959_), .ZN(G1346gat));
  OR3_X1    g759(.A1(new_n951_), .A2(G162gat), .A3(new_n294_), .ZN(new_n961_));
  OAI21_X1  g760(.A(G162gat), .B1(new_n951_), .B2(new_n704_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n771_), .A2(new_n707_), .ZN(new_n964_));
  INV_X1    g763(.A(new_n964_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n965_), .A2(new_n696_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n913_), .A2(new_n966_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G169gat), .B1(new_n967_), .B2(new_n672_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n969_));
  OR2_X1    g768(.A1(new_n968_), .A2(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n967_), .ZN(new_n971_));
  NAND4_X1  g770(.A1(new_n971_), .A2(new_n419_), .A3(new_n421_), .A4(new_n688_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n968_), .A2(new_n969_), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n970_), .A2(new_n972_), .A3(new_n973_), .ZN(G1348gat));
  AOI211_X1 g773(.A(new_n696_), .B(new_n965_), .C1(new_n927_), .C2(new_n854_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n622_), .A2(new_n394_), .ZN(new_n976_));
  AND3_X1   g775(.A1(new_n975_), .A2(KEYINPUT124), .A3(new_n976_), .ZN(new_n977_));
  AOI21_X1  g776(.A(KEYINPUT124), .B1(new_n975_), .B2(new_n976_), .ZN(new_n978_));
  AOI21_X1  g777(.A(G176gat), .B1(new_n971_), .B2(new_n623_), .ZN(new_n979_));
  NOR3_X1   g778(.A1(new_n977_), .A2(new_n978_), .A3(new_n979_), .ZN(G1349gat));
  AOI21_X1  g779(.A(new_n442_), .B1(new_n975_), .B2(new_n687_), .ZN(new_n981_));
  NOR4_X1   g780(.A1(new_n967_), .A2(new_n406_), .A3(new_n405_), .A4(new_n686_), .ZN(new_n982_));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n983_));
  OR3_X1    g782(.A1(new_n981_), .A2(new_n982_), .A3(new_n983_), .ZN(new_n984_));
  OAI21_X1  g783(.A(new_n983_), .B1(new_n981_), .B2(new_n982_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(G1350gat));
  OAI21_X1  g785(.A(G190gat), .B1(new_n967_), .B2(new_n704_), .ZN(new_n987_));
  NAND3_X1  g786(.A1(new_n293_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n988_));
  OAI21_X1  g787(.A(new_n987_), .B1(new_n967_), .B2(new_n988_), .ZN(G1351gat));
  INV_X1    g788(.A(new_n950_), .ZN(new_n990_));
  NOR2_X1   g789(.A1(new_n990_), .A2(new_n965_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n991_), .A2(new_n688_), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n992_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g792(.A1(new_n991_), .A2(new_n623_), .ZN(new_n994_));
  INV_X1    g793(.A(G204gat), .ZN(new_n995_));
  NOR2_X1   g794(.A1(new_n995_), .A2(KEYINPUT126), .ZN(new_n996_));
  AND2_X1   g795(.A1(new_n995_), .A2(KEYINPUT126), .ZN(new_n997_));
  OAI21_X1  g796(.A(new_n994_), .B1(new_n996_), .B2(new_n997_), .ZN(new_n998_));
  OAI21_X1  g797(.A(new_n998_), .B1(new_n994_), .B2(new_n996_), .ZN(G1353gat));
  INV_X1    g798(.A(KEYINPUT63), .ZN(new_n1000_));
  AOI21_X1  g799(.A(new_n686_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1001_));
  NAND3_X1  g800(.A1(new_n950_), .A2(new_n964_), .A3(new_n1001_), .ZN(new_n1002_));
  NAND2_X1  g801(.A1(new_n1002_), .A2(KEYINPUT127), .ZN(new_n1003_));
  INV_X1    g802(.A(G211gat), .ZN(new_n1004_));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n1005_));
  NAND4_X1  g804(.A1(new_n950_), .A2(new_n1005_), .A3(new_n964_), .A4(new_n1001_), .ZN(new_n1006_));
  AND4_X1   g805(.A1(new_n1000_), .A2(new_n1003_), .A3(new_n1004_), .A4(new_n1006_), .ZN(new_n1007_));
  AOI22_X1  g806(.A1(new_n1003_), .A2(new_n1006_), .B1(new_n1000_), .B2(new_n1004_), .ZN(new_n1008_));
  NOR2_X1   g807(.A1(new_n1007_), .A2(new_n1008_), .ZN(G1354gat));
  INV_X1    g808(.A(G218gat), .ZN(new_n1010_));
  NAND3_X1  g809(.A1(new_n991_), .A2(new_n1010_), .A3(new_n293_), .ZN(new_n1011_));
  NOR3_X1   g810(.A1(new_n990_), .A2(new_n704_), .A3(new_n965_), .ZN(new_n1012_));
  OAI21_X1  g811(.A(new_n1011_), .B1(new_n1010_), .B2(new_n1012_), .ZN(G1355gat));
endmodule


