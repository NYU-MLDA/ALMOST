//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G127gat), .B(G134gat), .Z(new_n203_));
  XOR2_X1   g002(.A(G113gat), .B(G120gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G127gat), .B(G134gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G113gat), .B(G120gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT31), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT84), .B1(new_n210_), .B2(KEYINPUT83), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(KEYINPUT84), .B2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(G183gat), .B2(G190gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n213_), .A2(KEYINPUT81), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n215_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n216_), .B1(new_n220_), .B2(KEYINPUT82), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n213_), .A2(KEYINPUT81), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT23), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT82), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT79), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n228_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(KEYINPUT79), .A3(new_n229_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n232_), .A2(new_n237_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n221_), .A2(new_n226_), .B1(new_n227_), .B2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n227_), .B1(G169gat), .B2(G176gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n232_), .A2(new_n237_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242_));
  INV_X1    g041(.A(G190gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT77), .B1(new_n243_), .B2(KEYINPUT26), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT25), .B(G183gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT26), .B(G190gat), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n244_), .B(new_n245_), .C1(new_n246_), .C2(KEYINPUT77), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n241_), .A2(new_n242_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n242_), .B1(new_n241_), .B2(new_n247_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n239_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(new_n234_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT23), .B1(new_n218_), .B2(new_n219_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n213_), .A2(new_n215_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n250_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT30), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G71gat), .B(G99gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n263_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G227gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(G15gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(G43gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n264_), .A2(new_n265_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n270_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n212_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n264_), .A2(new_n265_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n269_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(new_n211_), .A3(new_n271_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G85gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT0), .B(G57gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n209_), .A2(KEYINPUT4), .ZN(new_n283_));
  INV_X1    g082(.A(G155gat), .ZN(new_n284_));
  INV_X1    g083(.A(G162gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(KEYINPUT85), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT85), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(G155gat), .B2(G162gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT86), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n297_));
  INV_X1    g096(.A(G141gat), .ZN(new_n298_));
  INV_X1    g097(.A(G148gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT3), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT2), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT2), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n297_), .A3(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT88), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT88), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n301_), .A2(new_n306_), .A3(new_n312_), .A4(new_n309_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n296_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n302_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(new_n307_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n295_), .A2(KEYINPUT1), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n289_), .B1(new_n295_), .B2(KEYINPUT1), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n317_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n283_), .B1(new_n314_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT98), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(KEYINPUT97), .B(new_n209_), .C1(new_n314_), .C2(new_n321_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n296_), .ZN(new_n327_));
  AOI22_X1  g126(.A1(KEYINPUT3), .A2(new_n300_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n312_), .B1(new_n328_), .B2(new_n309_), .ZN(new_n329_));
  AND4_X1   g128(.A1(new_n312_), .A2(new_n301_), .A3(new_n306_), .A4(new_n309_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n327_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT97), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n205_), .A2(new_n332_), .A3(new_n208_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n209_), .A2(KEYINPUT97), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n295_), .A2(KEYINPUT1), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n290_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n316_), .B1(new_n336_), .B2(new_n318_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n331_), .A2(new_n333_), .A3(new_n334_), .A4(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n326_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n325_), .B1(new_n339_), .B2(KEYINPUT4), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n326_), .A2(new_n338_), .B1(G225gat), .B2(G233gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n282_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n323_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n326_), .B2(new_n338_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n343_), .B(new_n281_), .C1(new_n345_), .C2(new_n325_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n274_), .A2(new_n277_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT27), .ZN(new_n350_));
  INV_X1    g149(.A(G197gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G204gat), .ZN(new_n352_));
  INV_X1    g151(.A(G204gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G197gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT91), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G218gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G211gat), .ZN(new_n358_));
  INV_X1    g157(.A(G211gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G218gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n356_), .A2(KEYINPUT21), .A3(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G197gat), .B(G204gat), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(new_n355_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT21), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n365_), .B2(new_n363_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n352_), .A2(new_n354_), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n351_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(KEYINPUT21), .A3(new_n369_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n362_), .A2(new_n364_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n250_), .B2(new_n259_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n373_), .B1(G169gat), .B2(G176gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n237_), .A3(new_n232_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n236_), .A2(new_n229_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n376_), .A2(new_n373_), .B1(new_n246_), .B2(new_n245_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n255_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n256_), .B1(new_n221_), .B2(new_n226_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n234_), .A2(KEYINPUT22), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT22), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G169gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT95), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G169gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(KEYINPUT95), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n235_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n389_), .B(KEYINPUT94), .Z(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n371_), .B(new_n378_), .C1(new_n379_), .C2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT20), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT19), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n372_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n378_), .B1(new_n379_), .B2(new_n392_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n371_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n250_), .A2(new_n371_), .A3(new_n259_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n398_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n397_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n409_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n250_), .A2(new_n371_), .A3(new_n259_), .ZN(new_n412_));
  OAI22_X1  g211(.A1(new_n224_), .A2(new_n225_), .B1(new_n215_), .B2(new_n214_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n224_), .A2(new_n225_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n257_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n383_), .A2(new_n384_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n386_), .A2(KEYINPUT95), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n390_), .B1(new_n418_), .B2(new_n235_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n376_), .A2(new_n373_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n246_), .A2(new_n245_), .ZN(new_n421_));
  AND4_X1   g220(.A1(new_n254_), .A2(new_n420_), .A3(new_n253_), .A4(new_n421_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n415_), .A2(new_n419_), .B1(new_n422_), .B2(new_n375_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT20), .B1(new_n423_), .B2(new_n371_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n396_), .B1(new_n412_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n237_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT79), .B1(new_n236_), .B2(new_n229_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n227_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n414_), .B2(new_n413_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n241_), .A2(new_n247_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT80), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n241_), .A2(new_n242_), .A3(new_n247_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n401_), .B1(new_n433_), .B2(new_n258_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n399_), .B1(new_n423_), .B2(new_n371_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n398_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n411_), .B1(new_n425_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n350_), .B1(new_n410_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT102), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n409_), .B1(new_n397_), .B2(new_n404_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n425_), .A2(new_n411_), .A3(new_n436_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT102), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n350_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G228gat), .A2(G233gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT89), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n371_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT29), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(new_n331_), .B2(new_n337_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n451_), .B2(new_n371_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT29), .B1(new_n314_), .B2(new_n321_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n401_), .A3(new_n448_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G78gat), .B(G106gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT92), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n314_), .A2(new_n321_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G22gat), .B(G50gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT28), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n459_), .A2(new_n450_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n461_), .B1(new_n459_), .B2(new_n450_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n455_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n453_), .A2(new_n401_), .A3(new_n448_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n448_), .B1(new_n453_), .B2(new_n401_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n465_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n458_), .A2(new_n464_), .B1(new_n456_), .B2(new_n468_), .ZN(new_n469_));
  AND4_X1   g268(.A1(KEYINPUT92), .A2(new_n468_), .A3(new_n456_), .A4(new_n464_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT100), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n396_), .B1(new_n372_), .B2(new_n394_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n402_), .A2(new_n398_), .A3(new_n403_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n434_), .A2(new_n435_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT100), .B1(new_n477_), .B2(new_n396_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(KEYINPUT27), .B(new_n441_), .C1(new_n479_), .C2(new_n411_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n445_), .A2(new_n472_), .A3(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n349_), .A2(new_n481_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n469_), .A2(new_n470_), .A3(new_n347_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n443_), .B1(new_n442_), .B2(new_n350_), .ZN(new_n484_));
  AOI211_X1 g283(.A(KEYINPUT102), .B(KEYINPUT27), .C1(new_n440_), .C2(new_n441_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n483_), .B(new_n480_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT103), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT103), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n445_), .A2(new_n488_), .A3(new_n480_), .A4(new_n483_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n339_), .A2(KEYINPUT4), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT99), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n322_), .A2(new_n323_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n490_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT99), .B1(new_n345_), .B2(new_n492_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n281_), .B1(new_n339_), .B2(new_n324_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n440_), .A2(new_n497_), .A3(new_n441_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n346_), .B(KEYINPUT33), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n397_), .A2(new_n404_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n411_), .A2(KEYINPUT32), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n500_), .A2(new_n501_), .B1(new_n342_), .B2(new_n346_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n498_), .A2(new_n499_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT101), .B1(new_n505_), .B2(new_n471_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n504_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n500_), .A2(new_n501_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n347_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n340_), .A2(new_n341_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(KEYINPUT33), .A3(new_n281_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT33), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n346_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n440_), .A2(new_n497_), .A3(new_n441_), .ZN(new_n515_));
  OAI22_X1  g314(.A1(new_n507_), .A2(new_n509_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT101), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n472_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n487_), .A2(new_n489_), .A3(new_n506_), .A4(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n274_), .A2(new_n277_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n482_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G85gat), .A2(G92gat), .ZN(new_n522_));
  INV_X1    g321(.A(G85gat), .ZN(new_n523_));
  INV_X1    g322(.A(G92gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT9), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n522_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n528_));
  OR2_X1    g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT6), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n528_), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT10), .B(G99gat), .Z(new_n533_));
  INV_X1    g332(.A(G106gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n529_), .A2(new_n531_), .A3(new_n532_), .A4(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n525_), .A2(KEYINPUT66), .A3(new_n522_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT65), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n531_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n537_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n543_), .A2(KEYINPUT8), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(KEYINPUT8), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n536_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G29gat), .B(G36gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G43gat), .B(G50gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT15), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n546_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT35), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n543_), .B(KEYINPUT8), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(new_n549_), .A3(new_n536_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n551_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n555_), .A2(new_n556_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n563_));
  INV_X1    g362(.A(new_n561_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n551_), .A2(new_n559_), .A3(new_n564_), .A4(new_n557_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G190gat), .B(G218gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(KEYINPUT36), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n566_), .B(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n562_), .A2(new_n565_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(KEYINPUT36), .A3(new_n569_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G57gat), .B(G64gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT11), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT67), .ZN(new_n578_));
  XOR2_X1   g377(.A(G71gat), .B(G78gat), .Z(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(KEYINPUT11), .B2(new_n576_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n578_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G15gat), .B(G22gat), .ZN(new_n582_));
  INV_X1    g381(.A(G8gat), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G1gat), .B(G8gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n581_), .B(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT72), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT73), .ZN(new_n593_));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT17), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n592_), .A2(new_n593_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n593_), .B1(new_n592_), .B2(new_n599_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT17), .ZN(new_n603_));
  OAI22_X1  g402(.A1(new_n600_), .A2(new_n601_), .B1(new_n603_), .B2(new_n590_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n521_), .A2(new_n575_), .A3(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n578_), .A2(new_n580_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n578_), .A2(new_n580_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n546_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n558_), .A2(new_n581_), .A3(new_n536_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(KEYINPUT12), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT12), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n546_), .A2(new_n612_), .A3(new_n608_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n609_), .A2(new_n610_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT5), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n622_), .B(new_n623_), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n624_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n616_), .A2(new_n619_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT13), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n625_), .A2(KEYINPUT13), .A3(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(G113gat), .B(G141gat), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT74), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G169gat), .B(G197gat), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n634_), .B(new_n635_), .Z(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n550_), .A2(new_n587_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n549_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n587_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n587_), .B(new_n639_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT76), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(KEYINPUT75), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n646_), .B2(KEYINPUT75), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n637_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n650_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n648_), .A3(new_n636_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n632_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n605_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n202_), .B1(new_n656_), .B2(new_n347_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT104), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n575_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n572_), .A2(new_n574_), .A3(new_n659_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n604_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n632_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n521_), .A2(new_n654_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n202_), .A3(new_n347_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT38), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n658_), .A2(new_n671_), .ZN(G1324gat));
  NAND2_X1  g471(.A1(new_n445_), .A2(new_n480_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n583_), .B1(new_n656_), .B2(new_n673_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT105), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(KEYINPUT39), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n656_), .A2(new_n673_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(KEYINPUT39), .A3(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n669_), .A2(new_n583_), .A3(new_n673_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n676_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n676_), .A2(KEYINPUT40), .A3(new_n679_), .A4(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1325gat));
  INV_X1    g484(.A(new_n520_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n267_), .B1(new_n656_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT41), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n669_), .A2(new_n267_), .A3(new_n686_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1326gat));
  INV_X1    g489(.A(G22gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n656_), .B2(new_n471_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT42), .Z(new_n693_));
  NAND3_X1  g492(.A1(new_n669_), .A2(new_n691_), .A3(new_n471_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1327gat));
  NAND2_X1  g494(.A1(new_n604_), .A2(new_n575_), .ZN(new_n696_));
  NOR4_X1   g495(.A1(new_n521_), .A2(new_n696_), .A3(new_n654_), .A4(new_n632_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G29gat), .B1(new_n697_), .B2(new_n347_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n519_), .A2(new_n520_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n482_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n663_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n701_), .A2(KEYINPUT107), .A3(new_n702_), .A4(new_n663_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n663_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n521_), .B2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n705_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n604_), .A2(new_n655_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT106), .ZN(new_n711_));
  AOI211_X1 g510(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n709_), .C2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n521_), .A2(KEYINPUT43), .A3(new_n707_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n708_), .B1(new_n714_), .B2(KEYINPUT107), .ZN(new_n715_));
  INV_X1    g514(.A(new_n706_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n713_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n712_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT44), .B(new_n711_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n347_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n698_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  XNOR2_X1  g523(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n721_), .A2(new_n673_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n726_), .B1(new_n712_), .B2(new_n719_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G36gat), .ZN(new_n728_));
  INV_X1    g527(.A(G36gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n697_), .A2(new_n729_), .A3(new_n673_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT45), .Z(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n725_), .B1(new_n728_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n725_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n731_), .B(new_n734_), .C1(new_n727_), .C2(G36gat), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1329gat));
  AND2_X1   g535(.A1(new_n686_), .A2(G43gat), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n721_), .B(new_n737_), .C1(new_n712_), .C2(new_n719_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G43gat), .B1(new_n697_), .B2(new_n686_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT110), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT47), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n738_), .A2(new_n743_), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1330gat));
  AOI21_X1  g544(.A(G50gat), .B1(new_n697_), .B2(new_n471_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n471_), .A2(G50gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n722_), .B2(new_n747_), .ZN(G1331gat));
  INV_X1    g547(.A(new_n632_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n665_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n654_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n521_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n754_), .A2(KEYINPUT111), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(KEYINPUT111), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n347_), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n749_), .A2(new_n751_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n605_), .A2(KEYINPUT112), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT112), .B1(new_n605_), .B2(new_n759_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n348_), .A2(new_n758_), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n757_), .A2(new_n758_), .B1(new_n762_), .B2(new_n763_), .ZN(G1332gat));
  INV_X1    g563(.A(G64gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n754_), .A2(new_n765_), .A3(new_n673_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n762_), .A2(new_n673_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G64gat), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT48), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT48), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(G1333gat));
  OR3_X1    g570(.A1(new_n753_), .A2(G71gat), .A3(new_n520_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n762_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G71gat), .B1(new_n773_), .B2(new_n520_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(KEYINPUT49), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(G1334gat));
  OR3_X1    g576(.A1(new_n753_), .A2(G78gat), .A3(new_n472_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G78gat), .B1(new_n773_), .B2(new_n472_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT114), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(G78gat), .C1(new_n773_), .C2(new_n472_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n780_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n778_), .B1(new_n784_), .B2(new_n785_), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n715_), .A2(new_n716_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n759_), .A2(new_n604_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n348_), .ZN(new_n791_));
  NOR4_X1   g590(.A1(new_n521_), .A2(new_n696_), .A3(new_n751_), .A4(new_n749_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(new_n523_), .A3(new_n347_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1336gat));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n524_), .A3(new_n673_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n789_), .A2(new_n673_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n797_), .B2(new_n524_), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n790_), .B2(new_n520_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n792_), .A2(new_n533_), .A3(new_n686_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n801_), .B(new_n803_), .ZN(G1338gat));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n709_), .A2(new_n471_), .A3(new_n604_), .A4(new_n759_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n805_), .B1(new_n807_), .B2(new_n534_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n792_), .A2(new_n534_), .A3(new_n471_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT116), .Z(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g612(.A1(new_n520_), .A2(new_n481_), .A3(new_n348_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT120), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n611_), .A2(new_n618_), .A3(new_n613_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n616_), .A2(KEYINPUT55), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n618_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n626_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT56), .B1(new_n817_), .B2(new_n820_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n751_), .B(new_n627_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n638_), .A2(new_n640_), .A3(new_n644_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n643_), .A2(new_n641_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n636_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n646_), .B2(new_n636_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n824_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  INV_X1    g631(.A(new_n575_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(KEYINPUT57), .A4(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n627_), .A2(new_n651_), .A3(new_n653_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n817_), .A2(new_n820_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n835_), .B1(new_n838_), .B2(new_n821_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT57), .B(new_n833_), .C1(new_n839_), .C2(new_n829_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT118), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n834_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n627_), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n843_), .B(new_n828_), .C1(new_n838_), .C2(new_n821_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n844_), .A2(KEYINPUT58), .B1(new_n662_), .B2(new_n661_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n828_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n627_), .B(new_n846_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n845_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n842_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n831_), .A2(new_n833_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(KEYINPUT117), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n575_), .B1(new_n824_), .B2(new_n830_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(KEYINPUT57), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT119), .B1(new_n851_), .B2(new_n858_), .ZN(new_n859_));
  AOI22_X1  g658(.A1(new_n834_), .A2(new_n841_), .B1(new_n845_), .B2(new_n849_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n857_), .A4(new_n854_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n604_), .A3(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n664_), .A2(new_n654_), .A3(new_n749_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT54), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n815_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT59), .ZN(new_n868_));
  INV_X1    g667(.A(new_n815_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n870_));
  INV_X1    g669(.A(new_n865_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n604_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n852_), .A2(new_n853_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n860_), .B2(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n869_), .B(new_n870_), .C1(new_n871_), .C2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n868_), .A2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G113gat), .B1(new_n876_), .B2(new_n654_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n654_), .A2(G113gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n867_), .B2(new_n878_), .ZN(G1340gat));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n632_), .B(new_n875_), .C1(new_n866_), .C2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G120gat), .ZN(new_n882_));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n749_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n866_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n883_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n882_), .A2(new_n885_), .A3(KEYINPUT122), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1341gat));
  INV_X1    g689(.A(new_n876_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n872_), .A2(G127gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(G127gat), .B1(new_n866_), .B2(new_n872_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n893_), .A2(KEYINPUT123), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(KEYINPUT123), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n891_), .A2(new_n892_), .B1(new_n894_), .B2(new_n895_), .ZN(G1342gat));
  OAI21_X1  g695(.A(G134gat), .B1(new_n876_), .B2(new_n707_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n833_), .A2(G134gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n867_), .B2(new_n898_), .ZN(G1343gat));
  NAND2_X1  g698(.A1(new_n863_), .A2(new_n865_), .ZN(new_n900_));
  NOR4_X1   g699(.A1(new_n686_), .A2(new_n673_), .A3(new_n348_), .A4(new_n472_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n654_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n298_), .ZN(G1344gat));
  NOR2_X1   g703(.A1(new_n902_), .A2(new_n749_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n299_), .ZN(G1345gat));
  NOR2_X1   g705(.A1(new_n902_), .A2(new_n604_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT61), .B(G155gat), .Z(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n902_), .B2(new_n707_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n575_), .A2(new_n285_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n902_), .B2(new_n911_), .ZN(G1347gat));
  INV_X1    g711(.A(new_n349_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(new_n472_), .A3(new_n673_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n915_), .B1(new_n871_), .B2(new_n874_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916_), .B2(new_n654_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n919_));
  INV_X1    g718(.A(new_n916_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(new_n751_), .A3(new_n418_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n918_), .B1(new_n919_), .B2(new_n921_), .ZN(G1348gat));
  AOI21_X1  g721(.A(new_n914_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n923_), .A2(G176gat), .A3(new_n632_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n924_), .A2(KEYINPUT124), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n924_), .A2(KEYINPUT124), .ZN(new_n926_));
  AOI21_X1  g725(.A(G176gat), .B1(new_n920_), .B2(new_n632_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(G1349gat));
  AOI21_X1  g727(.A(G183gat), .B1(new_n923_), .B2(new_n872_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n916_), .A2(new_n245_), .A3(new_n604_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n916_), .B2(new_n707_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n575_), .A2(new_n246_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n916_), .B2(new_n933_), .ZN(G1351gat));
  NAND2_X1  g733(.A1(new_n520_), .A2(new_n483_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n673_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n937_), .B1(new_n936_), .B2(new_n935_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n900_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n751_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n632_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g742(.A1(new_n939_), .A2(new_n872_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n359_), .ZN(new_n946_));
  OAI21_X1  g745(.A(KEYINPUT127), .B1(new_n944_), .B2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n939_), .A2(new_n872_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n948_), .A2(new_n949_), .A3(new_n945_), .A4(new_n359_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT63), .B(G211gat), .Z(new_n951_));
  NAND3_X1  g750(.A1(new_n939_), .A2(new_n872_), .A3(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n939_), .A2(KEYINPUT126), .A3(new_n872_), .A4(new_n951_), .ZN(new_n955_));
  AOI22_X1  g754(.A1(new_n947_), .A2(new_n950_), .B1(new_n954_), .B2(new_n955_), .ZN(G1354gat));
  NAND3_X1  g755(.A1(new_n939_), .A2(new_n357_), .A3(new_n575_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n939_), .A2(new_n663_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n958_), .B2(new_n357_), .ZN(G1355gat));
endmodule


