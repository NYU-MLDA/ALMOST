//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n950_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n212_), .A2(new_n213_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n213_), .B1(new_n212_), .B2(new_n218_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT9), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G85gat), .A3(G92gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n209_), .A2(new_n223_), .A3(new_n210_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n216_), .A2(KEYINPUT9), .A3(new_n217_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT10), .B(G99gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n226_), .B2(G106gat), .ZN(new_n227_));
  OAI22_X1  g026(.A1(new_n220_), .A2(new_n221_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G29gat), .B(G36gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G50gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G43gat), .ZN(new_n232_));
  INV_X1    g031(.A(G43gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G50gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n230_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n233_), .A2(G50gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n231_), .A2(G43gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT69), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n229_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G232gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT34), .ZN(new_n246_));
  OAI22_X1  g045(.A1(new_n228_), .A2(new_n244_), .B1(KEYINPUT35), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT66), .B1(new_n227_), .B2(new_n224_), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT10), .B(G99gat), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n205_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n209_), .A2(new_n223_), .A3(new_n210_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .A4(new_n225_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(new_n221_), .B2(new_n220_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT15), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n244_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n238_), .A2(new_n243_), .A3(KEYINPUT15), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n256_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n248_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n246_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT35), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n256_), .A2(new_n260_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT70), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n256_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n267_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n248_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G190gat), .B(G218gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(G134gat), .B(G162gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT36), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT71), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n268_), .A2(new_n274_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n202_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n277_), .B(KEYINPUT36), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n273_), .B1(new_n272_), .B2(new_n248_), .ZN(new_n285_));
  AOI211_X1 g084(.A(new_n267_), .B(new_n247_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n281_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n287_), .B(new_n281_), .C1(new_n282_), .C2(new_n202_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  INV_X1    g092(.A(G1gat), .ZN(new_n294_));
  INV_X1    g093(.A(G8gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT14), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n300_), .B(KEYINPUT73), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n299_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT11), .ZN(new_n303_));
  INV_X1    g102(.A(G78gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G71gat), .ZN(new_n305_));
  INV_X1    g104(.A(G71gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G78gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G57gat), .B(G64gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G57gat), .ZN(new_n312_));
  INV_X1    g111(.A(G64gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G57gat), .A2(G64gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT64), .A3(new_n315_), .ZN(new_n316_));
  AOI211_X1 g115(.A(new_n303_), .B(new_n308_), .C1(new_n311_), .C2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n308_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n311_), .A2(new_n316_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(KEYINPUT11), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n311_), .A2(new_n303_), .A3(new_n316_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n317_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n302_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G127gat), .B(G155gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G211gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT16), .B(G183gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n327_), .A2(KEYINPUT17), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(KEYINPUT17), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n323_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT75), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n323_), .A2(KEYINPUT74), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n323_), .A2(KEYINPUT74), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n328_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n292_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT92), .ZN(new_n338_));
  INV_X1    g137(.A(G141gat), .ZN(new_n339_));
  INV_X1    g138(.A(G148gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT89), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n339_), .B(new_n340_), .C1(new_n341_), .C2(KEYINPUT3), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n343_), .B(KEYINPUT89), .C1(G141gat), .C2(G148gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT90), .B1(G141gat), .B2(G148gat), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n342_), .A2(new_n344_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G141gat), .A2(G148gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT90), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n350_), .A2(KEYINPUT2), .B1(new_n341_), .B2(KEYINPUT3), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G155gat), .ZN(new_n353_));
  INV_X1    g152(.A(G162gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(KEYINPUT88), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT88), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(G155gat), .B2(G162gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n352_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT91), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n355_), .A2(new_n357_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT1), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n358_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n339_), .A2(new_n340_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n348_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n361_), .A2(new_n362_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n359_), .B1(new_n347_), .B2(new_n351_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n368_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT91), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT28), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT28), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n371_), .A2(new_n375_), .A3(new_n378_), .A4(new_n372_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G22gat), .B(G50gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n338_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n377_), .A2(new_n379_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n380_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(KEYINPUT92), .A3(new_n381_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G78gat), .B(G106gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n390_), .B(KEYINPUT94), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G204gat), .ZN(new_n393_));
  AND2_X1   g192(.A1(KEYINPUT93), .A2(G197gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(KEYINPUT93), .A2(G197gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT21), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(G197gat), .B2(G204gat), .ZN(new_n398_));
  OR2_X1    g197(.A1(G211gat), .A2(G218gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G211gat), .A2(G218gat), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n396_), .A2(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(G204gat), .B1(new_n394_), .B2(new_n395_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n393_), .A2(G197gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n397_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n403_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n399_), .A2(KEYINPUT21), .A3(new_n400_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n401_), .A2(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G228gat), .ZN(new_n409_));
  INV_X1    g208(.A(G233gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n371_), .A2(new_n375_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(KEYINPUT29), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT29), .B1(new_n373_), .B2(new_n374_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n412_), .B1(new_n416_), .B2(new_n408_), .ZN(new_n417_));
  OAI211_X1 g216(.A(KEYINPUT95), .B(new_n392_), .C1(new_n415_), .C2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n392_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n417_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n372_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n420_), .B(new_n391_), .C1(new_n421_), .C2(new_n413_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT95), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n419_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n389_), .A2(new_n418_), .A3(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n382_), .A2(new_n383_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT96), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n422_), .A4(new_n419_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n387_), .A2(new_n419_), .A3(new_n381_), .A4(new_n422_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT96), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT87), .B(G113gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G127gat), .ZN(new_n434_));
  INV_X1    g233(.A(G134gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G127gat), .A2(G134gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(G120gat), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(G120gat), .B1(new_n436_), .B2(new_n437_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n433_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(new_n438_), .A3(new_n432_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G71gat), .B(G99gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT85), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n446_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G15gat), .B(G43gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT31), .ZN(new_n451_));
  XOR2_X1   g250(.A(KEYINPUT86), .B(KEYINPUT30), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G183gat), .A2(G190gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n454_), .A2(new_n455_), .A3(KEYINPUT23), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n455_), .B1(new_n454_), .B2(KEYINPUT23), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT23), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(G183gat), .A3(G190gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT83), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(new_n459_), .A3(G183gat), .A4(G190gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n458_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G190gat), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n466_), .A2(KEYINPUT79), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(KEYINPUT79), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT26), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT25), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(KEYINPUT78), .A3(G183gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT26), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(KEYINPUT80), .A3(G190gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(G190gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT80), .ZN(new_n476_));
  NAND2_X1  g275(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n475_), .A2(new_n476_), .B1(KEYINPUT25), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n469_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G169gat), .A2(G176gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT81), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n480_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n465_), .A2(new_n479_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n454_), .A2(KEYINPUT23), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n460_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n467_), .A2(new_n468_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n492_), .B2(G183gat), .ZN(new_n493_));
  INV_X1    g292(.A(G176gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n495_));
  INV_X1    g294(.A(G169gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(KEYINPUT22), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT22), .B(G169gat), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n494_), .B(new_n497_), .C1(new_n498_), .C2(new_n495_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n493_), .A2(new_n485_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n489_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n453_), .B(new_n501_), .Z(new_n502_));
  OR2_X1    g301(.A1(new_n449_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n449_), .A2(new_n502_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n425_), .A2(new_n431_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n444_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n444_), .A2(new_n374_), .A3(new_n373_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT4), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n362_), .B1(new_n361_), .B2(new_n370_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT91), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n444_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G225gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n509_), .A2(new_n510_), .A3(new_n519_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G29gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G85gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT0), .B(G57gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n520_), .A2(new_n522_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n518_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n526_), .B1(new_n529_), .B2(new_n521_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT20), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n501_), .B2(new_n408_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n481_), .A2(KEYINPUT24), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n534_), .A2(KEYINPUT99), .B1(new_n496_), .B2(new_n494_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(KEYINPUT99), .B2(new_n534_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n480_), .B1(new_n490_), .B2(new_n460_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT25), .B(G183gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT98), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n466_), .A2(KEYINPUT26), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n475_), .A2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n536_), .B(new_n537_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n498_), .A2(new_n494_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(G183gat), .A2(G190gat), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT100), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n543_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  AOI211_X1 g346(.A(KEYINPUT100), .B(new_n544_), .C1(new_n458_), .C2(new_n464_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n407_), .B(new_n542_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G226gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n533_), .A2(new_n549_), .A3(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G8gat), .B(G36gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(G92gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT18), .B(G64gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n489_), .A2(new_n407_), .A3(new_n500_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT20), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n542_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n408_), .B2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n554_), .B(new_n559_), .C1(new_n563_), .C2(new_n553_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n564_), .A2(KEYINPUT27), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n533_), .A2(new_n549_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n552_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n408_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n560_), .A2(KEYINPUT20), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n553_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n558_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n565_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n553_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n533_), .A2(new_n549_), .A3(new_n553_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n558_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n564_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n573_), .B1(KEYINPUT27), .B2(new_n578_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n507_), .A2(new_n531_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n531_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT27), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n565_), .A2(new_n572_), .B1(new_n577_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n429_), .B(new_n427_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n424_), .A2(new_n418_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n388_), .B2(new_n384_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n581_), .B(new_n583_), .C1(new_n584_), .C2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n521_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT33), .B1(new_n588_), .B2(new_n527_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n519_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n510_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n514_), .A2(new_n519_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n526_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n576_), .B(new_n564_), .C1(new_n590_), .C2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n589_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n588_), .A2(KEYINPUT33), .A3(new_n527_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n559_), .A2(KEYINPUT32), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n554_), .B(new_n597_), .C1(new_n563_), .C2(new_n553_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n567_), .B2(new_n570_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(KEYINPUT101), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n601_));
  AOI211_X1 g400(.A(new_n601_), .B(new_n597_), .C1(new_n567_), .C2(new_n570_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n595_), .A2(new_n596_), .B1(new_n603_), .B2(new_n531_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n425_), .A2(new_n431_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n587_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n580_), .B1(new_n606_), .B2(new_n505_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n260_), .A2(new_n299_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT77), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G229gat), .A2(G233gat), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n299_), .A2(new_n244_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT77), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n260_), .A2(new_n612_), .A3(new_n299_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .A4(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n299_), .A2(new_n244_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT76), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(KEYINPUT76), .A3(new_n615_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n610_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G169gat), .B(G197gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n614_), .A2(new_n621_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n614_), .B2(new_n621_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT102), .B1(new_n607_), .B2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n256_), .A2(KEYINPUT12), .A3(new_n322_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT12), .ZN(new_n632_));
  INV_X1    g431(.A(new_n316_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT64), .B1(new_n314_), .B2(new_n315_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT11), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n308_), .A3(new_n321_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n319_), .A2(KEYINPUT11), .A3(new_n318_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n227_), .A2(new_n224_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n221_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n640_), .B2(new_n219_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n632_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n631_), .A2(new_n642_), .A3(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n638_), .A2(new_n641_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT65), .B1(new_n322_), .B2(new_n228_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT65), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n638_), .A2(new_n641_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n647_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n646_), .B1(new_n651_), .B2(new_n643_), .ZN(new_n652_));
  XOR2_X1   g451(.A(G176gat), .B(G204gat), .Z(new_n653_));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n652_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n646_), .B(new_n657_), .C1(new_n651_), .C2(new_n643_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n627_), .A2(new_n628_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n603_), .A2(new_n531_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT33), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n528_), .A2(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n590_), .A2(new_n593_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n671_), .A2(new_n578_), .A3(new_n596_), .A4(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n669_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n584_), .A2(new_n586_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n506_), .B1(new_n676_), .B2(new_n587_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n667_), .B(new_n668_), .C1(new_n677_), .C2(new_n580_), .ZN(new_n678_));
  AND4_X1   g477(.A1(new_n337_), .A2(new_n630_), .A3(new_n666_), .A4(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n581_), .A2(G1gat), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT103), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n679_), .A2(new_n683_), .A3(new_n680_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n687_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n682_), .A2(new_n684_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n685_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n629_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n336_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n288_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n696_), .B2(new_n695_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n607_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G1gat), .B1(new_n701_), .B2(new_n581_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n688_), .A2(new_n689_), .A3(new_n692_), .A4(new_n702_), .ZN(G1324gat));
  NAND3_X1  g502(.A1(new_n679_), .A2(new_n295_), .A3(new_n579_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT39), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n700_), .A2(new_n579_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(G8gat), .ZN(new_n707_));
  AOI211_X1 g506(.A(KEYINPUT39), .B(new_n295_), .C1(new_n700_), .C2(new_n579_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n709_), .B(new_n710_), .Z(G1325gat));
  INV_X1    g510(.A(G15gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n700_), .B2(new_n506_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT41), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n679_), .A2(new_n712_), .A3(new_n506_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1326gat));
  INV_X1    g515(.A(G22gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n700_), .B2(new_n605_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT42), .Z(new_n719_));
  NAND3_X1  g518(.A1(new_n679_), .A2(new_n717_), .A3(new_n605_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1327gat));
  NOR2_X1   g520(.A1(new_n694_), .A2(new_n288_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n666_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n630_), .A2(new_n678_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G29gat), .B1(new_n726_), .B2(new_n531_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT110), .B1(KEYINPUT109), .B2(KEYINPUT44), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n607_), .B2(new_n291_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n730_), .B(new_n292_), .C1(new_n677_), .C2(new_n580_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n693_), .A2(new_n733_), .A3(new_n336_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n693_), .B2(new_n336_), .ZN(new_n735_));
  OAI22_X1  g534(.A1(new_n734_), .A2(new_n735_), .B1(KEYINPUT110), .B2(KEYINPUT44), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n728_), .B1(new_n732_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n728_), .ZN(new_n740_));
  AOI211_X1 g539(.A(new_n740_), .B(new_n736_), .C1(new_n729_), .C2(new_n731_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n531_), .A2(G29gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n727_), .B1(new_n743_), .B2(new_n744_), .ZN(G1328gat));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(KEYINPUT112), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(KEYINPUT112), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n583_), .A2(G36gat), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n630_), .A2(new_n678_), .A3(new_n725_), .A4(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT45), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT45), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(G36gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n579_), .B1(new_n738_), .B2(new_n741_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  OAI211_X1 g556(.A(KEYINPUT111), .B(new_n579_), .C1(new_n738_), .C2(new_n741_), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n747_), .B(new_n753_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n747_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n755_), .A2(new_n756_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(G36gat), .A3(new_n758_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n753_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n760_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n759_), .A2(new_n764_), .ZN(G1329gat));
  OAI21_X1  g564(.A(new_n506_), .B1(new_n738_), .B2(new_n741_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G43gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n726_), .A2(new_n233_), .A3(new_n506_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g569(.A1(new_n726_), .A2(new_n231_), .A3(new_n605_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n675_), .B1(new_n739_), .B2(new_n742_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT113), .ZN(new_n773_));
  OAI21_X1  g572(.A(G50gat), .B1(new_n772_), .B2(KEYINPUT113), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n773_), .B2(new_n774_), .ZN(G1331gat));
  NOR3_X1   g574(.A1(new_n607_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(new_n337_), .ZN(new_n777_));
  AOI21_X1  g576(.A(G57gat), .B1(new_n777_), .B2(new_n531_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n776_), .A2(new_n288_), .A3(new_n694_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n581_), .A2(new_n312_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(G1332gat));
  AOI21_X1  g580(.A(new_n313_), .B1(new_n779_), .B2(new_n579_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT48), .Z(new_n783_));
  NAND2_X1  g582(.A1(new_n579_), .A2(new_n313_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT114), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n777_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n786_), .ZN(G1333gat));
  AOI21_X1  g586(.A(new_n306_), .B1(new_n779_), .B2(new_n506_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT49), .Z(new_n789_));
  NAND3_X1  g588(.A1(new_n777_), .A2(new_n306_), .A3(new_n506_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1334gat));
  AOI21_X1  g590(.A(new_n304_), .B1(new_n779_), .B2(new_n605_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT50), .Z(new_n793_));
  NAND2_X1  g592(.A1(new_n605_), .A2(new_n304_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT115), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n777_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n796_), .ZN(G1335gat));
  NAND3_X1  g596(.A1(new_n724_), .A2(new_n336_), .A3(new_n629_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n799_), .A2(new_n531_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n776_), .A2(new_n722_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n531_), .A2(new_n214_), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n800_), .A2(new_n214_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT116), .ZN(G1336gat));
  INV_X1    g603(.A(new_n801_), .ZN(new_n805_));
  AOI21_X1  g604(.A(G92gat), .B1(new_n805_), .B2(new_n579_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n583_), .A2(new_n215_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n799_), .B2(new_n807_), .ZN(G1337gat));
  AND2_X1   g607(.A1(new_n799_), .A2(new_n506_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n506_), .A2(new_n250_), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n809_), .A2(new_n204_), .B1(new_n801_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g611(.A1(new_n805_), .A2(new_n205_), .A3(new_n605_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n799_), .A2(new_n605_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(G106gat), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT52), .B(new_n205_), .C1(new_n799_), .C2(new_n605_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g618(.A1(new_n291_), .A2(new_n694_), .A3(new_n666_), .A4(new_n629_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823_));
  INV_X1    g622(.A(new_n647_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n322_), .A2(new_n228_), .A3(KEYINPUT65), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n649_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n644_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n657_), .B1(new_n828_), .B2(new_n646_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n660_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n609_), .A2(new_n620_), .A3(new_n611_), .A4(new_n613_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n618_), .A2(new_n619_), .A3(new_n610_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n624_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n626_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n823_), .B1(new_n831_), .B2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n661_), .A2(KEYINPUT118), .A3(new_n626_), .A4(new_n834_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n660_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n825_), .A2(new_n826_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n631_), .A2(new_n642_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n644_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n631_), .A2(new_n642_), .A3(new_n645_), .A4(KEYINPUT55), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n646_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n842_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n658_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n846_), .A2(KEYINPUT56), .A3(new_n658_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n839_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT57), .B(new_n288_), .C1(new_n838_), .C2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT120), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n846_), .A2(KEYINPUT56), .A3(new_n658_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT56), .B1(new_n846_), .B2(new_n658_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n837_), .B(new_n836_), .C1(new_n856_), .C2(new_n839_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n857_), .A2(new_n858_), .A3(KEYINPUT57), .A4(new_n288_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n853_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n849_), .A2(new_n850_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n835_), .A2(new_n830_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT58), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n291_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(KEYINPUT58), .A3(new_n862_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n288_), .B1(new_n838_), .B2(new_n851_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n864_), .A2(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n694_), .B1(new_n860_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n822_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  AOI211_X1 g670(.A(KEYINPUT122), .B(new_n694_), .C1(new_n860_), .C2(new_n868_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n507_), .A2(new_n579_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n531_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n877_));
  NAND3_X1  g676(.A1(new_n873_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n864_), .A2(new_n865_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n864_), .A2(KEYINPUT119), .A3(new_n865_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n866_), .A2(new_n867_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n881_), .A2(new_n860_), .A3(new_n882_), .A4(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n336_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n885_), .A2(new_n822_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT59), .B1(new_n886_), .B2(new_n875_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n878_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(G113gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n629_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n886_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n668_), .A3(new_n876_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n888_), .A2(new_n890_), .B1(new_n889_), .B2(new_n892_), .ZN(G1340gat));
  NAND3_X1  g692(.A1(new_n878_), .A2(new_n724_), .A3(new_n887_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G120gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n891_), .A2(new_n876_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G120gat), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n666_), .A2(KEYINPUT60), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(G120gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n895_), .B1(new_n896_), .B2(new_n900_), .ZN(G1341gat));
  NOR2_X1   g700(.A1(new_n336_), .A2(new_n434_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n891_), .A2(new_n694_), .A3(new_n876_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n888_), .A2(new_n902_), .B1(new_n434_), .B2(new_n903_), .ZN(G1342gat));
  XOR2_X1   g703(.A(KEYINPUT123), .B(G134gat), .Z(new_n905_));
  NOR2_X1   g704(.A1(new_n291_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n288_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n891_), .A2(new_n907_), .A3(new_n876_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n888_), .A2(new_n906_), .B1(new_n435_), .B2(new_n908_), .ZN(G1343gat));
  NAND3_X1  g708(.A1(new_n605_), .A2(new_n531_), .A3(new_n505_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n886_), .A2(new_n579_), .A3(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n668_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n724_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g714(.A1(new_n911_), .A2(new_n694_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT61), .B(G155gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1346gat));
  AOI21_X1  g717(.A(G162gat), .B1(new_n911_), .B2(new_n907_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n291_), .A2(new_n354_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n911_), .B2(new_n920_), .ZN(G1347gat));
  NAND3_X1  g720(.A1(new_n579_), .A2(new_n581_), .A3(new_n506_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n605_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n668_), .B(new_n923_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G169gat), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n924_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n873_), .A2(new_n668_), .A3(new_n498_), .A4(new_n923_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n927_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(KEYINPUT124), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n927_), .A2(new_n929_), .A3(new_n932_), .A4(new_n928_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1348gat));
  AND2_X1   g733(.A1(new_n873_), .A2(new_n923_), .ZN(new_n935_));
  AOI21_X1  g734(.A(G176gat), .B1(new_n935_), .B2(new_n724_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n886_), .A2(new_n605_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n922_), .A2(new_n666_), .A3(new_n494_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(G1349gat));
  NOR2_X1   g738(.A1(new_n922_), .A2(new_n336_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G183gat), .B1(new_n937_), .B2(new_n940_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n694_), .A2(new_n539_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n935_), .B2(new_n942_), .ZN(G1350gat));
  NAND4_X1  g742(.A1(new_n935_), .A2(new_n907_), .A3(new_n475_), .A4(new_n540_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n935_), .A2(new_n292_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n944_), .B1(new_n946_), .B2(new_n466_), .ZN(G1351gat));
  NAND4_X1  g746(.A1(new_n605_), .A2(new_n581_), .A3(new_n579_), .A4(new_n505_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n886_), .A2(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(new_n668_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n724_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  NAND2_X1  g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  AND4_X1   g754(.A1(new_n694_), .A2(new_n949_), .A3(new_n954_), .A4(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n954_), .B1(new_n949_), .B2(new_n694_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1354gat));
  XOR2_X1   g757(.A(KEYINPUT125), .B(G218gat), .Z(new_n959_));
  AND3_X1   g758(.A1(new_n949_), .A2(new_n292_), .A3(new_n959_), .ZN(new_n960_));
  NOR3_X1   g759(.A1(new_n886_), .A2(new_n288_), .A3(new_n948_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(new_n959_), .ZN(new_n962_));
  OAI21_X1  g761(.A(KEYINPUT126), .B1(new_n960_), .B2(new_n962_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n949_), .A2(new_n292_), .A3(new_n959_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965_));
  OAI211_X1 g764(.A(new_n964_), .B(new_n965_), .C1(new_n961_), .C2(new_n959_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n963_), .A2(new_n966_), .ZN(G1355gat));
endmodule


