//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT100), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G8gat), .B(G36gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G226gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT19), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT20), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213_));
  XOR2_X1   g012(.A(G211gat), .B(G218gat), .Z(new_n214_));
  INV_X1    g013(.A(KEYINPUT92), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G197gat), .B(G204gat), .Z(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n213_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n217_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n216_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT81), .B(KEYINPUT23), .Z(new_n225_));
  INV_X1    g024(.A(G183gat), .ZN(new_n226_));
  INV_X1    g025(.A(G190gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT82), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n225_), .A2(new_n232_), .A3(new_n229_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G169gat), .ZN(new_n237_));
  INV_X1    g036(.A(G176gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT80), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(G169gat), .B2(G176gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT24), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT25), .B(G183gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT26), .B(G190gat), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n242_), .A2(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT24), .B1(new_n237_), .B2(new_n238_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n236_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n228_), .A2(KEYINPUT23), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n250_), .B1(new_n228_), .B2(new_n225_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n226_), .A2(new_n227_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G169gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n249_), .A2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n212_), .B1(new_n224_), .B2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n242_), .B1(KEYINPUT96), .B2(new_n247_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n247_), .A2(KEYINPUT96), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n230_), .A2(KEYINPUT82), .B1(new_n234_), .B2(new_n228_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n263_), .A2(new_n233_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT97), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n255_), .B(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n262_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT98), .B1(new_n267_), .B2(new_n222_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n266_), .B1(new_n252_), .B2(new_n236_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n261_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT98), .ZN(new_n272_));
  INV_X1    g071(.A(new_n222_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n258_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n210_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n211_), .B1(new_n224_), .B2(new_n257_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n222_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n208_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT101), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n222_), .B(KEYINPUT93), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n249_), .A2(new_n256_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n278_), .B(KEYINPUT20), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n210_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n208_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n274_), .A2(new_n268_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n285_), .B(new_n286_), .C1(new_n287_), .C2(new_n258_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n280_), .A2(new_n281_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT27), .ZN(new_n290_));
  OAI211_X1 g089(.A(KEYINPUT101), .B(new_n208_), .C1(new_n275_), .C2(new_n279_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(KEYINPUT27), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT103), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n295_));
  OAI211_X1 g094(.A(KEYINPUT103), .B(new_n262_), .C1(new_n264_), .C2(new_n266_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n273_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT104), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n298_), .A3(KEYINPUT20), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n282_), .A2(new_n283_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n298_), .B1(new_n297_), .B2(KEYINPUT20), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n210_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n277_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n293_), .B1(new_n305_), .B2(new_n208_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n292_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G78gat), .B(G106gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(G22gat), .B(G50gat), .Z(new_n309_));
  NAND3_X1  g108(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT89), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT3), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT85), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n311_), .B(new_n313_), .C1(KEYINPUT2), .C2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT86), .ZN(new_n318_));
  INV_X1    g117(.A(G155gat), .ZN(new_n319_));
  INV_X1    g118(.A(G162gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT90), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324_));
  OAI22_X1  g123(.A1(new_n318_), .A2(new_n324_), .B1(G155gat), .B2(G162gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n318_), .A2(new_n324_), .ZN(new_n328_));
  OAI221_X1 g127(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .C1(new_n318_), .C2(new_n324_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT88), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n315_), .A2(new_n312_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n323_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n309_), .B1(new_n335_), .B2(KEYINPUT29), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT90), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n322_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n330_), .A2(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT88), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n338_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343_));
  INV_X1    g142(.A(new_n309_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n336_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n336_), .B2(new_n345_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n308_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n336_), .A2(new_n345_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n346_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n308_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n336_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n358_), .B(new_n282_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n273_), .B1(new_n335_), .B2(KEYINPUT29), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n359_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT95), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n361_), .A2(KEYINPUT95), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n359_), .B(new_n362_), .C1(new_n358_), .C2(new_n360_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n350_), .B(new_n356_), .C1(new_n365_), .C2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n307_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G1gat), .B(G29gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G85gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT0), .B(G57gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G127gat), .B(G134gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G113gat), .B(G120gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT84), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n335_), .A2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n378_), .B(new_n323_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n375_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT4), .B1(new_n335_), .B2(new_n379_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n383_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n374_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n379_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n381_), .B1(new_n342_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n384_), .B1(new_n390_), .B2(KEYINPUT4), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n386_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n374_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n387_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n388_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G71gat), .B(G99gat), .ZN(new_n397_));
  INV_X1    g196(.A(G43gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT30), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n283_), .B(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(KEYINPUT83), .B(G15gat), .Z(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n379_), .B(KEYINPUT31), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n406_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n396_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n370_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n383_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n390_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n374_), .B1(new_n413_), .B2(new_n386_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n289_), .A2(new_n291_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT102), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(KEYINPUT33), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n387_), .B1(new_n391_), .B2(new_n386_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n393_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n417_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n374_), .B(new_n420_), .C1(new_n385_), .C2(new_n387_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n415_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n286_), .A2(KEYINPUT32), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n305_), .A2(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n285_), .B(new_n423_), .C1(new_n287_), .C2(new_n258_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n393_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n427_));
  AOI211_X1 g226(.A(new_n374_), .B(new_n387_), .C1(new_n391_), .C2(new_n386_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n425_), .B(new_n426_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n422_), .A2(new_n429_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n364_), .A2(new_n368_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n396_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n292_), .A2(new_n306_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n430_), .A2(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n409_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n411_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G232gat), .A2(G233gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n437_), .B(KEYINPUT34), .Z(new_n438_));
  INV_X1    g237(.A(KEYINPUT35), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G29gat), .B(G36gat), .Z(new_n441_));
  XOR2_X1   g240(.A(G43gat), .B(G50gat), .Z(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT15), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT65), .ZN(new_n446_));
  AND2_X1   g245(.A1(G85gat), .A2(G92gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G85gat), .A2(G92gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G85gat), .ZN(new_n450_));
  INV_X1    g249(.A(G92gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(KEYINPUT65), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT7), .ZN(new_n456_));
  INV_X1    g255(.A(G99gat), .ZN(new_n457_));
  INV_X1    g256(.A(G106gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G99gat), .A2(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT6), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(G99gat), .A3(G106gat), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n461_), .A2(KEYINPUT67), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n459_), .A2(new_n467_), .A3(new_n460_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n455_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT8), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT68), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n460_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT67), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n463_), .A2(new_n465_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n468_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n449_), .A2(new_n454_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT68), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(KEYINPUT8), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT66), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n475_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n470_), .A2(KEYINPUT64), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT64), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT8), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n449_), .A2(new_n454_), .A3(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n481_), .B1(new_n482_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n475_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n477_), .A2(KEYINPUT66), .A3(new_n489_), .A4(new_n486_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n471_), .A2(new_n480_), .A3(new_n488_), .A4(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT10), .B(G99gat), .Z(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n458_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n452_), .A2(KEYINPUT9), .A3(new_n453_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n453_), .A2(KEYINPUT9), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .A4(new_n475_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n445_), .B1(new_n491_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT72), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n440_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n491_), .A2(new_n443_), .A3(new_n496_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n438_), .A2(new_n439_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n496_), .ZN(new_n502_));
  AOI211_X1 g301(.A(KEYINPUT68), .B(new_n470_), .C1(new_n476_), .C2(new_n477_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n488_), .A2(new_n490_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n502_), .B1(new_n505_), .B2(new_n471_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n500_), .B(new_n501_), .C1(new_n506_), .C2(new_n445_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n499_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n497_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n509_), .A2(new_n498_), .A3(new_n440_), .A4(new_n500_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G190gat), .B(G218gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(G134gat), .B(G162gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT73), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT74), .B1(new_n511_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT74), .ZN(new_n519_));
  INV_X1    g318(.A(new_n517_), .ZN(new_n520_));
  AOI211_X1 g319(.A(new_n519_), .B(new_n520_), .C1(new_n508_), .C2(new_n510_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n511_), .A2(KEYINPUT76), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n514_), .B(KEYINPUT36), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT76), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n508_), .A2(new_n526_), .A3(new_n510_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n524_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n436_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G230gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n536_));
  XOR2_X1   g335(.A(G71gat), .B(G78gat), .Z(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n536_), .A2(new_n537_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n480_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n479_), .B1(new_n478_), .B2(KEYINPUT8), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n496_), .B(new_n540_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n491_), .B2(new_n496_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n543_), .B1(new_n544_), .B2(KEYINPUT69), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT69), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n506_), .A2(new_n546_), .A3(new_n540_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n531_), .B(new_n533_), .C1(new_n545_), .C2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G120gat), .B(G148gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G176gat), .B(G204gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n533_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT70), .ZN(new_n555_));
  INV_X1    g354(.A(new_n540_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n542_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n502_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT12), .A3(new_n543_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n560_), .B(new_n556_), .C1(new_n557_), .C2(new_n502_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n533_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n548_), .B(new_n553_), .C1(new_n555_), .C2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n543_), .A2(KEYINPUT12), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(new_n544_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n561_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n532_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(KEYINPUT70), .A3(new_n554_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n553_), .B1(new_n569_), .B2(new_n548_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n564_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n548_), .B1(new_n555_), .B2(new_n562_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n553_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT13), .B1(new_n575_), .B2(new_n563_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n443_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G15gat), .B(G22gat), .ZN(new_n580_));
  INV_X1    g379(.A(G8gat), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G1gat), .B(G8gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT78), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n579_), .A2(new_n585_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n445_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n585_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n590_), .A3(new_n586_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G169gat), .B(G197gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(new_n597_), .Z(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT79), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n592_), .A2(new_n595_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n540_), .B(new_n585_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n609_), .A2(new_n610_), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(KEYINPUT17), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n609_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n578_), .A2(new_n605_), .A3(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n530_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n202_), .B1(new_n621_), .B2(new_n396_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT75), .ZN(new_n623_));
  INV_X1    g422(.A(new_n525_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n511_), .B2(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n508_), .A2(KEYINPUT75), .A3(new_n510_), .A4(new_n525_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT37), .B1(new_n522_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n528_), .B(new_n629_), .C1(new_n518_), .C2(new_n521_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(KEYINPUT77), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT77), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n523_), .A2(new_n632_), .A3(new_n629_), .A4(new_n528_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n577_), .A2(new_n631_), .A3(new_n633_), .A4(new_n618_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n436_), .A2(new_n604_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n436_), .A2(KEYINPUT105), .A3(new_n604_), .A4(new_n635_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n396_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(G1gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT106), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n638_), .A2(new_n644_), .A3(new_n639_), .A4(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n622_), .B1(new_n647_), .B2(KEYINPUT38), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT38), .B1(new_n643_), .B2(new_n645_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n649_), .A2(KEYINPUT107), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(KEYINPUT107), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n650_), .A3(new_n651_), .ZN(G1324gat));
  XNOR2_X1  g451(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n530_), .A2(new_n620_), .A3(new_n307_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G8gat), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(KEYINPUT39), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n654_), .B2(G8gat), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n638_), .A2(new_n639_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n581_), .A3(new_n307_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n653_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n661_), .B(new_n653_), .C1(new_n656_), .C2(new_n658_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n621_), .B2(new_n435_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT41), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n660_), .A2(new_n666_), .A3(new_n435_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n621_), .A2(new_n369_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G22gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT109), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n674_), .A3(G22gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n660_), .A2(new_n679_), .A3(new_n369_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n673_), .A2(KEYINPUT42), .A3(new_n675_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(new_n680_), .A3(new_n681_), .ZN(G1327gat));
  INV_X1    g481(.A(new_n529_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n619_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n578_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n436_), .A2(new_n604_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT111), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n436_), .A2(new_n685_), .A3(new_n688_), .A4(new_n604_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n396_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n577_), .A2(new_n604_), .A3(new_n619_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT110), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n631_), .A2(new_n633_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n430_), .A2(new_n431_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n432_), .A2(new_n433_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n435_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n431_), .A2(new_n433_), .A3(new_n410_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n694_), .B(new_n695_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n694_), .B1(new_n436_), .B2(new_n695_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n693_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(KEYINPUT44), .B(new_n693_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n396_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n691_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  NAND3_X1  g508(.A1(new_n705_), .A2(new_n307_), .A3(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n433_), .A2(G36gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n687_), .A2(new_n689_), .A3(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT45), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n711_), .A2(new_n714_), .A3(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1329gat));
  NAND2_X1  g518(.A1(new_n690_), .A2(new_n435_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n398_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n705_), .A2(G43gat), .A3(new_n435_), .A4(new_n706_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n690_), .B2(new_n369_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n369_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n707_), .B2(new_n726_), .ZN(G1331gat));
  AND4_X1   g526(.A1(new_n603_), .A2(new_n436_), .A3(new_n600_), .A4(new_n578_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n631_), .A2(new_n633_), .A3(new_n618_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G57gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n396_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n577_), .A2(new_n604_), .A3(new_n619_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n530_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n640_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(G1332gat));
  OAI21_X1  g535(.A(G64gat), .B1(new_n734_), .B2(new_n433_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n730_), .A2(new_n740_), .A3(new_n307_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1333gat));
  OAI21_X1  g541(.A(G71gat), .B1(new_n734_), .B2(new_n409_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT49), .ZN(new_n744_));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n730_), .A2(new_n745_), .A3(new_n435_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1334gat));
  INV_X1    g546(.A(G78gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n730_), .A2(new_n748_), .A3(new_n369_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G78gat), .B1(new_n734_), .B2(new_n431_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT50), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT50), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT113), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n749_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1335gat));
  NOR3_X1   g556(.A1(new_n577_), .A2(new_n604_), .A3(new_n618_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n640_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n728_), .A2(new_n683_), .A3(new_n619_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n396_), .A2(new_n450_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(G1336gat));
  OAI21_X1  g562(.A(G92gat), .B1(new_n759_), .B2(new_n433_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n307_), .A2(new_n451_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n761_), .B2(new_n765_), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n759_), .B2(new_n409_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n435_), .A2(new_n492_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n761_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g569(.A(new_n369_), .B(new_n758_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(G106gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G106gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n369_), .A2(new_n458_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n773_), .A2(new_n774_), .B1(new_n761_), .B2(new_n775_), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(G1339gat));
  OAI21_X1  g577(.A(KEYINPUT54), .B1(new_n634_), .B2(new_n604_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n729_), .A2(new_n780_), .A3(new_n605_), .A4(new_n577_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n589_), .A2(new_n590_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n602_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n785_), .A2(KEYINPUT117), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(KEYINPUT117), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n594_), .A2(new_n591_), .A3(new_n586_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n600_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n563_), .B2(new_n575_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n568_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n562_), .A2(KEYINPUT55), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n559_), .A2(new_n533_), .A3(new_n561_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n559_), .A2(KEYINPUT115), .A3(new_n533_), .A4(new_n561_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n793_), .A2(new_n794_), .A3(new_n797_), .A4(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n553_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n553_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AOI211_X1 g603(.A(KEYINPUT116), .B(KEYINPUT56), .C1(new_n799_), .C2(new_n553_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n800_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n604_), .A2(new_n575_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n791_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n783_), .B1(new_n809_), .B2(new_n683_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n802_), .A2(new_n803_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n800_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n797_), .A2(new_n798_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n559_), .A2(new_n561_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT55), .B1(new_n815_), .B2(new_n532_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n792_), .B(new_n533_), .C1(new_n559_), .C2(new_n561_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n574_), .B1(new_n814_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n790_), .A2(new_n570_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n813_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(KEYINPUT58), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n824_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n813_), .A2(new_n820_), .A3(new_n826_), .A4(new_n821_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n695_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT116), .B1(new_n819_), .B2(KEYINPUT56), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n802_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n807_), .B1(new_n831_), .B2(new_n800_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT57), .B(new_n529_), .C1(new_n832_), .C2(new_n791_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n810_), .A2(new_n828_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n782_), .B1(new_n834_), .B2(new_n619_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n370_), .A2(new_n396_), .A3(new_n435_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(G113gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n604_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n619_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n782_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n836_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(KEYINPUT59), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n605_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n839_), .B1(new_n847_), .B2(new_n838_), .ZN(G1340gat));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n577_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n837_), .B(new_n850_), .C1(KEYINPUT60), .C2(new_n849_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n577_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n849_), .ZN(G1341gat));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n619_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT59), .B1(new_n842_), .B2(new_n843_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n835_), .A2(new_n845_), .A3(new_n836_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n837_), .A2(new_n618_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n854_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(new_n860_), .A3(KEYINPUT120), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862_));
  INV_X1    g661(.A(new_n855_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G127gat), .B1(new_n837_), .B2(new_n618_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n862_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n866_), .ZN(G1342gat));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n837_), .A2(new_n868_), .A3(new_n683_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n695_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n871_), .B2(new_n868_), .ZN(G1343gat));
  NOR4_X1   g671(.A1(new_n431_), .A2(new_n307_), .A3(new_n640_), .A4(new_n435_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n842_), .A2(KEYINPUT121), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875_));
  INV_X1    g674(.A(new_n873_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n835_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n605_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT122), .B(G141gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n878_), .B(new_n880_), .ZN(G1344gat));
  AOI21_X1  g680(.A(new_n577_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n882_));
  INV_X1    g681(.A(G148gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1345gat));
  AOI21_X1  g683(.A(new_n619_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n885_), .B(new_n887_), .ZN(G1346gat));
  NAND2_X1  g687(.A1(new_n874_), .A2(new_n877_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n320_), .A3(new_n683_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n870_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n320_), .ZN(G1347gat));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n307_), .A2(new_n410_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT123), .Z(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n369_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n835_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n604_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n893_), .B1(new_n899_), .B2(G169gat), .ZN(new_n900_));
  AOI211_X1 g699(.A(KEYINPUT62), .B(new_n237_), .C1(new_n898_), .C2(new_n604_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n842_), .B2(new_n896_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n835_), .A2(KEYINPUT124), .A3(new_n897_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT22), .B(G169gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n604_), .A2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT125), .ZN(new_n908_));
  OAI22_X1  g707(.A1(new_n900_), .A2(new_n901_), .B1(new_n905_), .B2(new_n908_), .ZN(G1348gat));
  NAND2_X1  g708(.A1(new_n842_), .A2(new_n896_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G176gat), .B1(new_n910_), .B2(new_n577_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n578_), .A2(new_n238_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n905_), .B2(new_n912_), .ZN(G1349gat));
  NOR2_X1   g712(.A1(new_n619_), .A2(new_n244_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n226_), .B1(new_n910_), .B2(new_n619_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n914_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n842_), .A2(new_n902_), .A3(new_n896_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT124), .B1(new_n835_), .B2(new_n897_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(G183gat), .B1(new_n898_), .B2(new_n618_), .ZN(new_n923_));
  OAI21_X1  g722(.A(KEYINPUT126), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n918_), .A2(new_n924_), .ZN(G1350gat));
  AOI21_X1  g724(.A(new_n870_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n683_), .A2(new_n245_), .ZN(new_n927_));
  OAI22_X1  g726(.A1(new_n227_), .A2(new_n926_), .B1(new_n905_), .B2(new_n927_), .ZN(G1351gat));
  AND3_X1   g727(.A1(new_n432_), .A2(new_n307_), .A3(new_n409_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n842_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(G197gat), .B1(new_n931_), .B2(new_n604_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n842_), .A2(G197gat), .A3(new_n604_), .A4(new_n929_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n933_), .A2(KEYINPUT127), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(KEYINPUT127), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n932_), .A2(new_n934_), .A3(new_n935_), .ZN(G1352gat));
  NAND2_X1  g735(.A1(new_n931_), .A2(new_n578_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g737(.A(KEYINPUT63), .B(G211gat), .C1(new_n931_), .C2(new_n618_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT63), .B(G211gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n930_), .A2(new_n619_), .A3(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1354gat));
  OR3_X1    g741(.A1(new_n930_), .A2(G218gat), .A3(new_n529_), .ZN(new_n943_));
  OAI21_X1  g742(.A(G218gat), .B1(new_n930_), .B2(new_n870_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1355gat));
endmodule


