//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G15gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n204_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  OR3_X1    g016(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n218_));
  AND4_X1   g017(.A1(new_n212_), .A2(new_n216_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT80), .B1(new_n214_), .B2(KEYINPUT81), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(KEYINPUT80), .B(KEYINPUT25), .C1(new_n214_), .C2(KEYINPUT81), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n214_), .A2(KEYINPUT80), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n216_), .B(new_n217_), .C1(G183gat), .C2(G190gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(G176gat), .B1(KEYINPUT82), .B2(KEYINPUT22), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G169gat), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n219_), .A2(new_n226_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n207_), .B1(new_n233_), .B2(KEYINPUT84), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT31), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(KEYINPUT84), .ZN(new_n236_));
  INV_X1    g035(.A(G134gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G127gat), .ZN(new_n238_));
  INV_X1    g037(.A(G127gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G134gat), .ZN(new_n240_));
  INV_X1    g039(.A(G120gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G113gat), .ZN(new_n242_));
  INV_X1    g041(.A(G113gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G120gat), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n238_), .A2(new_n240_), .A3(new_n242_), .A4(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT85), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n238_), .A2(new_n240_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n242_), .A2(new_n244_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G113gat), .B(G120gat), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n251_), .A2(KEYINPUT85), .A3(new_n238_), .A4(new_n240_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n247_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n236_), .B(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n235_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n235_), .A2(new_n254_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT94), .ZN(new_n258_));
  XOR2_X1   g057(.A(G211gat), .B(G218gat), .Z(new_n259_));
  INV_X1    g058(.A(KEYINPUT88), .ZN(new_n260_));
  INV_X1    g059(.A(G197gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G204gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT21), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(G197gat), .B2(G204gat), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n259_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT89), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n261_), .B2(G204gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n263_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n262_), .A2(G204gat), .A3(new_n264_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n266_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n268_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n273_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(new_n266_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n276_), .A2(KEYINPUT90), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT90), .B1(new_n276_), .B2(new_n278_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n275_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G141gat), .ZN(new_n282_));
  INV_X1    g081(.A(G148gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(KEYINPUT3), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(G141gat), .B2(G148gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT2), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n288_), .A2(KEYINPUT86), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT86), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n292_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n287_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n282_), .A2(new_n283_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n299_), .A2(new_n289_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n295_), .A2(new_n302_), .A3(new_n296_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT29), .ZN(new_n306_));
  INV_X1    g105(.A(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT87), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(G228gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(G228gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n307_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n281_), .A2(new_n306_), .A3(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n305_), .A2(KEYINPUT29), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT91), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n281_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT90), .ZN(new_n318_));
  AND2_X1   g117(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n321_), .A2(G204gat), .B1(new_n270_), .B2(new_n271_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n259_), .A2(KEYINPUT21), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n318_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n276_), .A2(KEYINPUT90), .A3(new_n278_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(KEYINPUT91), .A3(new_n275_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n315_), .B1(new_n317_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n314_), .B1(new_n328_), .B2(new_n313_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G78gat), .B(G106gat), .ZN(new_n332_));
  OAI211_X1 g131(.A(KEYINPUT92), .B(new_n314_), .C1(new_n328_), .C2(new_n313_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n331_), .A2(KEYINPUT93), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G22gat), .B(G50gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n305_), .A2(KEYINPUT29), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n337_), .A2(new_n338_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n336_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n341_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n339_), .A3(new_n335_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n329_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n332_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n334_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT93), .B1(new_n350_), .B2(new_n333_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n258_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n333_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT93), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n355_), .A2(KEYINPUT94), .A3(new_n334_), .A4(new_n348_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n329_), .B(new_n332_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n345_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n294_), .A2(new_n297_), .B1(new_n303_), .B2(new_n301_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n250_), .A2(new_n245_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT98), .B1(new_n305_), .B2(new_n253_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n247_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT98), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n361_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(KEYINPUT4), .B(new_n363_), .C1(new_n364_), .C2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT99), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n305_), .A2(new_n253_), .A3(KEYINPUT98), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n366_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT99), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(KEYINPUT4), .A4(new_n363_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n305_), .A2(new_n253_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(KEYINPUT4), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n369_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G85gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT0), .B(G57gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n372_), .A2(new_n363_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(new_n380_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n381_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n376_), .B1(new_n368_), .B2(KEYINPUT99), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n379_), .B1(new_n392_), .B2(new_n374_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n385_), .B1(new_n393_), .B2(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT25), .B(G183gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n225_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n211_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT22), .B(G169gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(new_n209_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n219_), .A2(new_n398_), .B1(new_n227_), .B2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n317_), .A2(new_n327_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n219_), .A2(new_n226_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n229_), .A2(new_n227_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n281_), .B2(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G226gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT101), .B1(new_n409_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT20), .B1(new_n281_), .B2(new_n407_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n402_), .B1(new_n326_), .B2(new_n275_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n412_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n412_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT101), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n413_), .A2(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G8gat), .B(G36gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT18), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n414_), .A2(new_n415_), .A3(new_n412_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n324_), .A2(new_n325_), .B1(new_n274_), .B2(new_n268_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n402_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n416_), .B1(new_n408_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n425_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n427_), .A2(KEYINPUT27), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT27), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT20), .B1(new_n429_), .B2(new_n230_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n219_), .A2(new_n398_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n401_), .A2(new_n227_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n281_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n412_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n429_), .A2(new_n230_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n281_), .A2(new_n438_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(KEYINPUT20), .A4(new_n416_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n440_), .A2(new_n443_), .A3(new_n426_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT96), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n440_), .A2(KEYINPUT96), .A3(new_n443_), .A4(new_n426_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n432_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n434_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n433_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n360_), .A2(new_n396_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n425_), .A2(KEYINPUT32), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(new_n421_), .B2(new_n453_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n395_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n389_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT33), .B1(new_n457_), .B2(new_n386_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n459_), .B(new_n385_), .C1(new_n393_), .C2(new_n389_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT97), .B1(new_n446_), .B2(new_n448_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n444_), .A2(new_n445_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT97), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n447_), .A4(new_n432_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n385_), .B1(new_n388_), .B2(new_n380_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n461_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n456_), .B1(new_n469_), .B2(KEYINPUT100), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT100), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n461_), .A2(new_n466_), .A3(new_n471_), .A4(new_n468_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n360_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT102), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n451_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  AOI211_X1 g274(.A(KEYINPUT102), .B(new_n360_), .C1(new_n470_), .C2(new_n472_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n257_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT103), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT103), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n479_), .B(new_n257_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n450_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n360_), .A2(new_n481_), .A3(new_n257_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n396_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT8), .ZN(new_n485_));
  XOR2_X1   g284(.A(G85gat), .B(G92gat), .Z(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT6), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n488_), .B(KEYINPUT67), .Z(new_n489_));
  INV_X1    g288(.A(G99gat), .ZN(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT68), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT7), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n485_), .B(new_n486_), .C1(new_n489_), .C2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n488_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n486_), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n496_), .A2(KEYINPUT69), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT8), .B1(new_n496_), .B2(KEYINPUT69), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT9), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n486_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT66), .B1(new_n502_), .B2(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(KEYINPUT66), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT10), .B(G99gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT65), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n504_), .B(new_n505_), .C1(G106gat), .C2(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n508_), .A2(new_n489_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G57gat), .B(G64gat), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n512_));
  XOR2_X1   g311(.A(G71gat), .B(G78gat), .Z(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n512_), .A2(new_n513_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n499_), .A2(new_n509_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n499_), .B2(new_n509_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT12), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT64), .Z(new_n522_));
  OR2_X1    g321(.A1(new_n519_), .A2(KEYINPUT12), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n499_), .A2(new_n509_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n516_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n517_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n522_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n524_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT70), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n524_), .A2(new_n533_), .A3(new_n530_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G120gat), .B(G148gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT5), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n524_), .A2(new_n530_), .A3(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(KEYINPUT71), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n532_), .A2(new_n543_), .A3(new_n534_), .A4(new_n538_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT72), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT13), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(KEYINPUT13), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(KEYINPUT13), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n542_), .A2(new_n548_), .A3(new_n544_), .A4(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G15gat), .B(G22gat), .Z(new_n552_));
  NAND2_X1  g351(.A1(G1gat), .A2(G8gat), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(KEYINPUT14), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT75), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT76), .ZN(new_n556_));
  XOR2_X1   g355(.A(G1gat), .B(G8gat), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT76), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n555_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n557_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G29gat), .B(G36gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n565_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT78), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n563_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT79), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n568_), .B(KEYINPUT15), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n571_), .B(new_n573_), .C1(new_n563_), .C2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n563_), .B(new_n569_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(new_n572_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G113gat), .B(G141gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G169gat), .B(G197gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n576_), .B(new_n581_), .C1(new_n577_), .C2(new_n572_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n551_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n484_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n516_), .B(new_n589_), .Z(new_n590_));
  OR2_X1    g389(.A1(new_n563_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G127gat), .B(G155gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT16), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n563_), .A2(new_n590_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n591_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT77), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n591_), .A2(new_n598_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n595_), .B(KEYINPUT17), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(KEYINPUT36), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n525_), .A2(new_n574_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT34), .ZN(new_n612_));
  INV_X1    g411(.A(new_n568_), .ZN(new_n613_));
  OAI221_X1 g412(.A(new_n610_), .B1(KEYINPUT35), .B2(new_n612_), .C1(new_n613_), .C2(new_n525_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n616_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT73), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n609_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n617_), .A2(KEYINPUT73), .A3(new_n618_), .A4(new_n608_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(KEYINPUT36), .A3(new_n607_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n625_), .B(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n588_), .A2(new_n604_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(G1gat), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n395_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n625_), .B(KEYINPUT105), .Z(new_n636_));
  NOR3_X1   g435(.A1(new_n588_), .A2(new_n604_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n630_), .B1(new_n637_), .B2(new_n395_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT106), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n631_), .A2(new_n632_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n631_), .A2(new_n632_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(KEYINPUT38), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n639_), .A3(new_n642_), .ZN(G1324gat));
  INV_X1    g442(.A(G8gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n629_), .A2(new_n644_), .A3(new_n481_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n636_), .A2(new_n604_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n484_), .A2(new_n587_), .A3(new_n481_), .A4(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n644_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n648_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n650_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n645_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n645_), .B(new_n656_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1325gat));
  INV_X1    g459(.A(G15gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n257_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n637_), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n629_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1326gat));
  INV_X1    g465(.A(G22gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n629_), .A2(new_n667_), .A3(new_n360_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n637_), .A2(new_n360_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(G22gat), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT42), .B(new_n667_), .C1(new_n637_), .C2(new_n360_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1327gat));
  INV_X1    g474(.A(new_n588_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n625_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n604_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n395_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n551_), .A2(new_n586_), .A3(new_n678_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n625_), .B(new_n626_), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n477_), .A2(KEYINPUT103), .B1(new_n396_), .B2(new_n482_), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT43), .B(new_n684_), .C1(new_n685_), .C2(new_n480_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n484_), .B2(new_n628_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n683_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT44), .B(new_n683_), .C1(new_n686_), .C2(new_n688_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n395_), .A2(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n682_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n691_), .A2(new_n481_), .A3(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n450_), .A2(G36gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n676_), .A2(new_n679_), .A3(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n697_), .A2(KEYINPUT46), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  NAND4_X1  g505(.A1(new_n691_), .A2(G43gat), .A3(new_n662_), .A4(new_n692_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n203_), .B1(new_n680_), .B2(new_n257_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n681_), .B2(new_n360_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n360_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n693_), .B2(new_n713_), .ZN(G1331gat));
  NAND3_X1  g513(.A1(new_n684_), .A2(new_n551_), .A3(new_n678_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT112), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n585_), .B1(new_n685_), .B2(new_n480_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT113), .Z(new_n719_));
  AOI21_X1  g518(.A(G57gat), .B1(new_n719_), .B2(new_n395_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n717_), .A2(new_n551_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n646_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(G57gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n395_), .B2(KEYINPUT114), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(KEYINPUT114), .B2(new_n724_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n720_), .B1(new_n723_), .B2(new_n726_), .ZN(G1332gat));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n719_), .A2(new_n728_), .A3(new_n481_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n723_), .B2(new_n481_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n730_), .A2(new_n731_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n722_), .B2(new_n257_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT49), .ZN(new_n737_));
  INV_X1    g536(.A(G71gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n719_), .A2(new_n738_), .A3(new_n662_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1334gat));
  INV_X1    g539(.A(new_n360_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G78gat), .B1(new_n722_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT50), .ZN(new_n743_));
  INV_X1    g542(.A(G78gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n719_), .A2(new_n744_), .A3(new_n360_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1335gat));
  NAND2_X1  g545(.A1(new_n721_), .A2(new_n679_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(G85gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n395_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n686_), .A2(new_n688_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n551_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n752_), .A2(new_n585_), .A3(new_n678_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n395_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n750_), .B1(new_n757_), .B2(new_n749_), .ZN(G1336gat));
  AOI21_X1  g557(.A(G92gat), .B1(new_n748_), .B2(new_n481_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n481_), .A2(G92gat), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT116), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n759_), .B1(new_n755_), .B2(new_n761_), .ZN(G1337gat));
  OAI21_X1  g561(.A(G99gat), .B1(new_n754_), .B2(new_n257_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n257_), .A2(new_n507_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n747_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT51), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n763_), .B(new_n767_), .C1(new_n747_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1338gat));
  OAI211_X1 g568(.A(new_n360_), .B(new_n753_), .C1(new_n686_), .C2(new_n688_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n491_), .B1(new_n771_), .B2(KEYINPUT52), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(KEYINPUT117), .A3(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n748_), .A2(new_n491_), .A3(new_n360_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n770_), .B(new_n772_), .C1(new_n771_), .C2(KEYINPUT52), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .A4(new_n779_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1339gat));
  NAND2_X1  g582(.A1(new_n482_), .A2(new_n395_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n784_), .A2(KEYINPUT59), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n678_), .A2(new_n586_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT119), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n752_), .A2(new_n787_), .A3(new_n684_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n519_), .A2(KEYINPUT12), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n528_), .B2(KEYINPUT12), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n793_), .B2(new_n522_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n520_), .A2(new_n523_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(KEYINPUT120), .A3(new_n529_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n524_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n793_), .A2(KEYINPUT55), .A3(new_n522_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n794_), .A2(new_n796_), .A3(new_n798_), .A4(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n538_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT56), .B1(new_n800_), .B2(new_n538_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n585_), .B(new_n541_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n573_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n571_), .B(new_n804_), .C1(new_n563_), .C2(new_n575_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n582_), .C1(new_n577_), .C2(new_n804_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n584_), .A2(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n524_), .A2(new_n533_), .A3(new_n530_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n533_), .B1(new_n524_), .B2(new_n530_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n540_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n541_), .A2(KEYINPUT71), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n807_), .B(new_n544_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT121), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n542_), .A2(new_n814_), .A3(new_n544_), .A4(new_n807_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n803_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n677_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n800_), .A2(new_n538_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n538_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n541_), .A3(new_n807_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n824_), .A2(KEYINPUT58), .A3(new_n541_), .A4(new_n807_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n628_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n816_), .A2(KEYINPUT57), .A3(new_n677_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n819_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n831_), .A2(new_n604_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n785_), .B1(new_n790_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n819_), .A2(new_n829_), .A3(KEYINPUT122), .A4(new_n830_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n604_), .A3(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n788_), .B(KEYINPUT54), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n784_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n833_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841_), .B2(new_n586_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n243_), .A3(new_n585_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1340gat));
  OAI211_X1 g643(.A(new_n551_), .B(new_n833_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(G120gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n241_), .B1(new_n752_), .B2(KEYINPUT60), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n839_), .B(new_n847_), .C1(KEYINPUT60), .C2(new_n241_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n846_), .A2(KEYINPUT123), .A3(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1341gat));
  OAI21_X1  g652(.A(G127gat), .B1(new_n841_), .B2(new_n604_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n839_), .A2(new_n239_), .A3(new_n678_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1342gat));
  OAI21_X1  g655(.A(G134gat), .B1(new_n841_), .B2(new_n684_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n839_), .A2(new_n237_), .A3(new_n636_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1343gat));
  NAND2_X1  g658(.A1(new_n837_), .A2(new_n838_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n360_), .ZN(new_n861_));
  NOR4_X1   g660(.A1(new_n861_), .A2(new_n396_), .A3(new_n662_), .A4(new_n481_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n585_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G141gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n282_), .A3(new_n585_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1344gat));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n551_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT124), .B(G148gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n862_), .A2(new_n551_), .A3(new_n868_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1345gat));
  NAND2_X1  g671(.A1(new_n862_), .A2(new_n678_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n874_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n862_), .A2(new_n678_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1346gat));
  INV_X1    g677(.A(G162gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n862_), .A2(new_n879_), .A3(new_n636_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n862_), .A2(new_n628_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n879_), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n790_), .A2(new_n832_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n450_), .A2(new_n395_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n741_), .A2(new_n662_), .A3(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n208_), .B1(new_n886_), .B2(new_n585_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n887_), .A2(KEYINPUT62), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(KEYINPUT62), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n585_), .A3(new_n400_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(G1348gat));
  AOI21_X1  g690(.A(G176gat), .B1(new_n886_), .B2(new_n551_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n360_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n884_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n257_), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n551_), .A2(G176gat), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n892_), .B1(new_n893_), .B2(new_n896_), .ZN(G1349gat));
  NAND3_X1  g696(.A1(new_n893_), .A2(new_n678_), .A3(new_n895_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n604_), .A2(new_n397_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n898_), .A2(new_n214_), .B1(new_n886_), .B2(new_n899_), .ZN(G1350gat));
  AND3_X1   g699(.A1(new_n886_), .A2(new_n225_), .A3(new_n636_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n215_), .B1(new_n886_), .B2(new_n628_), .ZN(new_n902_));
  OR3_X1    g701(.A1(new_n901_), .A2(new_n902_), .A3(KEYINPUT125), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT125), .B1(new_n901_), .B2(new_n902_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1351gat));
  NOR2_X1   g704(.A1(new_n894_), .A2(new_n662_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n860_), .A2(new_n360_), .A3(new_n906_), .ZN(new_n907_));
  OAI22_X1  g706(.A1(new_n907_), .A2(new_n586_), .B1(KEYINPUT126), .B2(new_n261_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n261_), .A2(KEYINPUT126), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n908_), .B(new_n909_), .Z(G1352gat));
  NOR2_X1   g709(.A1(new_n907_), .A2(new_n752_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n263_), .ZN(G1353gat));
  AOI21_X1  g711(.A(new_n604_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n860_), .A2(new_n360_), .A3(new_n906_), .A4(new_n913_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n914_), .A2(KEYINPUT127), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(KEYINPUT127), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n918_));
  INV_X1    g717(.A(G211gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n917_), .A2(new_n920_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n915_), .A2(new_n918_), .A3(new_n919_), .A4(new_n916_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1354gat));
  OAI21_X1  g722(.A(G218gat), .B1(new_n907_), .B2(new_n684_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n636_), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n925_), .A2(G218gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n924_), .B1(new_n907_), .B2(new_n926_), .ZN(G1355gat));
endmodule


