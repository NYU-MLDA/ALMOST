//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n969_, new_n970_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n994_, new_n995_, new_n996_, new_n997_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1005_, new_n1006_,
    new_n1007_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G57gat), .B(G64gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT11), .ZN(new_n208_));
  XOR2_X1   g007(.A(G71gat), .B(G78gat), .Z(new_n209_));
  OR2_X1    g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n209_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n207_), .A2(KEYINPUT11), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT12), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT69), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT10), .B(G99gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT64), .B1(new_n218_), .B2(G106gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n219_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT6), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT9), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(G85gat), .A3(G92gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G85gat), .B(G92gat), .Z(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(KEYINPUT9), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n226_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n236_), .B1(new_n226_), .B2(new_n235_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n217_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n226_), .A2(new_n235_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT65), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n226_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(KEYINPUT69), .A3(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n245_));
  NAND2_X1  g044(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n227_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT7), .ZN(new_n249_));
  INV_X1    g048(.A(G99gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n224_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n245_), .A2(new_n227_), .A3(new_n246_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n248_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n234_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n251_), .A2(new_n229_), .A3(new_n252_), .A4(new_n232_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n234_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n259_), .A2(KEYINPUT8), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n257_), .A2(KEYINPUT8), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n216_), .B1(new_n244_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n241_), .A2(new_n242_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n214_), .B1(new_n263_), .B2(new_n261_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT12), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n260_), .A2(new_n258_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n247_), .A2(new_n253_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n259_), .B1(new_n268_), .B2(new_n255_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT8), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n267_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n271_), .A2(new_n242_), .A3(new_n241_), .A4(new_n213_), .ZN(new_n272_));
  INV_X1    g071(.A(G230gat), .ZN(new_n273_));
  INV_X1    g072(.A(G233gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n262_), .A2(new_n266_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(KEYINPUT67), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n237_), .A2(new_n238_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n271_), .A4(new_n213_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n264_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n273_), .A2(new_n274_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n277_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n206_), .B1(new_n287_), .B2(KEYINPUT70), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n289_), .B(new_n277_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n288_), .A2(KEYINPUT71), .A3(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n277_), .B(new_n206_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT13), .B1(new_n291_), .B2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n261_), .B1(new_n239_), .B2(new_n243_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n213_), .B1(new_n279_), .B2(new_n271_), .ZN(new_n298_));
  OAI22_X1  g097(.A1(new_n297_), .A2(new_n215_), .B1(new_n298_), .B2(KEYINPUT12), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(new_n275_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n282_), .A2(new_n284_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT68), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n300_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT71), .B1(new_n304_), .B2(new_n206_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n205_), .B1(new_n304_), .B2(new_n289_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n290_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n305_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT13), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n288_), .A2(KEYINPUT71), .A3(new_n290_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n296_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT86), .B(G43gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(G15gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(G71gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(new_n250_), .ZN(new_n318_));
  INV_X1    g117(.A(G169gat), .ZN(new_n319_));
  INV_X1    g118(.A(G176gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT22), .B(G169gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n320_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT84), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(KEYINPUT84), .A3(new_n320_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(KEYINPUT85), .A3(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n329_), .A2(new_n332_), .A3(new_n330_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n325_), .A2(new_n326_), .A3(new_n333_), .A4(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT25), .B(G183gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT24), .B1(new_n319_), .B2(new_n320_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n319_), .A2(new_n320_), .A3(KEYINPUT83), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT83), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(G169gat), .B2(G176gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n340_), .B(new_n331_), .C1(new_n346_), .C2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n337_), .A2(KEYINPUT30), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT30), .B1(new_n337_), .B2(new_n349_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n318_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n317_), .B(G99gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n350_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n313_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n353_), .A2(new_n356_), .A3(new_n313_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n360_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT87), .B1(new_n362_), .B2(new_n357_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G127gat), .B(G134gat), .Z(new_n364_));
  XOR2_X1   g163(.A(G113gat), .B(G120gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT31), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n361_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  OAI211_X1 g168(.A(KEYINPUT87), .B(new_n369_), .C1(new_n362_), .C2(new_n357_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT88), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n368_), .A2(KEYINPUT88), .A3(new_n370_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G155gat), .B(G162gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G141gat), .ZN(new_n379_));
  INV_X1    g178(.A(G148gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT3), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(G141gat), .B2(G148gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G141gat), .A2(G148gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT2), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT89), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n378_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n377_), .A2(KEYINPUT1), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n379_), .A2(new_n380_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n385_), .A3(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT90), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n391_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n389_), .B(new_n399_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n381_), .A2(new_n383_), .B1(new_n386_), .B2(new_n385_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n377_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n392_), .A2(new_n395_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT90), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n398_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT28), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n406_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n376_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n410_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n376_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n408_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G22gat), .B(G50gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n398_), .A2(new_n404_), .A3(KEYINPUT29), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n418_), .A2(KEYINPUT91), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G197gat), .B(G204gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT21), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(G197gat), .A2(G204gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G197gat), .A2(G204gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(KEYINPUT21), .A3(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G211gat), .B(G218gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n425_), .A2(new_n426_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n418_), .B2(KEYINPUT91), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n419_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n432_), .B(KEYINPUT92), .Z(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n427_), .A2(new_n428_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n402_), .A2(new_n403_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n435_), .B(new_n436_), .C1(new_n437_), .C2(new_n407_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n417_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n435_), .B1(new_n419_), .B2(new_n430_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n438_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n440_), .A2(new_n441_), .A3(new_n416_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n415_), .B1(new_n439_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n415_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n434_), .A2(new_n438_), .A3(new_n417_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n416_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n366_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n398_), .A2(new_n404_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT96), .B1(new_n437_), .B2(new_n366_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n398_), .A2(new_n404_), .A3(KEYINPUT96), .A4(new_n450_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(KEYINPUT4), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n451_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n449_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n449_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n459_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G1gat), .B(G29gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(G85gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT0), .B(G57gat), .ZN(new_n464_));
  XOR2_X1   g263(.A(new_n463_), .B(new_n464_), .Z(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G8gat), .B(G36gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G64gat), .B(G92gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT19), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n340_), .A2(new_n331_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n342_), .A2(new_n344_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n345_), .B1(new_n478_), .B2(new_n347_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n321_), .B1(new_n322_), .B2(new_n320_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n477_), .A2(new_n479_), .B1(new_n334_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT93), .B1(new_n481_), .B2(new_n429_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n334_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n349_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n485_), .A3(new_n436_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n337_), .A2(new_n429_), .A3(new_n349_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n488_), .A2(KEYINPUT20), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n476_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n337_), .A2(new_n349_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n436_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(new_n484_), .B2(new_n436_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT20), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n475_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n481_), .A2(KEYINPUT94), .A3(new_n429_), .ZN(new_n497_));
  AND4_X1   g296(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .A4(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n473_), .B1(new_n490_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n473_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .A4(new_n497_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n488_), .A2(KEYINPUT20), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(new_n482_), .B2(new_n486_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n500_), .B(new_n501_), .C1(new_n503_), .C2(new_n476_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n465_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n453_), .A2(new_n454_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(new_n449_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n459_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n499_), .B(new_n504_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR4_X1   g309(.A1(new_n458_), .A2(new_n467_), .A3(new_n505_), .A4(new_n460_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n468_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n500_), .A2(KEYINPUT32), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n514_), .B(new_n501_), .C1(new_n503_), .C2(new_n476_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n495_), .B1(new_n481_), .B2(new_n429_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n476_), .B1(new_n492_), .B2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n503_), .B2(new_n476_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n515_), .B1(new_n518_), .B2(new_n514_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n505_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n458_), .A2(new_n505_), .A3(new_n460_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n520_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n448_), .B1(new_n513_), .B2(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n443_), .A2(new_n447_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n499_), .A2(new_n504_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT27), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n504_), .B(KEYINPUT27), .C1(new_n518_), .C2(new_n500_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n529_), .A2(new_n466_), .A3(new_n530_), .A4(new_n521_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n375_), .B1(new_n525_), .B2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n522_), .A2(new_n523_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(new_n371_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n529_), .A2(new_n530_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n448_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G169gat), .B(G197gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G1gat), .A2(G8gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT14), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(G1gat), .A2(G8gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n546_), .A2(new_n547_), .A3(new_n550_), .A4(new_n548_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(G36gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(G29gat), .ZN(new_n556_));
  INV_X1    g355(.A(G29gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(G36gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n558_), .A3(KEYINPUT72), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT72), .B1(new_n556_), .B2(new_n558_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G43gat), .B(G50gat), .Z(new_n562_));
  NOR3_X1   g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G43gat), .B(G50gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n556_), .A2(new_n558_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n564_), .B1(new_n567_), .B2(new_n559_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n554_), .B1(new_n563_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT80), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n562_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(new_n559_), .A3(new_n564_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n571_), .A2(new_n572_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n569_), .A2(new_n570_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n570_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n545_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT81), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n571_), .A2(new_n572_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n578_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n577_), .B(new_n544_), .C1(new_n579_), .C2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n576_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n544_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT81), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n543_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n586_), .A2(new_n576_), .A3(new_n583_), .A4(new_n543_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT82), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT82), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n584_), .A2(new_n590_), .A3(new_n586_), .A4(new_n543_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n587_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n540_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n312_), .B1(new_n594_), .B2(KEYINPUT97), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n580_), .B(new_n578_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n297_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n279_), .A2(new_n271_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n580_), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n604_), .A2(new_n605_), .B1(KEYINPUT35), .B2(new_n597_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n600_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n263_), .A2(new_n261_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n608_), .A2(new_n580_), .B1(new_n599_), .B2(new_n598_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n600_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n609_), .B(new_n610_), .C1(new_n297_), .C2(new_n602_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT76), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT76), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n607_), .A2(new_n611_), .A3(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT74), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT36), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n613_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n619_), .A2(KEYINPUT36), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n607_), .A2(new_n611_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n622_), .A2(new_n623_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n620_), .B1(new_n607_), .B2(new_n611_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT37), .B1(new_n625_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT75), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT75), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n631_), .B(KEYINPUT37), .C1(new_n625_), .C2(new_n628_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n627_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n554_), .B(KEYINPUT77), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G127gat), .B(G155gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n639_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT17), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT79), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(G231gat), .A3(G233gat), .ZN(new_n645_));
  INV_X1    g444(.A(G231gat), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n642_), .B(new_n643_), .C1(new_n646_), .C2(new_n274_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n214_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n214_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n635_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n650_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n634_), .A3(new_n648_), .ZN(new_n653_));
  OR3_X1    g452(.A1(new_n640_), .A2(new_n641_), .A3(KEYINPUT17), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n633_), .A2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT33), .B1(new_n461_), .B2(new_n465_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n658_), .A2(new_n511_), .A3(new_n509_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n519_), .B1(new_n466_), .B2(new_n521_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n526_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n537_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n448_), .A3(new_n534_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  AOI22_X1  g463(.A1(new_n664_), .A2(new_n375_), .B1(new_n538_), .B2(new_n536_), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n665_), .A2(KEYINPUT97), .A3(new_n592_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n595_), .A2(new_n657_), .A3(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT98), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(KEYINPUT98), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n534_), .A2(G1gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n312_), .A2(new_n656_), .A3(new_n592_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n622_), .A2(new_n626_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n665_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT99), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n678_), .A2(KEYINPUT99), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n535_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G1gat), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n671_), .A2(new_n684_), .A3(new_n672_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n673_), .B(new_n683_), .C1(new_n685_), .C2(new_n686_), .ZN(G1324gat));
  NOR2_X1   g486(.A1(new_n662_), .A2(G8gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n668_), .A2(new_n669_), .A3(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n674_), .A2(new_n677_), .A3(new_n537_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G8gat), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(KEYINPUT39), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(KEYINPUT39), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n689_), .B(KEYINPUT40), .C1(new_n693_), .C2(new_n692_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1325gat));
  INV_X1    g497(.A(new_n681_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n679_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n375_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n315_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(KEYINPUT41), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(KEYINPUT41), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n668_), .A2(new_n669_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n701_), .A2(new_n315_), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n703_), .A2(new_n704_), .B1(new_n705_), .B2(new_n706_), .ZN(G1326gat));
  NAND2_X1  g506(.A1(new_n700_), .A2(new_n448_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G22gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G22gat), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n526_), .A2(G22gat), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n710_), .A2(new_n711_), .B1(new_n705_), .B2(new_n712_), .ZN(G1327gat));
  NAND3_X1  g512(.A1(new_n627_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n665_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n540_), .A2(new_n716_), .A3(new_n633_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n296_), .A2(new_n656_), .A3(new_n311_), .A4(new_n593_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n722_), .B(new_n719_), .C1(new_n715_), .C2(new_n717_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n557_), .B1(new_n724_), .B2(new_n535_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n675_), .A2(new_n655_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n595_), .A2(new_n666_), .A3(new_n726_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n727_), .A2(G29gat), .A3(new_n534_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n725_), .A2(new_n728_), .A3(KEYINPUT101), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT101), .B1(new_n725_), .B2(new_n728_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1328gat));
  NOR2_X1   g530(.A1(new_n662_), .A2(G36gat), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n595_), .A2(new_n666_), .A3(new_n726_), .A4(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT45), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n724_), .B2(new_n537_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n716_), .B1(new_n540_), .B2(new_n633_), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT43), .B(new_n714_), .C1(new_n533_), .C2(new_n539_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n720_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n722_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n718_), .A2(KEYINPUT44), .A3(new_n720_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n735_), .A4(new_n537_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G36gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n734_), .B1(new_n736_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT46), .B(new_n734_), .C1(new_n736_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1329gat));
  INV_X1    g547(.A(G43gat), .ZN(new_n749_));
  INV_X1    g548(.A(new_n371_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n724_), .B2(new_n750_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n727_), .A2(G43gat), .A3(new_n375_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753_));
  OR3_X1    g552(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1330gat));
  OR3_X1    g555(.A1(new_n727_), .A2(G50gat), .A3(new_n526_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n724_), .A2(new_n448_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n758_), .A2(KEYINPUT103), .A3(G50gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT103), .B1(new_n758_), .B2(G50gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(G1331gat));
  NAND2_X1  g560(.A1(new_n312_), .A2(new_n592_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(new_n665_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n657_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT104), .ZN(new_n765_));
  INV_X1    g564(.A(G57gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n535_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n656_), .A2(new_n593_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n677_), .A2(new_n312_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n677_), .A2(KEYINPUT105), .A3(new_n312_), .A4(new_n768_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(new_n535_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n767_), .B1(new_n774_), .B2(new_n766_), .ZN(G1332gat));
  NOR2_X1   g574(.A1(new_n662_), .A2(G64gat), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT107), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n765_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n773_), .A2(new_n537_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT106), .B(KEYINPUT48), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(G64gat), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(G64gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(G1333gat));
  NOR2_X1   g582(.A1(new_n375_), .A2(G71gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT109), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n765_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n773_), .A2(new_n701_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n787_), .A2(G71gat), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n787_), .B2(G71gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(G1334gat));
  INV_X1    g590(.A(G78gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n765_), .A2(new_n792_), .A3(new_n448_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n771_), .A2(new_n448_), .A3(new_n772_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(G78gat), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n794_), .B2(G78gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n793_), .B(KEYINPUT111), .C1(new_n796_), .C2(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1335gat));
  AND2_X1   g601(.A1(new_n763_), .A2(new_n726_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G85gat), .B1(new_n803_), .B2(new_n535_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n312_), .A2(new_n656_), .A3(new_n592_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(KEYINPUT112), .Z(new_n807_));
  AND2_X1   g606(.A1(new_n535_), .A2(G85gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(G1336gat));
  AOI21_X1  g608(.A(G92gat), .B1(new_n803_), .B2(new_n537_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n537_), .A2(G92gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n807_), .B2(new_n811_), .ZN(G1337gat));
  INV_X1    g611(.A(new_n806_), .ZN(new_n813_));
  OAI21_X1  g612(.A(G99gat), .B1(new_n813_), .B2(new_n375_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n803_), .A2(new_n222_), .A3(new_n750_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI211_X1 g616(.A(new_n655_), .B(new_n593_), .C1(new_n296_), .C2(new_n311_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n448_), .B(new_n818_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820_));
  OAI21_X1  g619(.A(G106gat), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT113), .B1(new_n806_), .B2(new_n448_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT52), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n819_), .A2(new_n820_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n806_), .A2(KEYINPUT113), .A3(new_n448_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .A4(G106gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n803_), .A2(new_n224_), .A3(new_n448_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT53), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n832_), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1339gat));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n655_), .A2(new_n835_), .A3(new_n592_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n655_), .B2(new_n592_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n296_), .A2(new_n838_), .A3(new_n311_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n296_), .A2(new_n838_), .A3(new_n311_), .A4(KEYINPUT115), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n844_));
  OAI21_X1  g643(.A(new_n714_), .B1(KEYINPUT117), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n844_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n850_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n843_), .A2(new_n852_), .A3(new_n846_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n278_), .A2(new_n281_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n284_), .B1(new_n299_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n299_), .B2(new_n275_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n262_), .A2(KEYINPUT55), .A3(new_n266_), .A4(new_n276_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n856_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n205_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT56), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT56), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n860_), .A2(new_n863_), .A3(new_n205_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n292_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n589_), .A2(new_n591_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n544_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n543_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n545_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n866_), .A2(new_n867_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n867_), .B1(new_n866_), .B2(new_n871_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n854_), .B1(new_n865_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n866_), .A2(new_n871_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT118), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n866_), .A2(new_n867_), .A3(new_n871_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n864_), .A2(new_n292_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(KEYINPUT58), .A4(new_n862_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n875_), .A2(new_n633_), .A3(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n308_), .A2(new_n310_), .A3(new_n879_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n593_), .A3(new_n862_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n676_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n882_), .B1(new_n885_), .B2(KEYINPUT57), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887_));
  AOI211_X1 g686(.A(new_n887_), .B(new_n676_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n656_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n851_), .A2(new_n853_), .A3(new_n889_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n371_), .A2(new_n448_), .A3(new_n537_), .A4(new_n534_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(G113gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(new_n593_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n891_), .A2(new_n895_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n889_), .A2(new_n898_), .ZN(new_n899_));
  OAI211_X1 g698(.A(KEYINPUT119), .B(new_n656_), .C1(new_n886_), .C2(new_n888_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n852_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n850_), .B(new_n845_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n897_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n896_), .A2(new_n905_), .A3(new_n592_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n894_), .B1(new_n906_), .B2(new_n893_), .ZN(G1340gat));
  INV_X1    g706(.A(new_n312_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n896_), .A2(new_n905_), .A3(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(G120gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(KEYINPUT60), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n908_), .A2(KEYINPUT60), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n910_), .ZN(new_n913_));
  AOI21_X1  g712(.A(KEYINPUT120), .B1(new_n892_), .B2(new_n913_), .ZN(new_n914_));
  AND4_X1   g713(.A1(KEYINPUT120), .A2(new_n890_), .A3(new_n891_), .A4(new_n913_), .ZN(new_n915_));
  OAI22_X1  g714(.A1(new_n909_), .A2(new_n910_), .B1(new_n914_), .B2(new_n915_), .ZN(G1341gat));
  INV_X1    g715(.A(G127gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n892_), .A2(new_n917_), .A3(new_n655_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n896_), .A2(new_n905_), .A3(new_n656_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n917_), .ZN(G1342gat));
  AOI21_X1  g719(.A(G134gat), .B1(new_n892_), .B2(new_n676_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n896_), .A2(new_n905_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n633_), .A2(G134gat), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(KEYINPUT121), .Z(new_n924_));
  AOI21_X1  g723(.A(new_n921_), .B1(new_n922_), .B2(new_n924_), .ZN(G1343gat));
  NOR2_X1   g724(.A1(new_n701_), .A2(new_n526_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n890_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n537_), .A2(new_n534_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(new_n593_), .A3(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT122), .B(G141gat), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n927_), .A2(new_n593_), .A3(new_n928_), .A4(new_n930_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1344gat));
  NAND3_X1  g733(.A1(new_n927_), .A2(new_n312_), .A3(new_n928_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(G148gat), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n927_), .A2(new_n380_), .A3(new_n312_), .A4(new_n928_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1345gat));
  NAND3_X1  g737(.A1(new_n927_), .A2(new_n655_), .A3(new_n928_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT61), .B(G155gat), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n940_), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n927_), .A2(new_n655_), .A3(new_n928_), .A4(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1346gat));
  INV_X1    g743(.A(G162gat), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n714_), .A2(new_n945_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(KEYINPUT124), .ZN(new_n947_));
  AND4_X1   g746(.A1(new_n890_), .A2(new_n926_), .A3(new_n928_), .A4(new_n947_), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n890_), .A2(new_n676_), .A3(new_n926_), .A4(new_n928_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(new_n945_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n949_), .A2(KEYINPUT123), .A3(new_n945_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n948_), .B1(new_n952_), .B2(new_n953_), .ZN(G1347gat));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n662_), .A2(new_n535_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n701_), .A2(new_n526_), .A3(new_n956_), .ZN(new_n957_));
  AOI211_X1 g756(.A(new_n592_), .B(new_n957_), .C1(new_n901_), .C2(new_n904_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n955_), .B1(new_n958_), .B2(new_n319_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n957_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n593_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n961_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n958_), .A2(new_n322_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n959_), .A2(new_n962_), .A3(new_n963_), .ZN(G1348gat));
  AOI21_X1  g763(.A(G176gat), .B1(new_n960_), .B2(new_n312_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n957_), .B1(new_n904_), .B2(new_n889_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n908_), .A2(new_n320_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(G1349gat));
  AOI21_X1  g767(.A(G183gat), .B1(new_n966_), .B2(new_n655_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n656_), .A2(new_n338_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n969_), .B1(new_n960_), .B2(new_n970_), .ZN(G1350gat));
  NAND3_X1  g770(.A1(new_n960_), .A2(new_n676_), .A3(new_n339_), .ZN(new_n972_));
  INV_X1    g771(.A(G190gat), .ZN(new_n973_));
  AOI211_X1 g772(.A(KEYINPUT125), .B(new_n973_), .C1(new_n960_), .C2(new_n633_), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n975_));
  INV_X1    g774(.A(new_n957_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n883_), .A2(new_n884_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n977_), .A2(new_n675_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n978_), .A2(new_n887_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n885_), .A2(KEYINPUT57), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n979_), .A2(new_n980_), .A3(new_n882_), .ZN(new_n981_));
  AOI21_X1  g780(.A(KEYINPUT119), .B1(new_n981_), .B2(new_n656_), .ZN(new_n982_));
  INV_X1    g781(.A(new_n900_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(new_n982_), .A2(new_n983_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n851_), .A2(new_n853_), .ZN(new_n985_));
  OAI211_X1 g784(.A(new_n633_), .B(new_n976_), .C1(new_n984_), .C2(new_n985_), .ZN(new_n986_));
  AOI21_X1  g785(.A(new_n975_), .B1(new_n986_), .B2(G190gat), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n972_), .B1(new_n974_), .B2(new_n987_), .ZN(G1351gat));
  NAND4_X1  g787(.A1(new_n890_), .A2(new_n593_), .A3(new_n926_), .A4(new_n956_), .ZN(new_n989_));
  INV_X1    g788(.A(G197gat), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n989_), .B1(KEYINPUT126), .B2(new_n990_), .ZN(new_n991_));
  XOR2_X1   g790(.A(KEYINPUT126), .B(G197gat), .Z(new_n992_));
  AOI21_X1  g791(.A(new_n991_), .B1(new_n989_), .B2(new_n992_), .ZN(G1352gat));
  NAND2_X1  g792(.A1(new_n927_), .A2(new_n956_), .ZN(new_n994_));
  OAI21_X1  g793(.A(G204gat), .B1(new_n994_), .B2(new_n908_), .ZN(new_n995_));
  INV_X1    g794(.A(G204gat), .ZN(new_n996_));
  NAND4_X1  g795(.A1(new_n927_), .A2(new_n996_), .A3(new_n312_), .A4(new_n956_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n995_), .A2(new_n997_), .ZN(G1353gat));
  AOI21_X1  g797(.A(new_n656_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n999_));
  NAND4_X1  g798(.A1(new_n890_), .A2(new_n926_), .A3(new_n956_), .A4(new_n999_), .ZN(new_n1000_));
  NOR2_X1   g799(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1001_));
  AOI21_X1  g800(.A(new_n1000_), .B1(KEYINPUT127), .B2(new_n1001_), .ZN(new_n1002_));
  XNOR2_X1  g801(.A(new_n1001_), .B(KEYINPUT127), .ZN(new_n1003_));
  AOI21_X1  g802(.A(new_n1002_), .B1(new_n1000_), .B2(new_n1003_), .ZN(G1354gat));
  OAI21_X1  g803(.A(G218gat), .B1(new_n994_), .B2(new_n714_), .ZN(new_n1005_));
  NOR2_X1   g804(.A1(new_n675_), .A2(G218gat), .ZN(new_n1006_));
  NAND3_X1  g805(.A1(new_n927_), .A2(new_n956_), .A3(new_n1006_), .ZN(new_n1007_));
  NAND2_X1  g806(.A1(new_n1005_), .A2(new_n1007_), .ZN(G1355gat));
endmodule


