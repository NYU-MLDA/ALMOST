//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n205_), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT9), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(KEYINPUT9), .A3(new_n210_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n204_), .A2(new_n209_), .A3(new_n211_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(new_n203_), .ZN(new_n220_));
  OAI22_X1  g019(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n220_), .B(new_n221_), .C1(new_n206_), .C2(new_n208_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n210_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT66), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n214_), .A2(new_n226_), .A3(new_n210_), .ZN(new_n227_));
  AND4_X1   g026(.A1(new_n217_), .A2(new_n222_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n225_), .A2(new_n227_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n217_), .B1(new_n229_), .B2(new_n222_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n216_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G64gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G57gat), .ZN(new_n233_));
  INV_X1    g032(.A(G57gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G64gat), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n233_), .A2(new_n235_), .A3(KEYINPUT67), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT67), .B1(new_n233_), .B2(new_n235_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT11), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n234_), .A2(G64gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n232_), .A2(G57gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n233_), .A2(new_n235_), .A3(KEYINPUT67), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G71gat), .B(G78gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n238_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(KEYINPUT11), .B(new_n246_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n231_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n222_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT8), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n229_), .A2(new_n217_), .A3(new_n222_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n248_), .A2(new_n249_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n216_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n251_), .A2(KEYINPUT12), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT12), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n231_), .A2(new_n250_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT64), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n251_), .A2(new_n257_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT69), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G120gat), .B(G148gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G176gat), .B(G204gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n272_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n264_), .B(new_n274_), .C1(new_n263_), .C2(new_n265_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n276_), .B(KEYINPUT13), .Z(new_n277_));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n276_), .B(KEYINPUT13), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT70), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G43gat), .B(G50gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G29gat), .B(G36gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n285_), .A2(KEYINPUT71), .ZN(new_n286_));
  INV_X1    g085(.A(G36gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G29gat), .ZN(new_n288_));
  INV_X1    g087(.A(G29gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G36gat), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n288_), .A2(new_n290_), .A3(KEYINPUT71), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n284_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n290_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n285_), .A2(KEYINPUT71), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(new_n283_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT15), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n292_), .A2(KEYINPUT15), .A3(new_n297_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G1gat), .ZN(new_n302_));
  INV_X1    g101(.A(G8gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT14), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT77), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n306_), .B(KEYINPUT14), .C1(new_n302_), .C2(new_n303_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G15gat), .B(G22gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G1gat), .B(G8gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n301_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n292_), .A2(new_n297_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G229gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT83), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n311_), .B(new_n313_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G229gat), .A3(G233gat), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G113gat), .B(G141gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G169gat), .B(G197gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  NOR2_X1   g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n323_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT84), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n320_), .A2(KEYINPUT84), .A3(new_n323_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n324_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n282_), .A2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G8gat), .B(G36gat), .Z(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G64gat), .B(G92gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G204gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G197gat), .ZN(new_n341_));
  INV_X1    g140(.A(G197gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G204gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT21), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT95), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT95), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT21), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n341_), .A2(new_n343_), .A3(new_n345_), .A4(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G211gat), .B(G218gat), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n341_), .A2(new_n343_), .A3(KEYINPUT94), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT21), .B1(new_n341_), .B2(KEYINPUT94), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n348_), .B(new_n349_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n349_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n344_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT89), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT23), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(G183gat), .A3(G190gat), .ZN(new_n362_));
  AOI21_X1  g161(.A(KEYINPUT88), .B1(new_n360_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT88), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n359_), .B2(KEYINPUT23), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n358_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  OAI211_X1 g168(.A(KEYINPUT89), .B(new_n369_), .C1(new_n363_), .C2(new_n365_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT22), .B(G169gat), .ZN(new_n371_));
  INV_X1    g170(.A(G176gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n368_), .A2(new_n370_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n360_), .A2(new_n362_), .ZN(new_n379_));
  INV_X1    g178(.A(G169gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n372_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(KEYINPUT24), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G183gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT25), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G183gat), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT26), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G190gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT26), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n389_), .B(new_n393_), .C1(new_n396_), .C2(new_n392_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n379_), .B(KEYINPUT87), .C1(KEYINPUT24), .C2(new_n381_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n376_), .A2(KEYINPUT24), .A3(new_n381_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n384_), .A2(new_n397_), .A3(new_n398_), .A4(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n357_), .B1(new_n378_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n379_), .A2(new_n369_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n376_), .A3(new_n373_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT99), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(KEYINPUT24), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT24), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(KEYINPUT99), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n381_), .B(new_n374_), .C1(new_n405_), .C2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(KEYINPUT99), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n404_), .A2(KEYINPUT24), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n380_), .A4(new_n372_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n391_), .A2(new_n395_), .A3(new_n386_), .A4(new_n388_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n408_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n403_), .B1(new_n413_), .B2(new_n366_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n356_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n339_), .B1(new_n401_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT20), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n414_), .B2(new_n356_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n378_), .A2(new_n400_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n338_), .B(new_n418_), .C1(new_n419_), .C2(new_n356_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n336_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n418_), .B1(new_n419_), .B2(new_n356_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(new_n338_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT97), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n352_), .A2(new_n425_), .A3(new_n355_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n425_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n414_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT102), .B1(new_n428_), .B2(new_n417_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n401_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT102), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n356_), .A2(KEYINPUT97), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n352_), .A2(new_n425_), .A3(new_n355_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n431_), .B(KEYINPUT20), .C1(new_n434_), .C2(new_n414_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n429_), .A2(new_n430_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n424_), .B1(new_n436_), .B2(new_n338_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n336_), .B(KEYINPUT103), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT27), .B(new_n422_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT98), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G22gat), .B(G50gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT3), .ZN(new_n443_));
  INV_X1    g242(.A(G141gat), .ZN(new_n444_));
  INV_X1    g243(.A(G148gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G141gat), .A2(G148gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT2), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .A4(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G155gat), .ZN(new_n453_));
  INV_X1    g252(.A(G162gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G155gat), .A2(G162gat), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n444_), .A2(new_n445_), .A3(KEYINPUT91), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(G141gat), .B2(G148gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT1), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n455_), .A2(new_n464_), .A3(new_n456_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n466_), .A2(new_n447_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n458_), .A2(new_n459_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT92), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n458_), .A2(new_n468_), .A3(new_n471_), .A4(new_n459_), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n470_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n442_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n470_), .A2(new_n472_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n473_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n470_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n441_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n458_), .A2(new_n468_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT29), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT96), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(new_n487_), .A3(KEYINPUT96), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n487_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n490_), .A2(new_n491_), .B1(new_n492_), .B2(new_n484_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n440_), .B1(new_n482_), .B2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G78gat), .B(G106gat), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n482_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n482_), .B2(new_n493_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n494_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NOR3_X1   g299(.A1(new_n475_), .A2(new_n476_), .A3(new_n442_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n441_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n493_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n495_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n490_), .A2(new_n491_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n483_), .B1(new_n434_), .B2(new_n487_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n481_), .B(new_n477_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n504_), .A2(new_n440_), .A3(new_n507_), .A4(new_n497_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT104), .B(KEYINPUT27), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n416_), .A2(new_n420_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n336_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n512_), .B2(new_n421_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n439_), .A2(new_n500_), .A3(new_n508_), .A4(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G134gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(G127gat), .ZN(new_n516_));
  INV_X1    g315(.A(G127gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G134gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(G120gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G113gat), .ZN(new_n521_));
  INV_X1    g320(.A(G113gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G120gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT90), .B1(new_n519_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n524_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G127gat), .B(G134gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G113gat), .B(G120gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n525_), .B1(new_n530_), .B2(KEYINPUT90), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT4), .B1(new_n531_), .B2(new_n486_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(KEYINPUT90), .ZN(new_n533_));
  INV_X1    g332(.A(new_n525_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n486_), .A3(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n530_), .A2(new_n468_), .A3(new_n458_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n532_), .B1(new_n537_), .B2(KEYINPUT4), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G225gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G1gat), .B(G29gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(G85gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT0), .B(G57gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n540_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n541_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT4), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n551_), .A2(new_n539_), .A3(new_n532_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n545_), .B1(new_n552_), .B2(new_n547_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G227gat), .A2(G233gat), .ZN(new_n556_));
  INV_X1    g355(.A(G15gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT30), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n419_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n531_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G71gat), .B(G99gat), .ZN(new_n563_));
  INV_X1    g362(.A(G43gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT31), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n560_), .A2(new_n561_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n566_), .B1(new_n562_), .B2(new_n567_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n555_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n514_), .A2(new_n571_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n498_), .A2(new_n494_), .A3(new_n499_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n504_), .A2(new_n497_), .B1(new_n440_), .B2(new_n507_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n555_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n439_), .A2(new_n513_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n436_), .A2(new_n338_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n424_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n511_), .A2(KEYINPUT32), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n549_), .A2(new_n553_), .B1(new_n510_), .B2(new_n580_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n538_), .A2(new_n540_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n546_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT101), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(KEYINPUT33), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n547_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n589_), .B1(new_n590_), .B2(new_n546_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n545_), .B(new_n588_), .C1(new_n552_), .C2(new_n547_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n586_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n512_), .A2(new_n421_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n582_), .A2(new_n583_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n500_), .A2(new_n508_), .ZN(new_n596_));
  OAI22_X1  g395(.A1(new_n575_), .A2(new_n576_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n569_), .A2(new_n570_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n572_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n331_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n256_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT78), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n311_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT79), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT79), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT81), .ZN(new_n610_));
  XOR2_X1   g409(.A(G183gat), .B(G211gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n606_), .A2(new_n608_), .A3(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n614_), .B(KEYINPUT17), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n605_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT82), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT82), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n605_), .A2(new_n621_), .A3(new_n618_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n620_), .A3(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT74), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT36), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n255_), .A2(new_n216_), .A3(new_n313_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT34), .Z(new_n631_));
  INV_X1    g430(.A(KEYINPUT35), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT72), .ZN(new_n634_));
  INV_X1    g433(.A(new_n216_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n629_), .B(new_n634_), .C1(new_n301_), .C2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT73), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n638_), .B1(new_n301_), .B2(new_n636_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n631_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n637_), .A2(new_n639_), .A3(KEYINPUT35), .A4(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n633_), .B(KEYINPUT72), .Z(new_n642_));
  AND3_X1   g441(.A1(new_n292_), .A2(KEYINPUT15), .A3(new_n297_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n298_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n644_), .B2(new_n231_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT73), .B1(new_n644_), .B2(new_n231_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n640_), .A2(KEYINPUT35), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n645_), .B(new_n629_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n627_), .A2(KEYINPUT36), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n641_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n641_), .B2(new_n648_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n628_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT76), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT76), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n654_), .B(new_n628_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT37), .B1(new_n650_), .B2(KEYINPUT75), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n657_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n653_), .A2(new_n659_), .A3(new_n655_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n623_), .A2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n600_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(new_n302_), .A3(new_n554_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n279_), .A2(new_n281_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n329_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n623_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n599_), .A2(new_n652_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n302_), .B1(new_n671_), .B2(new_n554_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n666_), .A2(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n673_), .B1(new_n665_), .B2(new_n664_), .ZN(G1324gat));
  NAND3_X1  g473(.A1(new_n663_), .A2(new_n303_), .A3(new_n576_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT39), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n576_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(G8gat), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT39), .B(new_n303_), .C1(new_n671_), .C2(new_n576_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g480(.A(new_n598_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n663_), .A2(new_n557_), .A3(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n671_), .A2(new_n682_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n684_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT41), .B1(new_n684_), .B2(G15gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT105), .ZN(G1326gat));
  INV_X1    g487(.A(G22gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n663_), .A2(new_n689_), .A3(new_n596_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n671_), .A2(new_n596_), .ZN(new_n691_));
  XOR2_X1   g490(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n692_));
  AND3_X1   g491(.A1(new_n691_), .A2(G22gat), .A3(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n691_), .B2(G22gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT107), .ZN(G1327gat));
  INV_X1    g495(.A(new_n652_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n669_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n600_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G29gat), .B1(new_n700_), .B2(new_n554_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n653_), .A2(new_n659_), .A3(new_n655_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n659_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n599_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n439_), .A2(new_n513_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n554_), .B1(new_n500_), .B2(new_n508_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n573_), .A2(new_n574_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n593_), .A2(new_n594_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n583_), .B1(new_n580_), .B2(new_n437_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n682_), .B1(new_n711_), .B2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n661_), .B(new_n708_), .C1(new_n717_), .C2(new_n572_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n702_), .B1(new_n707_), .B2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n661_), .B1(new_n717_), .B2(new_n572_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT109), .B1(new_n720_), .B2(new_n703_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n668_), .B(new_n623_), .C1(new_n719_), .C2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n723_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n555_), .A2(new_n289_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n701_), .B1(new_n726_), .B2(new_n727_), .ZN(G1328gat));
  AND4_X1   g527(.A1(new_n287_), .A2(new_n600_), .A3(new_n576_), .A4(new_n698_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n724_), .A2(new_n576_), .A3(new_n725_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G36gat), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n731_), .A2(new_n733_), .A3(KEYINPUT46), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1329gat));
  NAND4_X1  g537(.A1(new_n724_), .A2(new_n725_), .A3(G43gat), .A4(new_n682_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n564_), .B1(new_n699_), .B2(new_n598_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g541(.A(G50gat), .B1(new_n700_), .B2(new_n596_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n596_), .A2(G50gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n726_), .B2(new_n744_), .ZN(G1331gat));
  NAND4_X1  g544(.A1(new_n617_), .A2(new_n620_), .A3(new_n622_), .A4(new_n329_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n282_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n670_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n748_), .A2(new_n234_), .A3(new_n555_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n282_), .A2(new_n599_), .A3(new_n330_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n662_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT110), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT110), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n554_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n749_), .B1(new_n754_), .B2(new_n234_), .ZN(G1332gat));
  OAI21_X1  g554(.A(G64gat), .B1(new_n748_), .B2(new_n709_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT48), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n751_), .A2(new_n232_), .A3(new_n576_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n748_), .B2(new_n598_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(G71gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n751_), .A2(new_n765_), .A3(new_n682_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1334gat));
  OAI21_X1  g566(.A(G78gat), .B1(new_n748_), .B2(new_n712_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT50), .ZN(new_n769_));
  INV_X1    g568(.A(G78gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n751_), .A2(new_n770_), .A3(new_n596_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1335gat));
  NAND3_X1  g571(.A1(new_n667_), .A2(new_n623_), .A3(new_n329_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n707_), .A2(new_n718_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT109), .ZN(new_n775_));
  INV_X1    g574(.A(new_n721_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n773_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n554_), .A2(G85gat), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT113), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n750_), .A2(new_n698_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n212_), .B1(new_n781_), .B2(new_n555_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT114), .Z(G1336gat));
  AOI21_X1  g583(.A(new_n213_), .B1(new_n777_), .B2(new_n576_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n781_), .A2(G92gat), .A3(new_n709_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT115), .Z(G1337gat));
  INV_X1    g587(.A(new_n781_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(new_n202_), .A3(new_n682_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n777_), .A2(new_n682_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n790_), .B1(new_n792_), .B2(new_n219_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n793_), .B(new_n794_), .Z(G1338gat));
  AND3_X1   g594(.A1(new_n667_), .A2(new_n623_), .A3(new_n329_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n596_), .B(new_n796_), .C1(new_n719_), .C2(new_n721_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(KEYINPUT117), .ZN(new_n798_));
  OAI21_X1  g597(.A(G106gat), .B1(new_n797_), .B2(KEYINPUT117), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n777_), .A2(new_n801_), .A3(new_n596_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(KEYINPUT117), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n802_), .A2(new_n803_), .A3(G106gat), .A4(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n800_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n789_), .A2(new_n203_), .A3(new_n596_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT53), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n810_), .A3(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1339gat));
  NOR3_X1   g611(.A1(new_n514_), .A2(new_n598_), .A3(new_n555_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n316_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n312_), .A2(new_n314_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n323_), .B1(new_n318_), .B2(new_n316_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n327_), .A2(new_n328_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n275_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT121), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT55), .B1(new_n263_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n820_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n261_), .A2(KEYINPUT55), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n821_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n272_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  AOI211_X1 g627(.A(KEYINPUT122), .B(new_n821_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n829_));
  OR3_X1    g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n818_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n661_), .B1(new_n832_), .B2(KEYINPUT58), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n834_), .B(new_n818_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT124), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n831_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT123), .B(new_n828_), .C1(new_n827_), .C2(new_n829_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n830_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n330_), .A2(new_n275_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n841_), .A2(new_n842_), .B1(new_n276_), .B2(new_n817_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n837_), .B1(new_n843_), .B2(new_n652_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n836_), .B1(new_n844_), .B2(KEYINPUT57), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n837_), .B(new_n846_), .C1(new_n843_), .C2(new_n652_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n669_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  AND4_X1   g647(.A1(new_n617_), .A2(new_n620_), .A3(new_n622_), .A4(new_n329_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT118), .B1(new_n849_), .B2(new_n280_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n746_), .A2(new_n277_), .A3(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n706_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT120), .Z(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n706_), .B(new_n855_), .C1(new_n850_), .C2(new_n852_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n813_), .B1(new_n848_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n522_), .A3(new_n330_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n848_), .B2(new_n859_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n860_), .A3(new_n865_), .ZN(new_n866_));
  OAI221_X1 g665(.A(new_n813_), .B1(new_n863_), .B2(KEYINPUT59), .C1(new_n848_), .C2(new_n859_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n329_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n862_), .B1(new_n868_), .B2(new_n522_), .ZN(G1340gat));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT126), .B1(new_n870_), .B2(G120gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(G120gat), .B1(new_n667_), .B2(new_n870_), .ZN(new_n872_));
  MUX2_X1   g671(.A(new_n871_), .B(KEYINPUT126), .S(new_n872_), .Z(new_n873_));
  NAND2_X1  g672(.A1(new_n861_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n282_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n520_), .ZN(G1341gat));
  NAND3_X1  g675(.A1(new_n861_), .A2(new_n517_), .A3(new_n669_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n623_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n517_), .ZN(G1342gat));
  NAND3_X1  g678(.A1(new_n861_), .A2(new_n515_), .A3(new_n652_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n706_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n515_), .ZN(G1343gat));
  OR2_X1    g681(.A1(new_n848_), .A2(new_n859_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n712_), .A2(new_n576_), .A3(new_n555_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n598_), .A3(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(G141gat), .B1(new_n885_), .B2(new_n329_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n848_), .A2(new_n859_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n682_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n888_), .A2(new_n444_), .A3(new_n330_), .A4(new_n884_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(G1344gat));
  OAI21_X1  g689(.A(G148gat), .B1(new_n885_), .B2(new_n282_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n888_), .A2(new_n445_), .A3(new_n667_), .A4(new_n884_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1345gat));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n894_), .B1(new_n885_), .B2(new_n623_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n894_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n888_), .A2(new_n669_), .A3(new_n884_), .A4(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n885_), .B2(new_n706_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n652_), .A2(new_n454_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n885_), .B2(new_n900_), .ZN(G1347gat));
  NOR3_X1   g700(.A1(new_n709_), .A2(new_n571_), .A3(new_n596_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n883_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(new_n371_), .A3(new_n330_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n330_), .B(new_n902_), .C1(new_n848_), .C2(new_n859_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(G169gat), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n904_), .A2(new_n906_), .A3(new_n909_), .ZN(G1348gat));
  NAND3_X1  g709(.A1(new_n883_), .A2(new_n667_), .A3(new_n902_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g711(.A1(new_n883_), .A2(new_n902_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n385_), .B1(new_n913_), .B2(new_n623_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n389_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n883_), .A2(new_n669_), .A3(new_n915_), .A4(new_n902_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n903_), .A2(new_n652_), .A3(new_n396_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G190gat), .B1(new_n913_), .B2(new_n706_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1351gat));
  NOR2_X1   g719(.A1(new_n575_), .A2(new_n709_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n598_), .B(new_n921_), .C1(new_n848_), .C2(new_n859_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n329_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n342_), .ZN(G1352gat));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n282_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n340_), .ZN(G1353gat));
  AOI21_X1  g725(.A(new_n623_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n922_), .A2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT127), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n929_), .B(new_n932_), .ZN(G1354gat));
  OAI21_X1  g732(.A(G218gat), .B1(new_n922_), .B2(new_n706_), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n697_), .A2(G218gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n922_), .B2(new_n935_), .ZN(G1355gat));
endmodule


