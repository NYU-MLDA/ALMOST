//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_;
  XNOR2_X1  g000(.A(KEYINPUT72), .B(G8gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT73), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G1gat), .B(G8gat), .Z(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n208_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G57gat), .B(G64gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n213_));
  XOR2_X1   g012(.A(G71gat), .B(G78gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n213_), .A2(new_n214_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n211_), .B(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G127gat), .B(G155gat), .Z(new_n224_));
  XNOR2_X1  g023(.A(G183gat), .B(G211gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT77), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT17), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n223_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT76), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n222_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT78), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT78), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n239_), .A3(new_n235_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT10), .B(G99gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT64), .B(G106gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G85gat), .B(G92gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n246_), .B1(KEYINPUT9), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G99gat), .A2(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT6), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT6), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(G99gat), .A3(G106gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G85gat), .A2(G92gat), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n249_), .B(new_n254_), .C1(KEYINPUT9), .C2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT8), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G99gat), .A2(G106gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n259_));
  NAND2_X1  g058(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n258_), .A2(new_n260_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n254_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n251_), .A2(new_n253_), .A3(KEYINPUT66), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n263_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n257_), .B1(new_n267_), .B2(new_n248_), .ZN(new_n268_));
  AOI211_X1 g067(.A(KEYINPUT8), .B(new_n247_), .C1(new_n263_), .C2(new_n254_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n256_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n256_), .B(KEYINPUT67), .C1(new_n268_), .C2(new_n269_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n219_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n272_), .A2(KEYINPUT12), .A3(new_n273_), .A4(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n256_), .B(new_n219_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT12), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n270_), .A2(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G230gat), .A2(G233gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n275_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n278_), .A2(new_n276_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n281_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G120gat), .B(G148gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(G176gat), .B(G204gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n283_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n283_), .A2(new_n289_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT13), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n290_), .A2(KEYINPUT13), .A3(new_n291_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G43gat), .B(G50gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n211_), .B(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(G229gat), .A3(G233gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n211_), .A2(new_n299_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n299_), .B(new_n303_), .Z(new_n304_));
  NAND3_X1  g103(.A1(new_n209_), .A2(new_n304_), .A3(new_n210_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G229gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT81), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G113gat), .B(G141gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G169gat), .B(G197gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n301_), .A2(new_n308_), .A3(new_n312_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n243_), .A2(new_n296_), .A3(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT106), .ZN(new_n319_));
  INV_X1    g118(.A(G218gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G211gat), .ZN(new_n321_));
  INV_X1    g120(.A(G211gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G218gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT94), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n321_), .A2(new_n323_), .A3(KEYINPUT94), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(KEYINPUT95), .A3(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G197gat), .B(G204gat), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(KEYINPUT21), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT21), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n321_), .A2(new_n323_), .A3(KEYINPUT94), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT94), .B1(new_n321_), .B2(new_n323_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n335_), .B2(KEYINPUT95), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n326_), .A2(new_n332_), .A3(new_n327_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n329_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n331_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G169gat), .ZN(new_n340_));
  INV_X1    g139(.A(G176gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT22), .B(G169gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n343_), .B2(new_n341_), .ZN(new_n344_));
  INV_X1    g143(.A(G183gat), .ZN(new_n345_));
  INV_X1    g144(.A(G190gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT23), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(G183gat), .A3(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT83), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n352_), .A2(new_n349_), .A3(G183gat), .A4(G190gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n348_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n345_), .A2(new_n346_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n344_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(G183gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n345_), .A2(KEYINPUT25), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n346_), .A2(KEYINPUT26), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT26), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G190gat), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT24), .B1(new_n340_), .B2(new_n341_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n347_), .A2(new_n350_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n366_), .A2(new_n369_), .A3(new_n370_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n357_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n339_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT95), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n333_), .A2(new_n334_), .A3(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n337_), .B(new_n329_), .C1(new_n377_), .C2(new_n332_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n340_), .A2(KEYINPUT22), .ZN(new_n379_));
  AOI21_X1  g178(.A(G176gat), .B1(new_n379_), .B2(KEYINPUT84), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT22), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT85), .B1(new_n381_), .B2(G169gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n383_), .A2(new_n340_), .A3(KEYINPUT22), .ZN(new_n384_));
  OAI221_X1 g183(.A(new_n380_), .B1(KEYINPUT84), .B2(new_n379_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n342_), .B1(new_n370_), .B2(new_n355_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(new_n358_), .B2(G183gat), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n389_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT82), .B1(new_n359_), .B2(new_n360_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n351_), .A2(new_n353_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n347_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n392_), .A2(new_n394_), .A3(new_n369_), .A4(new_n372_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n378_), .A2(new_n331_), .A3(new_n387_), .A4(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n375_), .A2(KEYINPUT20), .A3(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n395_), .A2(new_n387_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n339_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n378_), .A2(new_n331_), .A3(new_n357_), .A4(new_n373_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(KEYINPUT20), .A4(new_n400_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n402_), .A2(new_n407_), .A3(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT20), .B1(new_n339_), .B2(new_n374_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n378_), .A2(new_n331_), .B1(new_n395_), .B2(new_n387_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n401_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n339_), .B2(new_n374_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n400_), .A3(new_n396_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n407_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT102), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT102), .ZN(new_n422_));
  AOI211_X1 g221(.A(new_n422_), .B(new_n407_), .C1(new_n415_), .C2(new_n418_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT27), .B(new_n412_), .C1(new_n421_), .C2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT104), .ZN(new_n425_));
  INV_X1    g224(.A(new_n411_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n400_), .B1(new_n417_), .B2(new_n396_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n420_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n412_), .ZN(new_n429_));
  XOR2_X1   g228(.A(KEYINPUT103), .B(KEYINPUT27), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n425_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  AOI211_X1 g231(.A(KEYINPUT104), .B(new_n430_), .C1(new_n428_), .C2(new_n412_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n424_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n408_), .B(KEYINPUT30), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT87), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G43gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G227gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT86), .B(G15gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n436_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT31), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT31), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n436_), .A2(new_n445_), .A3(new_n442_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n435_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n449_));
  INV_X1    g248(.A(G134gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G127gat), .ZN(new_n451_));
  INV_X1    g250(.A(G127gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G134gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G120gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(G113gat), .ZN(new_n456_));
  INV_X1    g255(.A(G113gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G120gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n451_), .A2(new_n453_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT88), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n454_), .A2(new_n459_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n448_), .A2(new_n449_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n435_), .B2(KEYINPUT87), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n447_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G141gat), .ZN(new_n472_));
  INV_X1    g271(.A(G148gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G141gat), .A2(G148gat), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G155gat), .A2(G162gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT1), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT1), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G155gat), .A3(G162gat), .ZN(new_n480_));
  OR2_X1    g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n476_), .A2(new_n482_), .A3(KEYINPUT89), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n481_), .A2(KEYINPUT92), .A3(new_n477_), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT92), .B1(new_n481_), .B2(new_n477_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n474_), .A2(KEYINPUT3), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n475_), .A2(KEYINPUT2), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT2), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(G141gat), .A3(G148gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n496_));
  NOR4_X1   g295(.A1(new_n496_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(G141gat), .A2(G148gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT3), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT90), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n491_), .B(new_n495_), .C1(new_n497_), .C2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n490_), .B1(new_n501_), .B2(KEYINPUT91), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n496_), .B1(new_n474_), .B2(KEYINPUT3), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n498_), .A2(KEYINPUT90), .A3(new_n499_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n492_), .A2(new_n494_), .B1(new_n474_), .B2(KEYINPUT3), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n487_), .B1(new_n502_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n468_), .ZN(new_n510_));
  OAI221_X1 g309(.A(new_n487_), .B1(new_n461_), .B2(new_n460_), .C1(new_n502_), .C2(new_n508_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT4), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G225gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT100), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n501_), .A2(KEYINPUT91), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n506_), .A2(new_n503_), .A3(new_n507_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n490_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n466_), .B1(new_n518_), .B2(new_n487_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT4), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n515_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n512_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n510_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G1gat), .B(G29gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G85gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT0), .B(G57gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n522_), .A2(new_n523_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n444_), .A2(new_n467_), .A3(new_n446_), .A4(new_n469_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n471_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT29), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n487_), .B(new_n534_), .C1(new_n502_), .C2(new_n508_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT93), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n518_), .A2(KEYINPUT93), .A3(new_n534_), .A4(new_n487_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT28), .B(G22gat), .ZN(new_n539_));
  INV_X1    g338(.A(G50gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n538_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G78gat), .B(G106gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT96), .Z(new_n547_));
  NOR3_X1   g346(.A1(new_n544_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(KEYINPUT97), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n537_), .A2(new_n538_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n541_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n549_), .B1(new_n551_), .B2(new_n543_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n509_), .A2(KEYINPUT29), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n339_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G228gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n548_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n555_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n554_), .B(new_n558_), .ZN(new_n559_));
  OAI22_X1  g358(.A1(new_n544_), .A2(new_n545_), .B1(KEYINPUT97), .B2(new_n547_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n547_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n551_), .A2(new_n561_), .A3(new_n543_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n559_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n557_), .A2(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n434_), .A2(new_n533_), .A3(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n556_), .B1(new_n548_), .B2(new_n552_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n522_), .A2(new_n523_), .A3(new_n528_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT33), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(KEYINPUT101), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n522_), .A2(KEYINPUT33), .A3(new_n523_), .A4(new_n528_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n510_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n510_), .A2(KEYINPUT4), .A3(new_n511_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n513_), .B1(new_n510_), .B2(KEYINPUT4), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n527_), .B(new_n574_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n573_), .A2(new_n428_), .A3(new_n577_), .A4(new_n412_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT101), .B1(new_n569_), .B2(new_n570_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n572_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n522_), .A2(new_n523_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n527_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n569_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n407_), .A2(KEYINPUT32), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n426_), .A2(new_n427_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n568_), .B1(new_n580_), .B2(new_n589_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n426_), .A2(new_n427_), .A3(new_n420_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n407_), .B1(new_n402_), .B2(new_n411_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n431_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT104), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n429_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n566_), .A2(new_n531_), .A3(new_n567_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n424_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n590_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n471_), .A2(new_n532_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n565_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n272_), .A2(new_n304_), .A3(new_n273_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT35), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n256_), .B(new_n299_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n607_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n602_), .A2(new_n609_), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n609_), .B1(new_n602_), .B2(new_n612_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(KEYINPUT36), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n618_), .B(KEYINPUT36), .Z(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT107), .Z(new_n624_));
  NOR2_X1   g423(.A1(new_n601_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n319_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n531_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n237_), .A2(KEYINPUT79), .A3(new_n240_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT79), .B1(new_n237_), .B2(new_n240_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n296_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT37), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n622_), .B2(KEYINPUT71), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n623_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n620_), .B(new_n622_), .C1(KEYINPUT71), .C2(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n630_), .A2(new_n631_), .A3(new_n636_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT80), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n601_), .A2(new_n317_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(KEYINPUT80), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n643_));
  NOR2_X1   g442(.A1(new_n531_), .A2(G1gat), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n643_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n627_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT108), .Z(G1324gat));
  AND3_X1   g447(.A1(new_n642_), .A2(new_n434_), .A3(new_n202_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n434_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G8gat), .B1(new_n626_), .B2(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n654_), .B(new_n656_), .ZN(G1325gat));
  NOR3_X1   g456(.A1(new_n641_), .A2(G15gat), .A3(new_n600_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n659_), .A2(KEYINPUT110), .ZN(new_n660_));
  OAI21_X1  g459(.A(G15gat), .B1(new_n626_), .B2(new_n600_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(KEYINPUT41), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(KEYINPUT41), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(KEYINPUT110), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n660_), .A2(new_n662_), .A3(new_n663_), .A4(new_n664_), .ZN(G1326gat));
  OR3_X1    g464(.A1(new_n641_), .A2(G22gat), .A3(new_n568_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G22gat), .B1(new_n626_), .B2(new_n568_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT42), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT42), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n666_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT111), .ZN(G1327gat));
  INV_X1    g470(.A(new_n623_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n630_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n639_), .A2(new_n672_), .A3(new_n631_), .A4(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT114), .ZN(new_n675_));
  AOI21_X1  g474(.A(G29gat), .B1(new_n675_), .B2(new_n583_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  INV_X1    g476(.A(new_n636_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n600_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n590_), .B2(new_n598_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n677_), .B(new_n678_), .C1(new_n680_), .C2(new_n565_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT112), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n566_), .A2(new_n531_), .A3(new_n567_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n434_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n685_), .B1(new_n529_), .B2(KEYINPUT33), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n428_), .A2(new_n577_), .A3(new_n412_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n571_), .A4(new_n573_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n564_), .B1(new_n688_), .B2(new_n588_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n600_), .B1(new_n684_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n565_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n677_), .A4(new_n678_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n601_), .B2(new_n636_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n682_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n630_), .A2(new_n317_), .A3(new_n296_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT113), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT113), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n698_), .A2(new_n702_), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n696_), .A2(KEYINPUT44), .A3(new_n697_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n705_), .A2(G29gat), .A3(new_n583_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n676_), .B1(new_n704_), .B2(new_n706_), .ZN(G1328gat));
  NOR2_X1   g506(.A1(new_n650_), .A2(G36gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n675_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT45), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n675_), .A2(new_n711_), .A3(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n705_), .ZN(new_n714_));
  AOI211_X1 g513(.A(new_n650_), .B(new_n714_), .C1(new_n701_), .C2(new_n703_), .ZN(new_n715_));
  INV_X1    g514(.A(G36gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n713_), .B(KEYINPUT46), .C1(new_n715_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  NAND2_X1  g520(.A1(new_n675_), .A2(new_n679_), .ZN(new_n722_));
  INV_X1    g521(.A(G43gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n600_), .A2(new_n723_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n705_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT115), .B1(new_n704_), .B2(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n702_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT113), .B(KEYINPUT44), .C1(new_n696_), .C2(new_n697_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n726_), .B(KEYINPUT115), .C1(new_n728_), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n724_), .B1(new_n727_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT47), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n734_), .B(new_n724_), .C1(new_n727_), .C2(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1330gat));
  AOI21_X1  g535(.A(G50gat), .B1(new_n675_), .B2(new_n564_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n714_), .A2(new_n540_), .A3(new_n568_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n704_), .B2(new_n738_), .ZN(G1331gat));
  NAND4_X1  g538(.A1(new_n625_), .A2(new_n317_), .A3(new_n296_), .A4(new_n630_), .ZN(new_n740_));
  INV_X1    g539(.A(G57gat), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n531_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n630_), .A2(new_n296_), .A3(new_n636_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT116), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n601_), .A2(new_n316_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n747_), .A2(KEYINPUT117), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(KEYINPUT117), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n583_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n741_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT118), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(KEYINPUT118), .A3(new_n741_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n742_), .B1(new_n753_), .B2(new_n754_), .ZN(G1332gat));
  AND2_X1   g554(.A1(new_n748_), .A2(new_n749_), .ZN(new_n756_));
  INV_X1    g555(.A(G64gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n434_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G64gat), .B1(new_n740_), .B2(new_n650_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT48), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1333gat));
  INV_X1    g560(.A(G71gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n756_), .A2(new_n762_), .A3(new_n679_), .ZN(new_n763_));
  OAI21_X1  g562(.A(G71gat), .B1(new_n740_), .B2(new_n600_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT49), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1334gat));
  INV_X1    g565(.A(G78gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n756_), .A2(new_n767_), .A3(new_n564_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G78gat), .B1(new_n740_), .B2(new_n568_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT50), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1335gat));
  NOR3_X1   g570(.A1(new_n630_), .A2(new_n631_), .A3(new_n316_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT120), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n696_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT121), .ZN(new_n775_));
  INV_X1    g574(.A(G85gat), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n531_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n745_), .A2(new_n672_), .A3(new_n296_), .A4(new_n673_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n778_), .B2(new_n531_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT119), .Z(new_n780_));
  NOR2_X1   g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1336gat));
  OAI21_X1  g580(.A(G92gat), .B1(new_n775_), .B2(new_n650_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n650_), .A2(G92gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n778_), .B2(new_n783_), .ZN(G1337gat));
  OAI21_X1  g583(.A(G99gat), .B1(new_n774_), .B2(new_n600_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n600_), .A2(new_n244_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n778_), .B2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g587(.A1(new_n778_), .A2(new_n568_), .A3(new_n245_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n773_), .A2(new_n564_), .A3(new_n696_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(G106gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(G106gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g594(.A1(new_n630_), .A2(new_n631_), .A3(new_n317_), .A4(new_n636_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT54), .Z(new_n797_));
  NAND2_X1  g596(.A1(new_n316_), .A2(new_n290_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n275_), .A2(new_n279_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT122), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT122), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n275_), .A2(new_n279_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n280_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT123), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT123), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n800_), .A2(new_n806_), .A3(new_n803_), .A4(new_n802_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n281_), .B(KEYINPUT55), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n289_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(KEYINPUT56), .A3(new_n289_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n798_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n300_), .A2(new_n307_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n307_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n302_), .A2(new_n305_), .A3(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n313_), .A3(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n292_), .A2(new_n315_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n623_), .B1(new_n814_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT57), .B(new_n623_), .C1(new_n814_), .C2(new_n820_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n290_), .A2(new_n315_), .A3(new_n818_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n289_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n813_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n809_), .A2(KEYINPUT124), .A3(KEYINPUT56), .A4(new_n289_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n825_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n678_), .B1(new_n830_), .B2(KEYINPUT58), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n813_), .A2(new_n827_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n829_), .A3(new_n812_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n825_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n823_), .B(new_n824_), .C1(new_n831_), .C2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n797_), .B1(new_n836_), .B2(new_n243_), .ZN(new_n837_));
  NOR4_X1   g636(.A1(new_n434_), .A2(new_n600_), .A3(new_n564_), .A4(new_n531_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n457_), .A3(new_n316_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT59), .B1(new_n837_), .B2(new_n839_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT58), .B1(new_n833_), .B2(new_n834_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n835_), .A2(new_n843_), .A3(new_n636_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n823_), .A2(new_n824_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n673_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n797_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n839_), .A2(KEYINPUT59), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n842_), .A2(new_n316_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n841_), .B1(new_n852_), .B2(new_n457_), .ZN(G1340gat));
  AOI21_X1  g652(.A(new_n631_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n455_), .B1(new_n854_), .B2(new_n842_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT60), .ZN(new_n856_));
  AOI21_X1  g655(.A(G120gat), .B1(new_n296_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n856_), .B2(G120gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n840_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT125), .B1(new_n855_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n243_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n847_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n864_), .B2(new_n838_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n797_), .B1(new_n836_), .B2(new_n673_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n849_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n296_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G120gat), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n859_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n861_), .A2(new_n871_), .ZN(G1341gat));
  NAND3_X1  g671(.A1(new_n840_), .A2(new_n452_), .A3(new_n630_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n842_), .A2(new_n242_), .A3(new_n850_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n875_), .B2(new_n452_), .ZN(G1342gat));
  NAND3_X1  g675(.A1(new_n840_), .A2(new_n450_), .A3(new_n624_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n842_), .A2(new_n678_), .A3(new_n850_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n877_), .B1(new_n879_), .B2(new_n450_), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n679_), .A2(new_n568_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n650_), .A2(new_n583_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n823_), .A2(new_n824_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n843_), .A2(new_n636_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n835_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n242_), .B1(new_n884_), .B2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n881_), .B(new_n883_), .C1(new_n888_), .C2(new_n797_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n317_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n472_), .ZN(G1344gat));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n631_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n473_), .ZN(G1345gat));
  OAI21_X1  g692(.A(KEYINPUT126), .B1(new_n889_), .B2(new_n673_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n881_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n863_), .B2(new_n847_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(new_n630_), .A4(new_n883_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n898_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n894_), .A2(new_n898_), .A3(new_n900_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n889_), .B2(new_n636_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n624_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n906_), .A2(G162gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n889_), .B2(new_n907_), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n650_), .A2(new_n533_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n848_), .A2(new_n568_), .A3(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n317_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n909_), .B1(new_n912_), .B2(new_n340_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n343_), .ZN(new_n914_));
  OAI211_X1 g713(.A(KEYINPUT62), .B(G169gat), .C1(new_n911_), .C2(new_n317_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(G1348gat));
  INV_X1    g715(.A(new_n911_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G176gat), .B1(new_n917_), .B2(new_n296_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n837_), .A2(new_n564_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n296_), .A2(new_n910_), .A3(G176gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1349gat));
  NOR3_X1   g720(.A1(new_n911_), .A2(new_n361_), .A3(new_n243_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n919_), .A2(new_n630_), .A3(new_n910_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n345_), .B2(new_n923_), .ZN(G1350gat));
  OAI21_X1  g723(.A(G190gat), .B1(new_n911_), .B2(new_n636_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n624_), .A2(new_n365_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n911_), .B2(new_n926_), .ZN(G1351gat));
  NAND3_X1  g726(.A1(new_n896_), .A2(new_n531_), .A3(new_n434_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n317_), .ZN(new_n929_));
  INV_X1    g728(.A(G197gat), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1352gat));
  NOR2_X1   g730(.A1(new_n928_), .A2(new_n631_), .ZN(new_n932_));
  INV_X1    g731(.A(G204gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1353gat));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n242_), .B1(new_n935_), .B2(new_n322_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n928_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(KEYINPUT127), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n937_), .B(new_n939_), .ZN(G1354gat));
  OAI21_X1  g739(.A(G218gat), .B1(new_n928_), .B2(new_n636_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n624_), .A2(new_n320_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n928_), .B2(new_n942_), .ZN(G1355gat));
endmodule


