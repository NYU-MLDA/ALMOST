//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT18), .B(G64gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G8gat), .B(G36gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207_));
  INV_X1    g006(.A(G204gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G197gat), .ZN(new_n209_));
  INV_X1    g008(.A(G197gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G204gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n207_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(G211gat), .A2(G218gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G211gat), .A2(G218gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT88), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n212_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT89), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G197gat), .B(G204gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n217_), .B1(new_n218_), .B2(new_n207_), .ZN(new_n219_));
  AND4_X1   g018(.A1(new_n217_), .A2(new_n209_), .A3(new_n211_), .A4(new_n207_), .ZN(new_n220_));
  OAI22_X1  g019(.A1(new_n219_), .A2(new_n220_), .B1(new_n214_), .B2(new_n213_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AND3_X1   g022(.A1(KEYINPUT77), .A2(G183gat), .A3(G190gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT77), .B1(G183gat), .B2(G190gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT23), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  OR3_X1    g026(.A1(new_n227_), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT78), .B1(new_n227_), .B2(KEYINPUT23), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n226_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n231_));
  INV_X1    g030(.A(G169gat), .ZN(new_n232_));
  INV_X1    g031(.A(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n235_), .A3(KEYINPUT97), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT97), .B1(new_n230_), .B2(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n231_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT25), .B(G183gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT26), .B(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n237_), .A2(new_n238_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT22), .B(G169gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n233_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n239_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n227_), .A2(KEYINPUT23), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n224_), .A2(new_n225_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(KEYINPUT23), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n249_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n223_), .B1(new_n246_), .B2(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n234_), .A2(KEYINPUT24), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n240_), .A2(KEYINPUT24), .ZN(new_n258_));
  AND4_X1   g057(.A1(new_n257_), .A2(new_n252_), .A3(new_n244_), .A4(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n249_), .B1(new_n254_), .B2(new_n230_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n222_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n256_), .A2(new_n262_), .A3(KEYINPUT20), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n264_), .B(KEYINPUT95), .Z(new_n265_));
  XOR2_X1   g064(.A(new_n265_), .B(KEYINPUT19), .Z(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n230_), .A2(new_n235_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT97), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n245_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(new_n236_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n255_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n222_), .A3(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n223_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(KEYINPUT20), .A4(new_n266_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n206_), .B1(new_n268_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT20), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n273_), .A2(new_n274_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(new_n223_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n266_), .B1(new_n281_), .B2(new_n262_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n277_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n206_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n202_), .B1(new_n278_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n275_), .A2(new_n276_), .A3(KEYINPUT20), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n267_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(new_n263_), .B2(new_n267_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n284_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n268_), .A2(new_n206_), .A3(new_n277_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(KEYINPUT27), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n286_), .A2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT2), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n300_), .A2(G141gat), .A3(G148gat), .ZN(new_n301_));
  INV_X1    g100(.A(G141gat), .ZN(new_n302_));
  INV_X1    g101(.A(G148gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT3), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n299_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT84), .B1(new_n297_), .B2(new_n298_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT84), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n307_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n296_), .B1(new_n305_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n294_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n296_), .ZN(new_n314_));
  OAI221_X1 g113(.A(new_n313_), .B1(G141gat), .B2(G148gat), .C1(new_n314_), .C2(KEYINPUT1), .ZN(new_n315_));
  AND2_X1   g114(.A1(G127gat), .A2(G134gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G127gat), .A2(G134gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(G113gat), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G127gat), .ZN(new_n319_));
  INV_X1    g118(.A(G134gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G113gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G127gat), .A2(G134gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n318_), .A2(new_n324_), .A3(G120gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(G120gat), .B1(new_n318_), .B2(new_n324_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT3), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n300_), .B1(G141gat), .B2(G148gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n330_), .A2(new_n306_), .A3(new_n308_), .A4(new_n299_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(KEYINPUT85), .A3(new_n296_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n312_), .A2(new_n315_), .A3(new_n327_), .A4(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT98), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n312_), .A2(new_n315_), .A3(new_n332_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT81), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n318_), .A2(new_n324_), .ZN(new_n339_));
  INV_X1    g138(.A(G120gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n318_), .A2(new_n324_), .A3(G120gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(KEYINPUT81), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT98), .B1(new_n336_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n335_), .B1(new_n345_), .B2(new_n333_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n338_), .A2(new_n343_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n312_), .A2(new_n315_), .A3(new_n332_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT4), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n333_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT98), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n334_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(new_n352_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n351_), .B1(new_n355_), .B2(KEYINPUT4), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n347_), .B(KEYINPUT99), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n348_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G57gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G85gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(G1gat), .B(G29gat), .Z(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n348_), .B(new_n364_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n293_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT87), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n331_), .A2(KEYINPUT85), .A3(new_n296_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT85), .B1(new_n331_), .B2(new_n296_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n370_), .B1(new_n373_), .B2(new_n315_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n369_), .B1(new_n374_), .B2(new_n222_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n350_), .A2(KEYINPUT29), .ZN(new_n376_));
  INV_X1    g175(.A(new_n369_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n223_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT90), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n375_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT93), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n377_), .B1(new_n376_), .B2(new_n223_), .ZN(new_n384_));
  AOI211_X1 g183(.A(new_n369_), .B(new_n222_), .C1(new_n350_), .C2(KEYINPUT29), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n379_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G22gat), .B(G50gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n350_), .A2(KEYINPUT29), .A3(new_n391_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n390_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT92), .B(new_n379_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n388_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n383_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n380_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n384_), .A2(new_n385_), .A3(new_n380_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n403_), .B2(KEYINPUT91), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n381_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n382_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n398_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT94), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n401_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n388_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT93), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n382_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n398_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n405_), .B1(new_n406_), .B2(new_n382_), .ZN(new_n416_));
  AOI211_X1 g215(.A(KEYINPUT91), .B(new_n381_), .C1(new_n375_), .C2(new_n378_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT94), .B1(new_n414_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n367_), .B1(new_n410_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT101), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n409_), .B1(new_n401_), .B2(new_n408_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n414_), .A2(KEYINPUT94), .A3(new_n418_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n357_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n346_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n347_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n425_), .B(new_n362_), .C1(new_n356_), .C2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT100), .ZN(new_n428_));
  INV_X1    g227(.A(new_n351_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n429_), .B1(new_n346_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n347_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT100), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n362_), .A4(new_n425_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n278_), .A2(new_n285_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n428_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n365_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n431_), .A2(new_n424_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n439_), .A2(KEYINPUT33), .A3(new_n348_), .A4(new_n364_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n268_), .A2(new_n277_), .A3(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n289_), .A2(KEYINPUT32), .A3(new_n206_), .ZN(new_n445_));
  AOI211_X1 g244(.A(new_n444_), .B(new_n445_), .C1(new_n363_), .C2(new_n365_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n422_), .B(new_n423_), .C1(new_n442_), .C2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n422_), .A2(new_n423_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT101), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n367_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n421_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT31), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G15gat), .B(G43gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT79), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(G71gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n456_));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n455_), .B(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G99gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n261_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(G99gat), .B1(new_n259_), .B2(new_n260_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n459_), .A2(new_n463_), .A3(new_n462_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n452_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n468_), .A3(new_n452_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n344_), .A3(new_n471_), .ZN(new_n472_));
  AOI211_X1 g271(.A(KEYINPUT82), .B(KEYINPUT31), .C1(new_n465_), .C2(new_n466_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n349_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n472_), .A2(KEYINPUT83), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n467_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n451_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n293_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n422_), .A2(new_n482_), .A3(new_n423_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT102), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n366_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n422_), .A2(new_n482_), .A3(new_n423_), .A4(KEYINPUT102), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n479_), .A2(new_n485_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n481_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G190gat), .B(G218gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G134gat), .ZN(new_n492_));
  INV_X1    g291(.A(G162gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n494_), .A2(KEYINPUT36), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT34), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G29gat), .B(G36gat), .ZN(new_n498_));
  INV_X1    g297(.A(G43gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G50gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n498_), .B(G43gat), .ZN(new_n502_));
  INV_X1    g301(.A(G50gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT66), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT66), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n514_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n515_));
  INV_X1    g314(.A(G106gat), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n461_), .B(new_n516_), .C1(new_n512_), .C2(KEYINPUT66), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n511_), .A2(new_n513_), .A3(new_n515_), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G85gat), .ZN(new_n519_));
  INV_X1    g318(.A(G92gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(G85gat), .A2(G92gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT8), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n517_), .A2(new_n515_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n526_), .B(new_n523_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n531_));
  NOR2_X1   g330(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT65), .B1(new_n533_), .B2(new_n521_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n522_), .B1(new_n521_), .B2(KEYINPUT9), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT65), .ZN(new_n536_));
  OAI221_X1 g335(.A(new_n536_), .B1(new_n519_), .B2(new_n520_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT10), .B(G99gat), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n516_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n511_), .A3(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n506_), .A2(new_n530_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT15), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n505_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n501_), .A2(new_n504_), .A3(KEYINPUT15), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n545_), .A2(new_n546_), .B1(new_n530_), .B2(new_n541_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT35), .B(new_n497_), .C1(new_n543_), .C2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n546_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n526_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n529_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n541_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n497_), .A2(KEYINPUT35), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n497_), .A2(KEYINPUT35), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n542_), .A4(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n494_), .B1(new_n548_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n495_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n548_), .A2(new_n556_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(KEYINPUT71), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(KEYINPUT71), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n562_), .B(new_n495_), .C1(new_n558_), .C2(new_n557_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT72), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n490_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n561_), .A2(KEYINPUT72), .A3(new_n563_), .A4(KEYINPUT37), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G1gat), .A2(G8gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT14), .ZN(new_n570_));
  INV_X1    g369(.A(G15gat), .ZN(new_n571_));
  INV_X1    g370(.A(G22gat), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(G15gat), .A2(G22gat), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n570_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n575_), .A2(KEYINPUT73), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G1gat), .B(G8gat), .Z(new_n581_));
  OR2_X1    g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n581_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G57gat), .B(G64gat), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT11), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(KEYINPUT11), .ZN(new_n589_));
  XOR2_X1   g388(.A(G71gat), .B(G78gat), .Z(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n589_), .A2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT74), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n586_), .B(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G183gat), .B(G211gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n595_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n600_), .B(KEYINPUT17), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n595_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n568_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n489_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G229gat), .A2(G233gat), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n582_), .A2(new_n583_), .A3(new_n506_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n584_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n549_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n610_), .B(new_n611_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n610_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n611_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n506_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G113gat), .B(G141gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n232_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(new_n210_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(KEYINPUT76), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(KEYINPUT76), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n624_), .B1(new_n614_), .B2(new_n618_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n530_), .A2(new_n593_), .A3(new_n541_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n593_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n552_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n629_), .A3(KEYINPUT12), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT12), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n552_), .A2(new_n631_), .A3(new_n628_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n634_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n637_));
  XOR2_X1   g436(.A(G120gat), .B(G148gat), .Z(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(G176gat), .B(G204gat), .Z(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n636_), .A2(new_n637_), .A3(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(KEYINPUT68), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT69), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n648_), .B2(KEYINPUT13), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT70), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n609_), .A2(new_n626_), .A3(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n655_), .A2(G1gat), .A3(new_n486_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT38), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(KEYINPUT38), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n623_), .A2(new_n625_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n652_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n489_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n564_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n607_), .A2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n366_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G1gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n658_), .A3(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT103), .ZN(G1324gat));
  OR3_X1    g467(.A1(new_n655_), .A2(G8gat), .A3(new_n482_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n664_), .A2(new_n293_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(G8gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n670_), .B2(G8gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1325gat));
  AOI21_X1  g475(.A(new_n571_), .B1(new_n664_), .B2(new_n479_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT41), .ZN(new_n678_));
  INV_X1    g477(.A(new_n655_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(new_n571_), .A3(new_n479_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1326gat));
  AOI21_X1  g480(.A(new_n572_), .B1(new_n664_), .B2(new_n448_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT42), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n679_), .A2(new_n572_), .A3(new_n448_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1327gat));
  NOR2_X1   g484(.A1(new_n606_), .A2(new_n564_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n661_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(G29gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n366_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n568_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n566_), .A2(KEYINPUT104), .A3(new_n567_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n481_), .B2(new_n488_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n479_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n696_), .A2(new_n486_), .B1(new_n451_), .B2(new_n480_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n568_), .A2(new_n695_), .ZN(new_n698_));
  OAI22_X1  g497(.A1(new_n694_), .A2(new_n695_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n607_), .A3(new_n660_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n699_), .A2(KEYINPUT44), .A3(new_n607_), .A4(new_n660_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n366_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(G29gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n704_), .B2(G29gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n689_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT106), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n710_), .A2(KEYINPUT106), .ZN(new_n712_));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n661_), .A2(new_n713_), .A3(new_n293_), .A4(new_n686_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT45), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n482_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n713_), .B1(new_n717_), .B2(new_n703_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n711_), .B(new_n712_), .C1(new_n716_), .C2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n703_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n721_), .A2(KEYINPUT106), .A3(new_n710_), .A4(new_n715_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1329gat));
  NAND4_X1  g522(.A1(new_n702_), .A2(G43gat), .A3(new_n479_), .A4(new_n703_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n687_), .A2(new_n479_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(G43gat), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n687_), .B2(new_n448_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n703_), .A2(G50gat), .ZN(new_n729_));
  INV_X1    g528(.A(new_n448_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n728_), .B1(new_n729_), .B2(new_n731_), .ZN(G1331gat));
  INV_X1    g531(.A(new_n652_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n626_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n609_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n366_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT107), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n697_), .A2(new_n654_), .A3(new_n626_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n663_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(KEYINPUT108), .A3(new_n663_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT109), .B(G57gat), .Z(new_n744_));
  NOR2_X1   g543(.A1(new_n486_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n737_), .B1(new_n743_), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n741_), .A2(new_n293_), .A3(new_n742_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(G64gat), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n748_), .B2(G64gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n747_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n752_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(KEYINPUT48), .A3(new_n750_), .ZN(new_n755_));
  INV_X1    g554(.A(G64gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n735_), .A2(new_n756_), .A3(new_n293_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n753_), .A2(new_n755_), .A3(new_n757_), .ZN(G1333gat));
  INV_X1    g557(.A(G71gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n735_), .A2(new_n759_), .A3(new_n479_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n743_), .A2(new_n479_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(G71gat), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT49), .B(new_n759_), .C1(new_n743_), .C2(new_n479_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(G1334gat));
  INV_X1    g564(.A(G78gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n735_), .A2(new_n766_), .A3(new_n448_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n743_), .A2(new_n448_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(G78gat), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT50), .B(new_n766_), .C1(new_n743_), .C2(new_n448_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(G1335gat));
  AND2_X1   g571(.A1(new_n738_), .A2(new_n686_), .ZN(new_n773_));
  AOI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n366_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n699_), .A2(new_n607_), .A3(new_n734_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(new_n486_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n774_), .B1(new_n777_), .B2(G85gat), .ZN(G1336gat));
  NAND3_X1  g577(.A1(new_n775_), .A2(G92gat), .A3(new_n293_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n773_), .A2(new_n293_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(G92gat), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT111), .ZN(G1337gat));
  OAI21_X1  g581(.A(G99gat), .B1(new_n776_), .B2(new_n480_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n773_), .A2(new_n539_), .A3(new_n479_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g585(.A1(new_n699_), .A2(new_n607_), .A3(new_n448_), .A4(new_n734_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G106gat), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(KEYINPUT52), .A3(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n773_), .A2(new_n516_), .A3(new_n448_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n788_), .A2(new_n789_), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n792_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT53), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n792_), .A2(new_n798_), .A3(new_n793_), .A4(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1339gat));
  NAND2_X1  g599(.A1(new_n630_), .A2(new_n632_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT55), .B1(new_n801_), .B2(new_n634_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n803_), .B(new_n635_), .C1(new_n630_), .C2(new_n632_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n801_), .A2(new_n634_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n802_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT113), .B1(new_n806_), .B2(new_n644_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n626_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n803_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n633_), .A2(new_n635_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n801_), .A2(KEYINPUT55), .A3(new_n634_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n810_), .B1(new_n814_), .B2(new_n645_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n643_), .B1(new_n815_), .B2(KEYINPUT56), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT114), .B1(new_n809_), .B2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n659_), .B1(new_n815_), .B2(KEYINPUT56), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n807_), .A2(new_n808_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n818_), .A2(new_n819_), .A3(new_n643_), .A4(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n584_), .A2(new_n505_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n615_), .B1(new_n822_), .B2(new_n611_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n622_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT115), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n610_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n622_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n615_), .B(new_n611_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT116), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n825_), .A2(new_n828_), .A3(new_n832_), .A4(new_n829_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n619_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n831_), .A2(new_n833_), .B1(new_n824_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n647_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n817_), .A2(new_n821_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n564_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(KEYINPUT57), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n840_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n837_), .A2(new_n564_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n808_), .B1(new_n806_), .B2(new_n644_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n814_), .A2(KEYINPUT56), .A3(new_n645_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(KEYINPUT118), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n847_), .B(new_n808_), .C1(new_n806_), .C2(new_n644_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n846_), .A2(new_n643_), .A3(new_n835_), .A4(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n831_), .A2(new_n833_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n834_), .A2(new_n824_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n852_), .A2(new_n643_), .A3(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n854_), .A2(new_n846_), .A3(KEYINPUT58), .A4(new_n848_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n855_), .A3(new_n568_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n841_), .A2(new_n843_), .A3(new_n856_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n566_), .A2(new_n606_), .A3(new_n659_), .A4(new_n567_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT54), .B1(new_n858_), .B2(new_n652_), .ZN(new_n859_));
  OR3_X1    g658(.A1(new_n858_), .A2(KEYINPUT54), .A3(new_n652_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n857_), .A2(new_n607_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n696_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n861_), .A2(new_n486_), .A3(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n859_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n837_), .A2(new_n564_), .A3(new_n842_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n842_), .B1(new_n837_), .B2(new_n564_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n856_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n866_), .B1(new_n870_), .B2(new_n606_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n871_), .A2(new_n366_), .A3(new_n696_), .A4(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n865_), .A2(G113gat), .A3(new_n626_), .A4(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n863_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n322_), .B1(new_n876_), .B2(new_n659_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1340gat));
  OAI21_X1  g677(.A(new_n340_), .B1(new_n733_), .B2(KEYINPUT60), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n863_), .B(new_n879_), .C1(KEYINPUT60), .C2(new_n340_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n865_), .A2(new_n653_), .A3(new_n874_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n340_), .ZN(G1341gat));
  OAI211_X1 g681(.A(new_n606_), .B(new_n874_), .C1(new_n863_), .C2(new_n864_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G127gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n863_), .A2(new_n319_), .A3(new_n606_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT120), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n884_), .A2(new_n888_), .A3(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1342gat));
  NAND4_X1  g689(.A1(new_n865_), .A2(G134gat), .A3(new_n568_), .A4(new_n874_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n320_), .B1(new_n876_), .B2(new_n564_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1343gat));
  NOR2_X1   g692(.A1(new_n479_), .A2(new_n730_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n861_), .A2(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n366_), .A3(new_n482_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n659_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n302_), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n654_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT121), .B(G148gat), .Z(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1345gat));
  NOR2_X1   g701(.A1(new_n897_), .A2(new_n607_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT61), .B(G155gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  OAI21_X1  g704(.A(new_n493_), .B1(new_n897_), .B2(new_n564_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n691_), .A2(G162gat), .A3(new_n692_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n897_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT122), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n906_), .B(new_n910_), .C1(new_n897_), .C2(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1347gat));
  NAND2_X1  g711(.A1(new_n626_), .A2(new_n247_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n482_), .A2(new_n366_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n479_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n871_), .A2(new_n730_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n917_), .A2(new_n918_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n914_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n871_), .A2(new_n730_), .A3(new_n626_), .A4(new_n916_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(G169gat), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n924_), .A2(new_n923_), .A3(G169gat), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n922_), .B(KEYINPUT124), .C1(new_n925_), .C2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n926_), .A2(new_n925_), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n871_), .A2(new_n730_), .A3(new_n916_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(KEYINPUT123), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n913_), .B1(new_n931_), .B2(new_n919_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n928_), .B1(new_n929_), .B2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n927_), .A2(new_n933_), .ZN(G1348gat));
  NOR3_X1   g733(.A1(new_n917_), .A2(new_n233_), .A3(new_n654_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT125), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n931_), .A2(new_n919_), .ZN(new_n937_));
  AOI21_X1  g736(.A(G176gat), .B1(new_n937_), .B2(new_n652_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1349gat));
  AOI211_X1 g738(.A(new_n607_), .B(new_n242_), .C1(new_n931_), .C2(new_n919_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G183gat), .B1(new_n930_), .B2(new_n606_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n937_), .A2(new_n662_), .A3(new_n243_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n937_), .A2(new_n568_), .ZN(new_n944_));
  INV_X1    g743(.A(G190gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n943_), .B1(new_n944_), .B2(new_n945_), .ZN(G1351gat));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n947_), .B1(new_n896_), .B2(new_n915_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n871_), .A2(new_n894_), .A3(new_n915_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(KEYINPUT126), .ZN(new_n950_));
  OAI211_X1 g749(.A(G197gat), .B(new_n626_), .C1(new_n948_), .C2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(KEYINPUT127), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n896_), .A2(new_n947_), .A3(new_n915_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n949_), .A2(KEYINPUT126), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n626_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n210_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n955_), .A2(new_n958_), .A3(G197gat), .A4(new_n626_), .ZN(new_n959_));
  AND3_X1   g758(.A1(new_n952_), .A2(new_n957_), .A3(new_n959_), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n955_), .A2(new_n653_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g761(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n963_));
  NAND2_X1  g762(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n964_));
  AND4_X1   g763(.A1(new_n606_), .A2(new_n955_), .A3(new_n963_), .A4(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n963_), .B1(new_n955_), .B2(new_n606_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1354gat));
  AOI21_X1  g766(.A(G218gat), .B1(new_n955_), .B2(new_n662_), .ZN(new_n968_));
  AND2_X1   g767(.A1(new_n955_), .A2(new_n568_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n968_), .B1(G218gat), .B2(new_n969_), .ZN(G1355gat));
endmodule


