//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT19), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT77), .B(G190gat), .Z(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(G183gat), .B2(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT79), .ZN(new_n212_));
  INV_X1    g011(.A(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT23), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n210_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n212_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n209_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT22), .B(G169gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(new_n222_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n208_), .B2(KEYINPUT26), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT25), .B(G183gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n223_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT24), .ZN(new_n235_));
  INV_X1    g034(.A(new_n233_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n235_), .B1(KEYINPUT24), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT78), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n218_), .B1(new_n215_), .B2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n211_), .A2(KEYINPUT78), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n232_), .A2(new_n237_), .A3(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n227_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244_));
  INV_X1    g043(.A(G197gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(G204gat), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n244_), .B(KEYINPUT21), .C1(KEYINPUT84), .C2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G197gat), .B(G204gat), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n244_), .A2(KEYINPUT21), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n250_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT20), .B1(new_n243_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n252_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n225_), .B1(new_n241_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n257_));
  OR3_X1    g056(.A1(new_n257_), .A2(new_n223_), .A3(new_n233_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n230_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n233_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n258_), .A2(new_n219_), .A3(new_n260_), .A4(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT92), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n256_), .A2(new_n262_), .A3(KEYINPUT92), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n254_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n207_), .B1(new_n253_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n252_), .B1(new_n227_), .B2(new_n242_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n256_), .A2(new_n262_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n254_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n269_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n207_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n205_), .B1(new_n268_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT93), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n237_), .A2(new_n241_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n232_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n254_), .B1(new_n226_), .B2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n263_), .A2(new_n252_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT20), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n207_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n226_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n269_), .B1(new_n287_), .B2(new_n254_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n207_), .B1(new_n271_), .B2(new_n252_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(new_n205_), .A3(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT27), .B1(new_n279_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n205_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n273_), .A2(new_n274_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n288_), .A2(new_n289_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n291_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(KEYINPUT27), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n293_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G113gat), .B(G120gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n306_));
  XOR2_X1   g105(.A(G71gat), .B(G99gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G43gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G227gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(G15gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n308_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n243_), .A2(KEYINPUT30), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT30), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n287_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n315_), .A3(new_n312_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n306_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n318_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n320_), .A2(KEYINPUT31), .A3(new_n316_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n305_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT31), .B1(new_n320_), .B2(new_n316_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n317_), .A2(new_n306_), .A3(new_n318_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n304_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(KEYINPUT80), .A3(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(KEYINPUT80), .B2(new_n332_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335_));
  INV_X1    g134(.A(G141gat), .ZN(new_n336_));
  INV_X1    g135(.A(G148gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339_));
  OAI22_X1  g138(.A1(new_n339_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n343_));
  OR3_X1    g142(.A1(new_n334_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n343_), .B1(new_n334_), .B2(new_n342_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n330_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n336_), .A2(new_n337_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n329_), .B1(new_n327_), .B2(KEYINPUT1), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n329_), .A2(KEYINPUT1), .ZN(new_n349_));
  AOI211_X1 g148(.A(new_n347_), .B(new_n331_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n304_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n305_), .B1(new_n346_), .B2(new_n350_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT87), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n352_), .A2(KEYINPUT87), .A3(new_n353_), .A4(new_n354_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT86), .B(KEYINPUT4), .Z(new_n360_));
  OAI211_X1 g159(.A(new_n305_), .B(new_n360_), .C1(new_n346_), .C2(new_n350_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n361_), .A2(G225gat), .A3(G233gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n352_), .A2(KEYINPUT4), .A3(new_n353_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT0), .ZN(new_n367_));
  INV_X1    g166(.A(G57gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G85gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n365_), .A2(new_n371_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n357_), .A2(new_n358_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n371_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n326_), .A2(new_n376_), .ZN(new_n377_));
  OR3_X1    g176(.A1(new_n346_), .A2(KEYINPUT29), .A3(new_n350_), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT28), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT29), .B1(new_n346_), .B2(new_n350_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n254_), .ZN(new_n382_));
  INV_X1    g181(.A(G233gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n384_), .A2(G228gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(G228gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT83), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n382_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n381_), .A2(new_n254_), .A3(new_n388_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n395_));
  XOR2_X1   g194(.A(G22gat), .B(G50gat), .Z(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n394_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n390_), .A2(new_n391_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n392_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n396_), .B1(new_n401_), .B2(new_n393_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n380_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n397_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n379_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n301_), .A2(new_n377_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT95), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n301_), .A2(new_n377_), .A3(new_n407_), .A4(KEYINPUT95), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT94), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n373_), .B(new_n371_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n403_), .A2(new_n414_), .A3(new_n406_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n285_), .A2(new_n207_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n265_), .A2(new_n266_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n252_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n274_), .B1(new_n418_), .B2(new_n288_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n294_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT93), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(new_n278_), .A3(new_n291_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n299_), .B1(new_n422_), .B2(KEYINPUT27), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n413_), .B1(new_n415_), .B2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n403_), .A2(new_n406_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n425_), .A2(new_n301_), .A3(KEYINPUT94), .A4(new_n414_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n268_), .B2(new_n275_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n286_), .A2(new_n290_), .A3(new_n427_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT91), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n286_), .A2(KEYINPUT91), .A3(new_n290_), .A4(new_n427_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n428_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n376_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(KEYINPUT89), .A2(KEYINPUT33), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n437_));
  AND4_X1   g236(.A1(new_n359_), .A2(new_n364_), .A3(new_n374_), .A4(new_n436_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT88), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT33), .ZN(new_n441_));
  OAI22_X1  g240(.A1(new_n439_), .A2(new_n440_), .B1(new_n375_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n363_), .A2(new_n354_), .A3(new_n361_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n352_), .A2(new_n353_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n443_), .B(new_n371_), .C1(new_n444_), .C2(new_n354_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n445_), .A2(KEYINPUT90), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(KEYINPUT90), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n298_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n435_), .B1(new_n442_), .B2(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n424_), .B(new_n426_), .C1(new_n449_), .C2(new_n425_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n412_), .B1(new_n450_), .B2(new_n326_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT64), .B(G106gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n456_), .A2(new_n458_), .B1(KEYINPUT9), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT9), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n462_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT8), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT65), .B1(new_n459_), .B2(new_n460_), .ZN(new_n472_));
  INV_X1    g271(.A(G92gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n370_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G85gat), .A2(G92gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n472_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT7), .ZN(new_n479_));
  INV_X1    g278(.A(G99gat), .ZN(new_n480_));
  INV_X1    g279(.A(G106gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n482_), .A2(new_n467_), .A3(new_n468_), .A4(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n471_), .B1(new_n478_), .B2(new_n484_), .ZN(new_n485_));
  AND4_X1   g284(.A1(new_n471_), .A2(new_n484_), .A3(new_n472_), .A4(new_n477_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n470_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT66), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G57gat), .B(G64gat), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n490_), .A2(KEYINPUT11), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(KEYINPUT11), .ZN(new_n492_));
  XOR2_X1   g291(.A(G71gat), .B(G78gat), .Z(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n492_), .A2(new_n493_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n484_), .A2(new_n472_), .A3(new_n477_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT8), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n484_), .A2(new_n471_), .A3(new_n472_), .A4(new_n477_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(KEYINPUT66), .A3(new_n470_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n489_), .A2(new_n497_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G230gat), .A2(G233gat), .ZN(new_n506_));
  AOI221_X4 g305(.A(new_n488_), .B1(new_n462_), .B2(new_n469_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT66), .B1(new_n501_), .B2(new_n470_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n496_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n497_), .A2(KEYINPUT12), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT67), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G85gat), .B(G92gat), .ZN(new_n513_));
  OAI22_X1  g312(.A1(new_n455_), .A2(new_n457_), .B1(new_n513_), .B2(new_n463_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n512_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n453_), .A2(new_n517_), .A3(new_n454_), .A4(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n461_), .A2(KEYINPUT9), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n469_), .A2(KEYINPUT67), .A3(new_n519_), .A4(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT68), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n522_), .A2(new_n501_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n522_), .B2(new_n501_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n511_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n505_), .A2(new_n506_), .A3(new_n509_), .A4(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n509_), .A2(new_n503_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n506_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G120gat), .B(G148gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(G176gat), .B(G204gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n534_), .B(new_n535_), .Z(new_n536_));
  OR2_X1    g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n536_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(KEYINPUT13), .A3(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT70), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546_));
  INV_X1    g345(.A(G1gat), .ZN(new_n547_));
  INV_X1    g346(.A(G8gat), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT14), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G1gat), .B(G8gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G29gat), .B(G36gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G43gat), .B(G50gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G43gat), .B(G50gat), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n553_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n552_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n559_), .B(new_n561_), .Z(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n562_), .B2(new_n552_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n559_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n552_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT76), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n566_), .B1(new_n569_), .B2(new_n564_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G169gat), .B(G197gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n566_), .B(new_n573_), .C1(new_n569_), .C2(new_n564_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G190gat), .B(G218gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT72), .ZN(new_n580_));
  XOR2_X1   g379(.A(G134gat), .B(G162gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n507_), .A2(new_n508_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(new_n559_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n559_), .B(new_n561_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n522_), .A2(new_n501_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT68), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n522_), .A2(new_n501_), .A3(new_n523_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n589_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(KEYINPUT35), .B(new_n586_), .C1(new_n588_), .C2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n489_), .A2(new_n502_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n567_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n595_), .A2(new_n596_), .A3(new_n598_), .A4(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n594_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n582_), .A2(new_n583_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n584_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n601_), .B(new_n604_), .C1(new_n584_), .C2(new_n602_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT74), .B(KEYINPUT37), .Z(new_n608_));
  AND3_X1   g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n496_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n552_), .B(KEYINPUT75), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT16), .ZN(new_n617_));
  XOR2_X1   g416(.A(G183gat), .B(G211gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT17), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n615_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT17), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n615_), .B1(new_n622_), .B2(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n611_), .A2(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n545_), .A2(new_n578_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n452_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n547_), .A3(new_n376_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT38), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n543_), .A2(new_n578_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n451_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n606_), .A2(new_n607_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT96), .ZN(new_n635_));
  INV_X1    g434(.A(new_n624_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n639_), .B2(new_n414_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n630_), .A2(new_n640_), .ZN(G1324gat));
  AOI21_X1  g440(.A(new_n548_), .B1(new_n638_), .B2(new_n423_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT39), .Z(new_n643_));
  NAND3_X1  g442(.A1(new_n628_), .A2(new_n548_), .A3(new_n423_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g445(.A(new_n326_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n310_), .B1(new_n638_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n649_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n628_), .A2(new_n310_), .A3(new_n647_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(new_n651_), .A3(new_n652_), .ZN(G1326gat));
  OAI21_X1  g452(.A(G22gat), .B1(new_n639_), .B2(new_n407_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT97), .B(KEYINPUT42), .Z(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n655_), .ZN(new_n657_));
  OR3_X1    g456(.A1(new_n627_), .A2(G22gat), .A3(new_n407_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(G1327gat));
  INV_X1    g458(.A(new_n634_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n624_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n633_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G29gat), .B1(new_n662_), .B2(new_n376_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n426_), .A2(new_n424_), .ZN(new_n665_));
  OAI22_X1  g464(.A1(new_n365_), .A2(new_n371_), .B1(KEYINPUT89), .B2(KEYINPUT33), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n373_), .A2(new_n374_), .A3(new_n436_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n440_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n375_), .A2(new_n441_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n448_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n425_), .B1(new_n670_), .B2(new_n434_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n326_), .B1(new_n665_), .B2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n410_), .A2(new_n411_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n611_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n664_), .B1(new_n674_), .B2(KEYINPUT98), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(KEYINPUT43), .C1(new_n451_), .C2(new_n611_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n631_), .A2(new_n636_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT44), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n682_), .B(new_n679_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n376_), .A2(G29gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n663_), .B1(new_n684_), .B2(new_n685_), .ZN(G1328gat));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(KEYINPUT101), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n678_), .A2(new_n680_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n682_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n678_), .A2(KEYINPUT44), .A3(new_n680_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n423_), .A4(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n692_), .B1(new_n684_), .B2(new_n423_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT100), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n691_), .A2(new_n423_), .A3(new_n693_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT99), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(G36gat), .A4(new_n694_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(G36gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n662_), .A2(new_n703_), .A3(new_n423_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT45), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n687_), .A2(KEYINPUT101), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n689_), .B1(new_n702_), .B2(new_n708_), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n707_), .B(new_n688_), .C1(new_n697_), .C2(new_n701_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1329gat));
  XNOR2_X1  g510(.A(KEYINPUT102), .B(G43gat), .ZN(new_n712_));
  INV_X1    g511(.A(new_n662_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n326_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT103), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n684_), .A2(G43gat), .A3(new_n647_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g517(.A1(new_n713_), .A2(G50gat), .A3(new_n407_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n684_), .A2(KEYINPUT104), .A3(new_n425_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G50gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT104), .B1(new_n684_), .B2(new_n425_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(G1331gat));
  NOR3_X1   g522(.A1(new_n451_), .A2(new_n577_), .A3(new_n544_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n637_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G57gat), .B1(new_n725_), .B2(new_n414_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n543_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n577_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n625_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n452_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n376_), .A2(new_n368_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n726_), .B1(new_n731_), .B2(new_n732_), .ZN(G1332gat));
  OAI21_X1  g532(.A(G64gat), .B1(new_n725_), .B2(new_n301_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n301_), .A2(G64gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n731_), .B2(new_n736_), .ZN(G1333gat));
  OAI21_X1  g536(.A(G71gat), .B1(new_n725_), .B2(new_n326_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT49), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n326_), .A2(G71gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n731_), .B2(new_n740_), .ZN(G1334gat));
  OAI21_X1  g540(.A(G78gat), .B1(new_n725_), .B2(new_n407_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT50), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n407_), .A2(G78gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n731_), .B2(new_n744_), .ZN(G1335gat));
  OR2_X1    g544(.A1(new_n678_), .A2(KEYINPUT105), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n678_), .A2(KEYINPUT105), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n729_), .A2(new_n624_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n746_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750_), .B2(new_n414_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n724_), .A2(new_n661_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n370_), .A3(new_n376_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n754_), .ZN(G1336gat));
  OAI21_X1  g554(.A(G92gat), .B1(new_n750_), .B2(new_n301_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(new_n473_), .A3(new_n423_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n750_), .B2(new_n326_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n753_), .A2(new_n456_), .A3(new_n647_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT51), .ZN(G1338gat));
  AND3_X1   g561(.A1(new_n678_), .A2(new_n425_), .A3(new_n748_), .ZN(new_n763_));
  OR3_X1    g562(.A1(new_n763_), .A2(KEYINPUT106), .A3(new_n481_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT106), .B1(new_n763_), .B2(new_n481_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(KEYINPUT52), .A3(new_n765_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n753_), .A2(new_n458_), .A3(new_n425_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n768_), .A2(new_n769_), .A3(new_n773_), .A4(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  NOR2_X1   g574(.A1(new_n636_), .A2(new_n577_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n541_), .A2(new_n542_), .A3(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n611_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n777_), .A2(new_n778_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT108), .B(KEYINPUT54), .Z(new_n781_));
  OR3_X1    g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n569_), .A2(new_n564_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n574_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n570_), .A2(new_n574_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n539_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n527_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n591_), .A2(new_n592_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n793_), .A2(new_n511_), .B1(new_n597_), .B2(new_n496_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n794_), .A2(KEYINPUT55), .A3(new_n506_), .A4(new_n505_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n526_), .A2(new_n509_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT12), .B1(new_n587_), .B2(new_n497_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n529_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n792_), .A2(new_n795_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT110), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n792_), .A2(new_n795_), .A3(new_n798_), .A4(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n536_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n803_), .A2(new_n804_), .A3(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n577_), .A2(new_n538_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT109), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n577_), .A2(new_n538_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n805_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n800_), .A2(new_n802_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n536_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT111), .B1(new_n803_), .B2(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n790_), .B1(new_n811_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n785_), .B1(new_n819_), .B2(new_n634_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n803_), .A2(KEYINPUT56), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n815_), .B(new_n536_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n821_), .A2(new_n822_), .A3(KEYINPUT111), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n814_), .A2(KEYINPUT111), .A3(new_n815_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n807_), .A2(new_n809_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n789_), .B1(new_n823_), .B2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(KEYINPUT57), .A3(new_n660_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n538_), .A2(new_n788_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n611_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT58), .B(new_n829_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n803_), .A2(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n816_), .A2(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n837_), .A2(KEYINPUT112), .A3(KEYINPUT58), .A4(new_n829_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n832_), .A2(new_n835_), .A3(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n820_), .A2(new_n828_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n784_), .B1(new_n840_), .B2(new_n636_), .ZN(new_n841_));
  NOR4_X1   g640(.A1(new_n425_), .A2(new_n423_), .A3(new_n414_), .A4(new_n326_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(KEYINPUT115), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(KEYINPUT115), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT114), .B(KEYINPUT59), .Z(new_n845_));
  OR4_X1    g644(.A1(new_n841_), .A2(new_n843_), .A3(new_n844_), .A4(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n839_), .B(KEYINPUT113), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n820_), .A2(new_n828_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n636_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n784_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n852_), .A2(new_n842_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n846_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n578_), .ZN(new_n856_));
  INV_X1    g655(.A(G113gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n853_), .A2(new_n857_), .A3(new_n577_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1340gat));
  OAI21_X1  g658(.A(G120gat), .B1(new_n855_), .B2(new_n544_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n861_));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n543_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n853_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT116), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n860_), .A2(new_n868_), .A3(new_n865_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(G1341gat));
  OAI21_X1  g669(.A(G127gat), .B1(new_n855_), .B2(new_n636_), .ZN(new_n871_));
  INV_X1    g670(.A(G127gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n853_), .A2(new_n872_), .A3(new_n624_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1342gat));
  AOI21_X1  g673(.A(G134gat), .B1(new_n853_), .B2(new_n635_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n855_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n611_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G134gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT117), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n876_), .B2(new_n879_), .ZN(G1343gat));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n423_), .A2(new_n407_), .A3(new_n647_), .A4(new_n414_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n852_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n784_), .B1(new_n849_), .B2(new_n636_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n882_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT118), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n883_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n577_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT119), .B(G141gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1344gat));
  NAND2_X1  g689(.A1(new_n887_), .A2(new_n545_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g691(.A(new_n887_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT120), .B1(new_n893_), .B2(new_n636_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n887_), .A2(new_n895_), .A3(new_n624_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT61), .B(G155gat), .Z(new_n897_));
  AND3_X1   g696(.A1(new_n894_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n894_), .B2(new_n896_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1346gat));
  AOI21_X1  g699(.A(G162gat), .B1(new_n887_), .B2(new_n635_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n877_), .A2(G162gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT121), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n887_), .B2(new_n903_), .ZN(G1347gat));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n377_), .A2(new_n423_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n407_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n840_), .A2(new_n636_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n851_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n905_), .B1(new_n909_), .B2(new_n577_), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n841_), .A2(KEYINPUT122), .A3(new_n578_), .A4(new_n907_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G169gat), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n912_), .A2(new_n913_), .A3(KEYINPUT62), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n912_), .B2(KEYINPUT62), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n916_), .B(G169gat), .C1(new_n910_), .C2(new_n911_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n914_), .A2(new_n915_), .A3(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n909_), .A2(new_n577_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n224_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(KEYINPUT124), .B1(new_n919_), .B2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n912_), .A2(KEYINPUT62), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n917_), .B1(new_n926_), .B2(new_n913_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n925_), .B(new_n922_), .C1(new_n927_), .C2(new_n914_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n924_), .A2(new_n928_), .ZN(G1348gat));
  INV_X1    g728(.A(new_n909_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n222_), .B1(new_n930_), .B2(new_n727_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n884_), .A2(new_n425_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT125), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n545_), .A2(G176gat), .A3(new_n906_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n931_), .B1(new_n933_), .B2(new_n934_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT126), .ZN(G1349gat));
  NAND3_X1  g735(.A1(new_n909_), .A2(new_n624_), .A3(new_n231_), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT127), .Z(new_n938_));
  NAND2_X1  g737(.A1(new_n906_), .A2(new_n624_), .ZN(new_n939_));
  OR2_X1    g738(.A1(new_n933_), .A2(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n940_), .B2(new_n213_), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n930_), .B2(new_n611_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n909_), .A2(new_n635_), .A3(new_n259_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1351gat));
  NOR4_X1   g743(.A1(new_n884_), .A2(new_n647_), .A3(new_n415_), .A4(new_n301_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n577_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n545_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g748(.A(new_n636_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n945_), .A2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  XOR2_X1   g751(.A(new_n951_), .B(new_n952_), .Z(G1354gat));
  INV_X1    g752(.A(G218gat), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n945_), .A2(new_n954_), .A3(new_n635_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n945_), .A2(new_n877_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n954_), .ZN(G1355gat));
endmodule


