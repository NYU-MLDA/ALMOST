//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_;
  XNOR2_X1  g000(.A(KEYINPUT87), .B(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT26), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204_));
  INV_X1    g003(.A(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n203_), .A2(KEYINPUT88), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(new_n202_), .B2(new_n204_), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT86), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT25), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(new_n209_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(new_n210_), .B2(new_n205_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT89), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT89), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(G169gat), .B2(G176gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n218_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n213_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n218_), .B1(G183gat), .B2(new_n202_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n220_), .A2(new_n221_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n233_), .B2(new_n221_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT30), .ZN(new_n237_));
  INV_X1    g036(.A(G43gat), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n213_), .A2(new_n229_), .B1(new_n234_), .B2(new_n231_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT30), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n238_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n238_), .B1(new_n237_), .B2(new_n241_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G227gat), .A2(G233gat), .ZN(new_n245_));
  INV_X1    g044(.A(G15gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n241_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n239_), .A2(new_n240_), .ZN(new_n251_));
  OAI21_X1  g050(.A(G43gat), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n247_), .B1(new_n252_), .B2(new_n242_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G71gat), .B(G99gat), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n249_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n254_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n248_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n252_), .A2(new_n247_), .A3(new_n242_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT90), .ZN(new_n260_));
  INV_X1    g059(.A(G120gat), .ZN(new_n261_));
  OR2_X1    g060(.A1(G127gat), .A2(G134gat), .ZN(new_n262_));
  INV_X1    g061(.A(G113gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G127gat), .A2(G134gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n263_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n261_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(G120gat), .A3(new_n265_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT91), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT31), .ZN(new_n273_));
  OAI22_X1  g072(.A1(new_n255_), .A2(new_n259_), .B1(new_n260_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n254_), .B1(new_n249_), .B2(new_n253_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n273_), .A2(new_n260_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n257_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281_));
  INV_X1    g080(.A(G141gat), .ZN(new_n282_));
  INV_X1    g081(.A(G148gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n284_), .A2(new_n287_), .A3(new_n288_), .A4(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT92), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n291_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n294_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(KEYINPUT92), .A3(new_n292_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n290_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(new_n299_), .A3(new_n292_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n282_), .A2(new_n283_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(KEYINPUT1), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .A4(new_n285_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n298_), .A2(new_n303_), .A3(KEYINPUT93), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT93), .B1(new_n298_), .B2(new_n303_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT29), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT21), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G197gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(G204gat), .ZN(new_n311_));
  INV_X1    g110(.A(G204gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n312_), .A2(G197gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT21), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n309_), .A2(new_n314_), .A3(KEYINPUT96), .A4(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(KEYINPUT96), .ZN(new_n317_));
  INV_X1    g116(.A(new_n307_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(KEYINPUT21), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G228gat), .A2(G233gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT95), .Z(new_n322_));
  NAND3_X1  g121(.A1(new_n306_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT97), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n298_), .A2(new_n303_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT29), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n320_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n322_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n324_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  AOI211_X1 g128(.A(KEYINPUT97), .B(new_n322_), .C1(new_n326_), .C2(new_n320_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n323_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT98), .B(G78gat), .ZN(new_n332_));
  INV_X1    g131(.A(G106gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n323_), .B(new_n334_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(KEYINPUT94), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT93), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n325_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n298_), .A2(new_n303_), .A3(KEYINPUT93), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(KEYINPUT29), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n336_), .A2(KEYINPUT94), .A3(new_n345_), .A4(new_n337_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G22gat), .B(G50gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT28), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n344_), .A2(new_n349_), .A3(new_n346_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n342_), .A2(new_n356_), .A3(new_n271_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n271_), .A2(new_n325_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n342_), .B2(new_n271_), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT101), .B1(new_n359_), .B2(KEYINPUT4), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n271_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n271_), .A2(new_n325_), .ZN(new_n362_));
  AND4_X1   g161(.A1(KEYINPUT101), .A2(new_n361_), .A3(new_n362_), .A4(KEYINPUT4), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n355_), .B(new_n357_), .C1(new_n360_), .C2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT102), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n359_), .A2(new_n354_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT101), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n362_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(new_n356_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n359_), .A2(KEYINPUT101), .A3(KEYINPUT4), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT102), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n355_), .A4(new_n357_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n365_), .A2(new_n366_), .A3(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT0), .B(G57gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G85gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(G1gat), .B(G29gat), .Z(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n365_), .A2(new_n380_), .A3(new_n366_), .A4(new_n373_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n316_), .A2(new_n319_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT26), .B(G190gat), .ZN(new_n384_));
  OR2_X1    g183(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT99), .ZN(new_n386_));
  NAND2_X1  g185(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n384_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n217_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT100), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n232_), .B2(new_n225_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n227_), .A2(KEYINPUT100), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n390_), .A2(new_n391_), .A3(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n234_), .B1(new_n217_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n383_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(KEYINPUT20), .C1(new_n239_), .C2(new_n383_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT19), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n239_), .A2(new_n383_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n396_), .A2(new_n398_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n320_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n405_), .A2(new_n407_), .A3(KEYINPUT20), .A4(new_n402_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT18), .B(G64gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G92gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G8gat), .B(G36gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT32), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n400_), .A2(new_n402_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n405_), .A2(new_n407_), .A3(KEYINPUT20), .A4(new_n403_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n415_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT103), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n416_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n409_), .A2(KEYINPUT103), .A3(new_n415_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n382_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n365_), .A2(new_n373_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n424_), .A2(KEYINPUT33), .A3(new_n380_), .A4(new_n366_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n378_), .B1(new_n368_), .B2(new_n354_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n357_), .A2(new_n354_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n371_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n413_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n404_), .A2(new_n413_), .A3(new_n408_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n381_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n425_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n353_), .B1(new_n423_), .B2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n414_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n429_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n430_), .B2(new_n429_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT104), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(KEYINPUT104), .B(new_n437_), .C1(new_n430_), .C2(new_n429_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n438_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n344_), .A2(new_n349_), .A3(new_n346_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n349_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n444_), .A2(new_n447_), .A3(new_n382_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n280_), .B1(new_n435_), .B2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n379_), .A2(new_n381_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n450_), .A2(new_n447_), .A3(new_n279_), .A4(new_n443_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT105), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n443_), .A2(new_n352_), .A3(new_n351_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT105), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n450_), .A4(new_n279_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n449_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT65), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT65), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT6), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n459_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G85gat), .B(G92gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT9), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT10), .B(G99gat), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n467_), .B(new_n470_), .C1(G106gat), .C2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT9), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G85gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n472_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT69), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(KEYINPUT6), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n460_), .A2(KEYINPUT69), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n458_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G99gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n333_), .A3(KEYINPUT66), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT7), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT7), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(new_n485_), .A3(new_n333_), .A4(KEYINPUT66), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n460_), .A2(KEYINPUT69), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n481_), .A2(KEYINPUT6), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n459_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n484_), .A2(new_n487_), .A3(new_n489_), .A4(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT70), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n469_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n494_), .B1(new_n493_), .B2(new_n469_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n467_), .A2(KEYINPUT67), .A3(new_n487_), .A4(new_n489_), .ZN(new_n499_));
  OR2_X1    g298(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n500_));
  NAND2_X1  g299(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n468_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n461_), .A2(new_n463_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n458_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n504_), .A2(new_n464_), .A3(new_n487_), .A4(new_n489_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT67), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n499_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n480_), .B1(new_n498_), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G57gat), .B(G64gat), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G71gat), .B(G78gat), .ZN(new_n513_));
  OR3_X1    g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n513_), .A3(KEYINPUT11), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n509_), .A2(KEYINPUT12), .A3(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n493_), .A2(new_n469_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT70), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n493_), .A2(new_n494_), .A3(new_n469_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(KEYINPUT8), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n499_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n479_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n519_), .B1(new_n525_), .B2(new_n516_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G230gat), .A2(G233gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n525_), .B2(new_n516_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n518_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT73), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n526_), .A2(new_n518_), .A3(new_n529_), .A4(KEYINPUT73), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT71), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n523_), .A2(new_n524_), .ZN(new_n536_));
  AND4_X1   g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n480_), .A4(new_n516_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n535_), .B1(new_n525_), .B2(new_n516_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n525_), .A2(new_n516_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n528_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G120gat), .B(G148gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(new_n312_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT5), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n221_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n534_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n534_), .B2(new_n541_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT13), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n534_), .A2(new_n541_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n545_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n534_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT13), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n548_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT77), .B(G1gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT78), .B(G8gat), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT14), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G1gat), .B(G8gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n564_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n559_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n562_), .A2(new_n565_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n563_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(new_n558_), .A3(new_n566_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G29gat), .B(G36gat), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(G43gat), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(G43gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(G50gat), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(G50gat), .B1(new_n575_), .B2(new_n576_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n573_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n569_), .A2(new_n580_), .A3(new_n572_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n557_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT84), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(new_n220_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n310_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT15), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n579_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(KEYINPUT15), .A3(new_n577_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n569_), .A2(new_n572_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n557_), .B(new_n583_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n596_), .A2(KEYINPUT84), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n585_), .B(new_n589_), .C1(new_n597_), .C2(new_n584_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n582_), .A2(new_n583_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n557_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n596_), .A2(KEYINPUT84), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n599_), .A2(KEYINPUT84), .A3(new_n600_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n588_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n598_), .A2(new_n603_), .A3(KEYINPUT85), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT85), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n605_), .B(new_n588_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n556_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n569_), .A2(new_n572_), .A3(new_n610_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n517_), .A3(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n569_), .A2(new_n572_), .A3(new_n610_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n516_), .B1(new_n615_), .B2(new_n611_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT17), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n614_), .A2(new_n616_), .A3(new_n617_), .A4(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT82), .B1(new_n614_), .B2(new_n616_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n617_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  AOI211_X1 g426(.A(KEYINPUT82), .B(new_n627_), .C1(new_n614_), .C2(new_n616_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n623_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT83), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT83), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n631_), .B(new_n623_), .C1(new_n626_), .C2(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(G134gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(G162gat), .Z(new_n637_));
  INV_X1    g436(.A(KEYINPUT36), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n525_), .A2(new_n594_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT35), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G232gat), .A2(G233gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT74), .Z(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT34), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n525_), .A2(new_n580_), .B1(new_n641_), .B2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n641_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT75), .Z(new_n647_));
  NAND4_X1  g446(.A1(new_n640_), .A2(new_n645_), .A3(KEYINPUT76), .A4(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT76), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(new_n641_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n650_), .B(new_n651_), .C1(new_n509_), .C2(new_n581_), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n652_), .A2(new_n647_), .B1(new_n640_), .B2(new_n645_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n639_), .B1(new_n649_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n647_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n640_), .A2(new_n645_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n637_), .B(new_n638_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n648_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT37), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n654_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n654_), .B2(new_n659_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n609_), .A2(new_n634_), .A3(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n457_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT106), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(new_n457_), .B2(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n560_), .A3(new_n382_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT107), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n669_), .A2(new_n672_), .A3(new_n560_), .A4(new_n382_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n654_), .A2(new_n659_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT108), .Z(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n457_), .A2(new_n633_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n609_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n382_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n674_), .A2(KEYINPUT38), .B1(G1gat), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n683_), .B1(new_n674_), .B2(KEYINPUT38), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n671_), .A2(new_n673_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT38), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(KEYINPUT109), .A3(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n682_), .A2(new_n684_), .A3(new_n687_), .ZN(G1324gat));
  NAND3_X1  g487(.A1(new_n669_), .A2(new_n444_), .A3(new_n561_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G8gat), .B1(new_n679_), .B2(new_n443_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(KEYINPUT39), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(KEYINPUT39), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1325gat));
  NAND3_X1  g494(.A1(new_n665_), .A2(new_n246_), .A3(new_n279_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n680_), .A2(new_n279_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n697_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT41), .B1(new_n697_), .B2(G15gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT110), .B(new_n696_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1326gat));
  OAI21_X1  g503(.A(G22gat), .B1(new_n679_), .B2(new_n447_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT42), .ZN(new_n706_));
  INV_X1    g505(.A(G22gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n665_), .A2(new_n707_), .A3(new_n353_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1327gat));
  INV_X1    g508(.A(new_n675_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n449_), .B2(new_n456_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n556_), .A2(new_n608_), .A3(new_n634_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n713_), .A2(G29gat), .A3(new_n450_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n449_), .A2(new_n456_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n663_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  AOI211_X1 g517(.A(KEYINPUT43), .B(new_n663_), .C1(new_n449_), .C2(new_n456_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n712_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n712_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n382_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n714_), .B1(new_n725_), .B2(G29gat), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT111), .B(new_n714_), .C1(new_n725_), .C2(G29gat), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1328gat));
  NAND3_X1  g529(.A1(new_n722_), .A2(new_n444_), .A3(new_n723_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G36gat), .ZN(new_n732_));
  INV_X1    g531(.A(G36gat), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n711_), .A2(new_n712_), .A3(new_n733_), .A4(new_n444_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n732_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT112), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n732_), .A2(new_n740_), .A3(new_n737_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(KEYINPUT46), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n740_), .B1(new_n732_), .B2(new_n737_), .ZN(new_n744_));
  AOI211_X1 g543(.A(KEYINPUT112), .B(new_n736_), .C1(new_n731_), .C2(G36gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n742_), .A2(new_n746_), .ZN(G1329gat));
  NAND3_X1  g546(.A1(new_n724_), .A2(G43gat), .A3(new_n279_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n238_), .B1(new_n713_), .B2(new_n280_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g550(.A(G50gat), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n447_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n711_), .A2(new_n353_), .A3(new_n712_), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n724_), .A2(new_n753_), .B1(new_n752_), .B2(new_n754_), .ZN(G1331gat));
  NOR2_X1   g554(.A1(new_n555_), .A2(new_n607_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n633_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n716_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G57gat), .B1(new_n758_), .B2(new_n382_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n678_), .A2(new_n756_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(new_n382_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n759_), .B1(new_n761_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g561(.A(G64gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n760_), .B2(new_n444_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT48), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n758_), .A2(new_n763_), .A3(new_n444_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1333gat));
  INV_X1    g566(.A(G71gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n760_), .B2(new_n279_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT49), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n758_), .A2(new_n768_), .A3(new_n279_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1334gat));
  NAND2_X1  g571(.A1(new_n760_), .A2(new_n353_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G78gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT113), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n776_), .A3(G78gat), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(G78gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n758_), .A2(new_n781_), .A3(new_n353_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n775_), .A2(KEYINPUT50), .A3(new_n777_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(new_n782_), .A3(new_n783_), .ZN(G1335gat));
  NAND2_X1  g583(.A1(new_n756_), .A2(new_n633_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n711_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(G85gat), .B1(new_n787_), .B2(new_n382_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n718_), .A2(new_n719_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(new_n382_), .A3(new_n786_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n788_), .B1(new_n791_), .B2(G85gat), .ZN(G1336gat));
  NAND2_X1  g591(.A1(new_n789_), .A2(new_n786_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n444_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n787_), .A2(new_n444_), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n793_), .A2(new_n794_), .B1(G92gat), .B2(new_n795_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT114), .Z(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n793_), .B2(new_n280_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n471_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n787_), .A2(new_n279_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n787_), .A2(new_n333_), .A3(new_n353_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n789_), .A2(new_n353_), .A3(new_n786_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n804_), .A2(new_n805_), .A3(G106gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n804_), .B2(G106gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n534_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n530_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n526_), .B(new_n518_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(KEYINPUT55), .A2(new_n813_), .B1(new_n814_), .B2(new_n528_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n810_), .B1(new_n816_), .B2(new_n550_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT55), .B1(new_n532_), .B2(new_n533_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n518_), .A2(new_n526_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n528_), .B1(new_n539_), .B2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n526_), .A2(new_n518_), .A3(new_n529_), .A4(KEYINPUT55), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n810_), .B(new_n550_), .C1(new_n818_), .C2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n817_), .A2(new_n824_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n601_), .A2(new_n602_), .A3(new_n588_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n599_), .A2(new_n557_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n600_), .B(new_n583_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n828_), .A2(new_n588_), .A3(new_n829_), .ZN(new_n830_));
  OR3_X1    g629(.A1(new_n826_), .A2(new_n827_), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n825_), .A2(KEYINPUT58), .A3(new_n552_), .A4(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n550_), .B1(new_n818_), .B2(new_n822_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT56), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(new_n833_), .A3(new_n552_), .A4(new_n823_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n834_), .A2(new_n717_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT119), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n836_), .A2(new_n607_), .A3(new_n552_), .A4(new_n823_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n833_), .B1(new_n547_), .B2(new_n546_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n710_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n675_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n834_), .A2(new_n850_), .A3(new_n839_), .A4(new_n717_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n841_), .A2(new_n849_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n633_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n757_), .A2(new_n555_), .A3(new_n608_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT54), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT116), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n857_), .A3(KEYINPUT54), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n854_), .B2(KEYINPUT54), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n607_), .B1(new_n548_), .B2(new_n554_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n861_), .A2(KEYINPUT115), .A3(new_n862_), .A4(new_n757_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n856_), .A2(new_n858_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n853_), .A2(new_n865_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n453_), .A2(new_n382_), .A3(new_n279_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G113gat), .B1(new_n869_), .B2(new_n607_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n634_), .B1(new_n849_), .B2(new_n840_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n871_), .A2(new_n864_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n867_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n869_), .B2(new_n873_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n263_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n870_), .B1(new_n876_), .B2(new_n607_), .ZN(G1340gat));
  OAI21_X1  g676(.A(G120gat), .B1(new_n875_), .B2(new_n555_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n261_), .B1(new_n555_), .B2(KEYINPUT60), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n869_), .B(new_n879_), .C1(KEYINPUT60), .C2(new_n261_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1341gat));
  AOI21_X1  g680(.A(G127gat), .B1(new_n869_), .B2(new_n634_), .ZN(new_n882_));
  INV_X1    g681(.A(G127gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n875_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n884_), .B2(new_n634_), .ZN(G1342gat));
  AOI21_X1  g684(.A(G134gat), .B1(new_n869_), .B2(new_n677_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n875_), .A2(new_n663_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g687(.A1(new_n280_), .A2(new_n353_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n889_), .A2(new_n450_), .A3(new_n444_), .ZN(new_n890_));
  XOR2_X1   g689(.A(new_n890_), .B(KEYINPUT120), .Z(new_n891_));
  NAND2_X1  g690(.A1(new_n866_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n608_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n282_), .ZN(G1344gat));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n555_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n283_), .ZN(G1345gat));
  XOR2_X1   g695(.A(KEYINPUT61), .B(G155gat), .Z(new_n897_));
  OR3_X1    g696(.A1(new_n892_), .A2(new_n633_), .A3(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT121), .B(KEYINPUT122), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n892_), .B2(new_n633_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n898_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1346gat));
  INV_X1    g702(.A(new_n892_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G162gat), .B1(new_n904_), .B2(new_n677_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n892_), .A2(new_n663_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(G162gat), .B2(new_n906_), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n382_), .A2(new_n443_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n280_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n447_), .B(new_n910_), .C1(new_n871_), .C2(new_n864_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n911_), .A2(new_n608_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G169gat), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n912_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n916_));
  INV_X1    g715(.A(new_n233_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n915_), .B(new_n916_), .C1(new_n917_), .C2(new_n912_), .ZN(G1348gat));
  AOI21_X1  g717(.A(new_n864_), .B1(new_n852_), .B2(new_n633_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n353_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n920_), .A2(G176gat), .A3(new_n556_), .A4(new_n910_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n872_), .A2(new_n447_), .A3(new_n556_), .A4(new_n910_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n221_), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n922_), .B(new_n221_), .C1(new_n911_), .C2(new_n555_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n921_), .B1(new_n924_), .B2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT124), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n929_), .B(new_n921_), .C1(new_n924_), .C2(new_n926_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1349gat));
  OR4_X1    g730(.A1(new_n389_), .A2(new_n911_), .A3(new_n388_), .A4(new_n633_), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n920_), .A2(new_n634_), .A3(new_n910_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(G183gat), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n932_), .B(KEYINPUT125), .C1(G183gat), .C2(new_n933_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1350gat));
  OAI21_X1  g737(.A(G190gat), .B1(new_n911_), .B2(new_n663_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n677_), .A2(new_n384_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n911_), .B2(new_n940_), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n889_), .A2(new_n909_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n866_), .A2(KEYINPUT126), .A3(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944_));
  INV_X1    g743(.A(new_n942_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n919_), .B2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n943_), .A2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n607_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n556_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n952_), .B1(new_n947_), .B2(new_n634_), .ZN(new_n953_));
  XOR2_X1   g752(.A(KEYINPUT63), .B(G211gat), .Z(new_n954_));
  AOI211_X1 g753(.A(new_n633_), .B(new_n954_), .C1(new_n943_), .C2(new_n946_), .ZN(new_n955_));
  OAI21_X1  g754(.A(KEYINPUT127), .B1(new_n953_), .B2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n954_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n947_), .A2(new_n634_), .A3(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n633_), .B1(new_n943_), .B2(new_n946_), .ZN(new_n960_));
  OAI211_X1 g759(.A(new_n958_), .B(new_n959_), .C1(new_n960_), .C2(new_n952_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n956_), .A2(new_n961_), .ZN(G1354gat));
  AOI21_X1  g761(.A(G218gat), .B1(new_n947_), .B2(new_n677_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n663_), .B1(new_n943_), .B2(new_n946_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n963_), .B1(G218gat), .B2(new_n964_), .ZN(G1355gat));
endmodule


