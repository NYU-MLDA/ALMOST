//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n821_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G43gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G227gat), .A2(G233gat), .ZN(new_n204_));
  INV_X1    g003(.A(G15gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n203_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(new_n209_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT84), .ZN(new_n213_));
  MUX2_X1   g012(.A(new_n209_), .B(new_n212_), .S(new_n213_), .Z(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(G183gat), .B2(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT82), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT22), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(KEYINPUT22), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n216_), .B(new_n219_), .C1(new_n220_), .C2(new_n217_), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n221_), .A2(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n215_), .B(new_n222_), .C1(KEYINPUT83), .C2(new_n221_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n216_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT81), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT24), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT25), .B(G183gat), .ZN(new_n231_));
  INV_X1    g030(.A(G190gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT80), .B1(new_n232_), .B2(KEYINPUT26), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT26), .B(G190gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n231_), .B(new_n233_), .C1(new_n234_), .C2(KEYINPUT80), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n228_), .A2(new_n230_), .A3(new_n212_), .A4(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n223_), .A2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT30), .Z(new_n238_));
  INV_X1    g037(.A(KEYINPUT85), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n207_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n207_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n245_), .A2(KEYINPUT86), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(KEYINPUT86), .ZN(new_n247_));
  XOR2_X1   g046(.A(G113gat), .B(G120gat), .Z(new_n248_));
  OR3_X1    g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n248_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OR3_X1    g053(.A1(new_n242_), .A2(new_n244_), .A3(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G155gat), .A2(G162gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT88), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(KEYINPUT2), .ZN(new_n262_));
  OR2_X1    g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT3), .ZN(new_n264_));
  OR3_X1    g063(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT2), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n264_), .B(new_n265_), .C1(new_n266_), .C2(new_n260_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n258_), .B(new_n259_), .C1(new_n262_), .C2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n263_), .B(KEYINPUT89), .ZN(new_n269_));
  INV_X1    g068(.A(new_n261_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n258_), .A2(KEYINPUT1), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n258_), .A2(KEYINPUT1), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(new_n259_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n268_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n275_), .A2(KEYINPUT29), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT28), .ZN(new_n277_));
  XOR2_X1   g076(.A(G22gat), .B(G50gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT90), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G197gat), .B(G204gat), .Z(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(KEYINPUT21), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(KEYINPUT21), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G211gat), .B(G218gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n275_), .B2(KEYINPUT29), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G228gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G78gat), .B(G106gat), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n293_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n279_), .A2(new_n280_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n281_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n295_), .A2(KEYINPUT91), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(KEYINPUT91), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(new_n279_), .A3(new_n294_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n275_), .A2(new_n251_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n275_), .A2(new_n251_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(KEYINPUT4), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n307_), .B(KEYINPUT99), .Z(new_n308_));
  AND2_X1   g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n275_), .A2(new_n251_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT100), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n304_), .A2(new_n305_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n309_), .A2(new_n313_), .B1(new_n314_), .B2(new_n307_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G1gat), .B(G29gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(G85gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT0), .B(G57gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  OR2_X1    g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n319_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n237_), .A2(new_n288_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n212_), .B1(G183gat), .B2(G190gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT93), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT22), .B(G169gat), .Z(new_n327_));
  OAI21_X1  g126(.A(new_n226_), .B1(new_n327_), .B2(G176gat), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n234_), .A2(new_n231_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n228_), .A2(new_n230_), .A3(new_n214_), .A4(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n289_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n323_), .A2(new_n332_), .A3(KEYINPUT20), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n331_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n326_), .A2(new_n328_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n288_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n340_), .B(KEYINPUT20), .C1(new_n288_), .C2(new_n237_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n337_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT96), .ZN(new_n344_));
  XOR2_X1   g143(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n342_), .A2(KEYINPUT32), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n341_), .A2(new_n336_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT94), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n332_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT20), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n336_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n329_), .A2(KEYINPUT94), .A3(new_n289_), .A4(new_n331_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .A4(new_n323_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n348_), .A2(KEYINPUT32), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n350_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n322_), .A2(new_n349_), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n313_), .A2(new_n307_), .A3(new_n306_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n319_), .B1(new_n314_), .B2(new_n308_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n315_), .A2(new_n363_), .A3(new_n319_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n362_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n350_), .A2(new_n356_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n348_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n350_), .A2(new_n356_), .A3(new_n348_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(KEYINPUT97), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT97), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n368_), .A2(new_n373_), .A3(new_n369_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT98), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n372_), .A2(KEYINPUT98), .A3(new_n374_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n367_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT101), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n359_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n365_), .A2(new_n366_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n372_), .A2(KEYINPUT98), .A3(new_n374_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT98), .B1(new_n372_), .B2(new_n374_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n362_), .B(new_n382_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(KEYINPUT101), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n303_), .B1(new_n381_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n322_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n302_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT27), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n372_), .A2(new_n390_), .A3(new_n374_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n342_), .A2(new_n369_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(KEYINPUT27), .A3(new_n371_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n257_), .B1(new_n387_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n322_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT102), .B1(new_n391_), .B2(new_n393_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n391_), .A2(KEYINPUT102), .A3(new_n393_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n398_), .B(new_n303_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT103), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT10), .B(G99gat), .Z(new_n404_));
  INV_X1    g203(.A(G106gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407_));
  INV_X1    g206(.A(G99gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(new_n405_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G85gat), .A2(G92gat), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n412_), .A2(KEYINPUT9), .ZN(new_n413_));
  INV_X1    g212(.A(G85gat), .ZN(new_n414_));
  INV_X1    g213(.A(G92gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(KEYINPUT9), .A3(new_n412_), .ZN(new_n417_));
  AND4_X1   g216(.A1(new_n406_), .A2(new_n411_), .A3(new_n413_), .A4(new_n417_), .ZN(new_n418_));
  OR3_X1    g217(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(new_n409_), .A3(new_n410_), .A4(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n416_), .A2(new_n412_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT8), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT8), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n421_), .A2(new_n425_), .A3(new_n422_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n418_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT11), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT64), .ZN(new_n429_));
  INV_X1    g228(.A(G57gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n430_), .A2(G64gat), .ZN(new_n431_));
  INV_X1    g230(.A(G64gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(G57gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n429_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(G57gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n430_), .A2(G64gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(KEYINPUT64), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n428_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n434_), .A2(new_n428_), .A3(new_n437_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT65), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G71gat), .B(G78gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n440_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n441_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n439_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n435_), .A2(new_n436_), .A3(KEYINPUT64), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT64), .B1(new_n435_), .B2(new_n436_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT11), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT65), .B1(new_n449_), .B2(new_n442_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n440_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n438_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n427_), .B1(new_n446_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT68), .B1(new_n453_), .B2(KEYINPUT12), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n424_), .A2(new_n426_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n418_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n444_), .A2(new_n445_), .A3(new_n439_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n438_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT68), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(KEYINPUT12), .B(new_n457_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n453_), .A2(KEYINPUT67), .A3(KEYINPUT12), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n454_), .A2(new_n463_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n446_), .A2(new_n452_), .A3(new_n427_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G230gat), .A2(G233gat), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT66), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n469_), .B(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n474_), .A2(new_n460_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n472_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(G120gat), .B(G148gat), .Z(new_n477_));
  XNOR2_X1  g276(.A(G176gat), .B(G204gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n476_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT13), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n483_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G29gat), .B(G36gat), .Z(new_n487_));
  XOR2_X1   g286(.A(G43gat), .B(G50gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n489_), .B(KEYINPUT79), .Z(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G8gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT75), .ZN(new_n492_));
  INV_X1    g291(.A(G22gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n205_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G15gat), .A2(G22gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G1gat), .A2(G8gat), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n494_), .A2(new_n495_), .B1(KEYINPUT14), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n492_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n490_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G229gat), .A2(G233gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n489_), .B(KEYINPUT15), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n498_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n502_), .B1(new_n490_), .B2(new_n499_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n500_), .A2(new_n502_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G113gat), .B(G141gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n506_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n486_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n403_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n458_), .A2(new_n459_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G231gat), .A2(G233gat), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n515_), .A2(new_n516_), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n499_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n499_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G127gat), .B(G155gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(G183gat), .B(G211gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .A4(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT77), .B1(new_n519_), .B2(new_n521_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n526_), .A2(new_n520_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n528_), .A2(new_n529_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n527_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT78), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n503_), .A2(new_n457_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n427_), .A2(new_n489_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n537_), .B2(KEYINPUT71), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n540_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT72), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT73), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n549_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n553_), .B(KEYINPUT36), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n546_), .A2(new_n548_), .A3(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(KEYINPUT37), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n558_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT74), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(new_n549_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n563_), .B2(new_n549_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n557_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n561_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n536_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n514_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(G1gat), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n572_), .A3(new_n322_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT38), .ZN(new_n574_));
  INV_X1    g373(.A(new_n566_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n257_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n359_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n385_), .B2(KEYINPUT101), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n379_), .A2(new_n380_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n302_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n576_), .B1(new_n580_), .B2(new_n395_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT103), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n401_), .B(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n575_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n513_), .A2(new_n536_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT104), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G1gat), .B1(new_n588_), .B2(new_n388_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n574_), .A2(new_n589_), .ZN(G1324gat));
  INV_X1    g389(.A(G8gat), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n400_), .A2(new_n399_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n571_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n594_));
  INV_X1    g393(.A(new_n586_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n592_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n594_), .B1(new_n596_), .B2(G8gat), .ZN(new_n597_));
  AOI211_X1 g396(.A(KEYINPUT39), .B(new_n591_), .C1(new_n595_), .C2(new_n592_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n593_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g399(.A(new_n205_), .B1(new_n587_), .B2(new_n257_), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n571_), .A2(new_n205_), .A3(new_n257_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(G1326gat));
  NAND3_X1  g405(.A1(new_n571_), .A2(new_n493_), .A3(new_n302_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G22gat), .B1(new_n588_), .B2(new_n303_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n608_), .A2(KEYINPUT42), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(KEYINPUT42), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(G1327gat));
  INV_X1    g410(.A(new_n536_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(new_n566_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n512_), .B(new_n613_), .C1(new_n397_), .C2(new_n402_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT108), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n615_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(G29gat), .B1(new_n618_), .B2(new_n322_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n512_), .A2(new_n536_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n568_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT43), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n622_), .A2(KEYINPUT106), .A3(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n569_), .B1(new_n397_), .B2(new_n402_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT106), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT43), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT44), .B(new_n621_), .C1(new_n624_), .C2(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n628_), .A2(G29gat), .A3(new_n322_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n623_), .B1(new_n622_), .B2(KEYINPUT106), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n625_), .A2(new_n626_), .A3(KEYINPUT43), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n620_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n619_), .B1(new_n629_), .B2(new_n634_), .ZN(G1328gat));
  OAI211_X1 g434(.A(new_n628_), .B(new_n592_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G36gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n592_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(G36gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n616_), .A2(new_n617_), .A3(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT45), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n637_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT46), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n637_), .A2(new_n641_), .A3(KEYINPUT46), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1329gat));
  NAND2_X1  g445(.A1(new_n616_), .A2(new_n617_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n647_), .A2(G43gat), .A3(new_n576_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n628_), .B(new_n257_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n649_), .B2(G43gat), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT47), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT47), .B(new_n648_), .C1(new_n649_), .C2(G43gat), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1330gat));
  AND4_X1   g453(.A1(G50gat), .A2(new_n634_), .A3(new_n302_), .A4(new_n628_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G50gat), .B1(new_n618_), .B2(new_n302_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1331gat));
  INV_X1    g456(.A(new_n486_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n534_), .A2(new_n535_), .A3(new_n511_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n584_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n584_), .A2(KEYINPUT109), .A3(new_n660_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n322_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G57gat), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n403_), .A2(new_n510_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n667_), .A2(new_n486_), .A3(new_n570_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(new_n430_), .A3(new_n322_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT110), .Z(G1332gat));
  NAND3_X1  g470(.A1(new_n668_), .A2(new_n432_), .A3(new_n592_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT48), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n663_), .A2(new_n664_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n592_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n675_), .B2(G64gat), .ZN(new_n676_));
  AOI211_X1 g475(.A(KEYINPUT48), .B(new_n432_), .C1(new_n674_), .C2(new_n592_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n676_), .B2(new_n677_), .ZN(G1333gat));
  INV_X1    g477(.A(G71gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n668_), .A2(new_n679_), .A3(new_n257_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n663_), .A2(new_n257_), .A3(new_n664_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT49), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(G71gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G71gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT111), .ZN(G1334gat));
  INV_X1    g485(.A(G78gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n668_), .A2(new_n687_), .A3(new_n302_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT50), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n674_), .A2(new_n302_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(G78gat), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT50), .B(new_n687_), .C1(new_n674_), .C2(new_n302_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(G1335gat));
  NOR3_X1   g492(.A1(new_n658_), .A2(new_n612_), .A3(new_n510_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n388_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n667_), .A2(new_n486_), .A3(new_n613_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n414_), .A3(new_n322_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1336gat));
  OAI21_X1  g500(.A(G92gat), .B1(new_n697_), .B2(new_n638_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n415_), .A3(new_n592_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1337gat));
  NAND3_X1  g503(.A1(new_n699_), .A2(new_n257_), .A3(new_n404_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n257_), .B(new_n694_), .C1(new_n624_), .C2(new_n627_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n706_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT112), .B1(new_n706_), .B2(G99gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT51), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT51), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n711_), .B(new_n705_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1338gat));
  INV_X1    g512(.A(KEYINPUT113), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT52), .ZN(new_n715_));
  OAI21_X1  g514(.A(G106gat), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n696_), .B2(new_n302_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n715_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n699_), .A2(new_n405_), .A3(new_n302_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n721_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT53), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n717_), .A2(new_n718_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT53), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(new_n719_), .A4(new_n721_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1339gat));
  NOR2_X1   g526(.A1(new_n592_), .A2(new_n302_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n576_), .A2(new_n388_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT119), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n463_), .A2(new_n454_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n466_), .A2(new_n467_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n474_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT117), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT117), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n468_), .A2(new_n736_), .A3(new_n474_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n470_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n741_));
  AND4_X1   g540(.A1(new_n733_), .A2(new_n732_), .A3(new_n471_), .A4(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n481_), .B1(new_n738_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT56), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n476_), .A2(new_n481_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n481_), .C1(new_n738_), .C2(new_n743_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n745_), .A2(new_n510_), .A3(new_n747_), .A4(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n509_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n490_), .A2(new_n499_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(new_n504_), .A3(new_n502_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n506_), .A2(new_n509_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n482_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n750_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(KEYINPUT57), .A3(new_n566_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n745_), .A2(new_n747_), .A3(new_n754_), .A4(new_n749_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n746_), .B1(new_n744_), .B2(KEYINPUT56), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n761_), .A2(KEYINPUT58), .A3(new_n754_), .A4(new_n749_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n569_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n757_), .A2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n756_), .B2(new_n566_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n731_), .B1(new_n764_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n756_), .A2(new_n566_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n765_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n770_), .A2(KEYINPUT119), .A3(new_n757_), .A4(new_n763_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n536_), .A3(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n484_), .A2(new_n485_), .A3(new_n568_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n659_), .A2(KEYINPUT114), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n534_), .A2(new_n775_), .A3(new_n535_), .A4(new_n511_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n773_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n777_), .B(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n730_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G113gat), .B1(new_n781_), .B2(new_n510_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT120), .Z(new_n783_));
  NOR2_X1   g582(.A1(new_n730_), .A2(KEYINPUT59), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n777_), .B(new_n778_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n764_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n612_), .B1(new_n786_), .B2(new_n770_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n784_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT59), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n781_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n788_), .B(KEYINPUT121), .C1(new_n781_), .C2(new_n789_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(G113gat), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n511_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n783_), .B1(new_n794_), .B2(new_n796_), .ZN(G1340gat));
  OAI21_X1  g596(.A(G120gat), .B1(new_n790_), .B2(new_n658_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n781_), .ZN(new_n799_));
  INV_X1    g598(.A(G120gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n658_), .B2(KEYINPUT60), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(KEYINPUT60), .B2(new_n800_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n799_), .B2(new_n802_), .ZN(G1341gat));
  NAND3_X1  g602(.A1(new_n792_), .A2(new_n612_), .A3(new_n793_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(G127gat), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n536_), .A2(G127gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n799_), .B2(new_n806_), .ZN(G1342gat));
  INV_X1    g606(.A(G134gat), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n568_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n792_), .A2(new_n793_), .A3(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n799_), .B2(new_n566_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT122), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(KEYINPUT122), .A3(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1343gat));
  AOI21_X1  g615(.A(new_n257_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n817_));
  AND4_X1   g616(.A1(new_n322_), .A2(new_n817_), .A3(new_n302_), .A4(new_n638_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n510_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n486_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n612_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT61), .B(G155gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1346gat));
  AOI21_X1  g624(.A(G162gat), .B1(new_n818_), .B2(new_n575_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n569_), .A2(G162gat), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT123), .Z(new_n828_));
  AOI21_X1  g627(.A(new_n826_), .B1(new_n818_), .B2(new_n828_), .ZN(G1347gat));
  NOR2_X1   g628(.A1(new_n785_), .A2(new_n787_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n592_), .A2(new_n398_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT124), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n303_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n218_), .B1(new_n834_), .B2(new_n510_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n835_), .A2(KEYINPUT62), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n510_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n836_), .B(new_n838_), .C1(new_n327_), .C2(new_n837_), .ZN(G1348gat));
  AOI21_X1  g638(.A(G176gat), .B1(new_n834_), .B2(new_n486_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n302_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n832_), .A2(G176gat), .A3(new_n486_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(G1349gat));
  INV_X1    g642(.A(new_n834_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n844_), .A2(new_n231_), .A3(new_n536_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(new_n612_), .A3(new_n832_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G183gat), .B1(new_n846_), .B2(new_n847_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n845_), .B1(new_n848_), .B2(new_n849_), .ZN(G1350gat));
  OAI21_X1  g649(.A(G190gat), .B1(new_n844_), .B2(new_n568_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n834_), .A2(new_n234_), .A3(new_n575_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1351gat));
  NOR2_X1   g652(.A1(new_n638_), .A2(new_n389_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n817_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n510_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n486_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g659(.A1(new_n855_), .A2(new_n536_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  OR3_X1    g662(.A1(new_n861_), .A2(KEYINPUT126), .A3(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT126), .B1(new_n861_), .B2(new_n863_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT63), .B(G211gat), .Z(new_n866_));
  AOI22_X1  g665(.A1(new_n864_), .A2(new_n865_), .B1(new_n861_), .B2(new_n866_), .ZN(G1354gat));
  OR3_X1    g666(.A1(new_n855_), .A2(G218gat), .A3(new_n566_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G218gat), .B1(new_n855_), .B2(new_n568_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1355gat));
endmodule


