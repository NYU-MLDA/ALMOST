//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_;
  XOR2_X1   g000(.A(G1gat), .B(G8gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT70), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT71), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205_));
  INV_X1    g004(.A(G1gat), .ZN(new_n206_));
  INV_X1    g005(.A(G8gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G15gat), .ZN(new_n209_));
  INV_X1    g008(.A(G22gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G15gat), .A2(G22gat), .ZN(new_n212_));
  OAI22_X1  g011(.A1(new_n205_), .A2(new_n208_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n204_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT71), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n203_), .B(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(new_n213_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G29gat), .B(G36gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G43gat), .B(G50gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n222_), .B(KEYINPUT74), .Z(new_n223_));
  XNOR2_X1  g022(.A(new_n219_), .B(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT75), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(KEYINPUT15), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n222_), .B(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n215_), .A2(new_n218_), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT76), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n219_), .A2(new_n223_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n225_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G113gat), .B(G141gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT77), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT78), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G169gat), .B(G197gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n228_), .A2(new_n234_), .A3(new_n240_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(G197gat), .A2(G204gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G197gat), .A2(G204gat), .ZN(new_n247_));
  AND2_X1   g046(.A1(KEYINPUT89), .A2(KEYINPUT21), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G211gat), .B(G218gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n246_), .A2(new_n247_), .ZN(new_n252_));
  OAI22_X1  g051(.A1(new_n249_), .A2(new_n251_), .B1(new_n252_), .B2(KEYINPUT21), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n250_), .B1(new_n252_), .B2(new_n248_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G141gat), .A2(G148gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT2), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n259_), .A2(new_n262_), .A3(new_n263_), .A4(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(KEYINPUT1), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(G155gat), .A3(G162gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n272_), .A3(new_n266_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G141gat), .B(G148gat), .Z(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n256_), .B1(KEYINPUT29), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  NOR2_X1   g078(.A1(new_n276_), .A2(KEYINPUT29), .ZN(new_n280_));
  XOR2_X1   g079(.A(G22gat), .B(G50gat), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n280_), .A2(new_n282_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G228gat), .A2(G233gat), .ZN(new_n287_));
  INV_X1    g086(.A(G78gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G106gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n286_), .A2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n279_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AND3_X1   g096(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT22), .B(G169gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(KEYINPUT83), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT84), .B(G176gat), .ZN(new_n303_));
  INV_X1    g102(.A(G169gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT83), .B1(new_n304_), .B2(KEYINPUT22), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n300_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT85), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n309_), .B(new_n300_), .C1(new_n302_), .C2(new_n306_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT23), .ZN(new_n312_));
  INV_X1    g111(.A(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT79), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT79), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G190gat), .ZN(new_n316_));
  INV_X1    g115(.A(G183gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n308_), .A2(new_n310_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323_));
  NOR4_X1   g122(.A1(new_n298_), .A2(new_n299_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n314_), .A2(new_n316_), .A3(KEYINPUT26), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT26), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G190gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT25), .B(G183gat), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n326_), .A2(KEYINPUT80), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n317_), .A2(KEYINPUT25), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(G183gat), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n328_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT80), .B1(new_n335_), .B2(new_n326_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n325_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT82), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n314_), .A2(new_n316_), .A3(KEYINPUT26), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n328_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n330_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT82), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n325_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n311_), .A2(KEYINPUT23), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(G183gat), .A3(G190gat), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n347_), .A2(new_n349_), .B1(new_n323_), .B2(new_n322_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n321_), .B1(new_n346_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(G71gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(G99gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n351_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G134gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G127gat), .ZN(new_n358_));
  INV_X1    g157(.A(G127gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G134gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G127gat), .B(G134gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT87), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G113gat), .B(G120gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n361_), .A2(new_n362_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n364_), .A2(KEYINPUT87), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n356_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n344_), .B1(new_n343_), .B2(new_n325_), .ZN(new_n373_));
  AOI211_X1 g172(.A(KEYINPUT82), .B(new_n324_), .C1(new_n342_), .C2(new_n330_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n350_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n320_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(new_n355_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n367_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n366_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n372_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G15gat), .B(G43gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT86), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT30), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT31), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n381_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n372_), .A2(new_n380_), .A3(new_n385_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n265_), .A2(new_n268_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n276_), .A2(new_n371_), .A3(new_n367_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(KEYINPUT4), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n276_), .A2(new_n371_), .A3(new_n395_), .A4(new_n367_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n392_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n390_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n399_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(new_n398_), .A3(new_n404_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n387_), .A2(new_n388_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT100), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n375_), .A2(new_n320_), .A3(new_n256_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n313_), .A2(KEYINPUT26), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n329_), .A2(new_n328_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT90), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(KEYINPUT24), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(G169gat), .B2(G176gat), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n416_), .B2(KEYINPUT24), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n415_), .B(new_n350_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n301_), .A2(new_n303_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n347_), .A2(new_n349_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(G183gat), .A2(G190gat), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n422_), .B(new_n300_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n255_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT91), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n255_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n413_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n412_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT19), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT92), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n256_), .B1(new_n375_), .B2(new_n320_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n426_), .A2(new_n255_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n434_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(KEYINPUT20), .A3(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n436_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n442_), .B(KEYINPUT92), .C1(new_n351_), .C2(new_n256_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n435_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G8gat), .B(G36gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT18), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G64gat), .B(G92gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n435_), .A2(new_n441_), .A3(new_n443_), .A4(new_n448_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT27), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n376_), .A2(new_n255_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT97), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n255_), .B1(new_n426_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n421_), .A2(new_n425_), .A3(KEYINPUT97), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n413_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n439_), .B1(new_n453_), .B2(new_n457_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n412_), .A2(new_n439_), .A3(new_n431_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n449_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(KEYINPUT27), .A3(new_n451_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n411_), .B1(new_n452_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT27), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n440_), .B1(new_n376_), .B2(new_n255_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(KEYINPUT92), .A2(new_n465_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n448_), .B1(new_n466_), .B2(new_n441_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n451_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n464_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(KEYINPUT100), .A3(new_n461_), .ZN(new_n470_));
  AOI211_X1 g269(.A(new_n297_), .B(new_n410_), .C1(new_n463_), .C2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n387_), .A2(new_n388_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n296_), .A2(new_n408_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n469_), .A2(new_n461_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475_));
  OR3_X1    g274(.A1(new_n407_), .A2(KEYINPUT94), .A3(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT94), .B1(new_n407_), .B2(new_n475_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT95), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT33), .B1(new_n407_), .B2(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n397_), .A2(KEYINPUT95), .A3(new_n398_), .A4(new_n404_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n392_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n390_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n405_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT96), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n482_), .A2(new_n486_), .A3(new_n405_), .A4(new_n483_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n480_), .A2(new_n481_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n450_), .A2(new_n451_), .A3(new_n478_), .A4(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n448_), .A2(KEYINPUT32), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n435_), .A2(new_n441_), .A3(new_n443_), .A4(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n458_), .A2(new_n459_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n491_), .B(new_n408_), .C1(new_n492_), .C2(new_n490_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n297_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n474_), .B1(new_n494_), .B2(KEYINPUT98), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT98), .ZN(new_n496_));
  AOI211_X1 g295(.A(new_n496_), .B(new_n297_), .C1(new_n489_), .C2(new_n493_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n472_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n471_), .B1(new_n498_), .B2(KEYINPUT99), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT99), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n500_), .B(new_n472_), .C1(new_n495_), .C2(new_n497_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n245_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G85gat), .B(G92gat), .Z(new_n503_));
  NOR2_X1   g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT7), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n503_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT8), .B1(new_n503_), .B2(KEYINPUT65), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n503_), .A2(KEYINPUT9), .ZN(new_n513_));
  INV_X1    g312(.A(G85gat), .ZN(new_n514_));
  INV_X1    g313(.A(G92gat), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT9), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT10), .B(G99gat), .Z(new_n518_));
  AND3_X1   g317(.A1(new_n518_), .A2(KEYINPUT64), .A3(new_n290_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT64), .B1(new_n518_), .B2(new_n290_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n513_), .B(new_n517_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n510_), .A2(new_n511_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n512_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n526_));
  XOR2_X1   g325(.A(G71gat), .B(G78gat), .Z(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n526_), .A2(new_n527_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n523_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT12), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT12), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n523_), .A2(new_n533_), .A3(new_n529_), .A4(new_n528_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G230gat), .A2(G233gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n536_), .B2(new_n531_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT5), .ZN(new_n540_));
  XOR2_X1   g339(.A(G176gat), .B(G204gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(KEYINPUT66), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n538_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n546_), .A2(KEYINPUT13), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(KEYINPUT13), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n523_), .A2(new_n230_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT67), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n512_), .A2(new_n222_), .A3(new_n521_), .A4(new_n522_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n555_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n559_));
  OAI22_X1  g358(.A1(new_n558_), .A2(new_n559_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n553_), .A2(new_n550_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n557_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n560_), .A2(new_n563_), .A3(KEYINPUT36), .A4(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT69), .B1(new_n560_), .B2(new_n563_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(KEYINPUT36), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  AOI211_X1 g370(.A(KEYINPUT69), .B(new_n571_), .C1(new_n560_), .C2(new_n563_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n567_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT37), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n576_), .B(new_n567_), .C1(new_n570_), .C2(new_n572_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n530_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n219_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585_));
  XOR2_X1   g384(.A(G127gat), .B(G155gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n584_), .A2(new_n585_), .A3(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT73), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n590_), .B(KEYINPUT17), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n584_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n580_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n502_), .A2(new_n549_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT101), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(new_n206_), .A3(new_n408_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n573_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n549_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n603_), .A2(new_n245_), .A3(new_n595_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n206_), .B1(new_n605_), .B2(new_n408_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n600_), .B2(new_n599_), .ZN(G1324gat));
  INV_X1    g407(.A(new_n463_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n470_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n207_), .B1(new_n605_), .B2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT39), .Z(new_n613_));
  NAND3_X1  g412(.A1(new_n598_), .A2(new_n207_), .A3(new_n611_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g415(.A(new_n472_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n209_), .B1(new_n605_), .B2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT41), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n598_), .A2(new_n209_), .A3(new_n617_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1326gat));
  AOI21_X1  g420(.A(new_n210_), .B1(new_n605_), .B2(new_n297_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT42), .Z(new_n623_));
  NAND3_X1  g422(.A1(new_n598_), .A2(new_n210_), .A3(new_n297_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1327gat));
  NAND2_X1  g424(.A1(new_n498_), .A2(KEYINPUT99), .ZN(new_n626_));
  INV_X1    g425(.A(new_n471_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n501_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n595_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n573_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AND4_X1   g430(.A1(new_n628_), .A2(new_n244_), .A3(new_n549_), .A4(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(G29gat), .B1(new_n632_), .B2(new_n408_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n574_), .A2(KEYINPUT103), .A3(new_n577_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT103), .B1(new_n574_), .B2(new_n577_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n628_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT43), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n628_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n641_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT104), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n639_), .A2(new_n645_), .A3(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n549_), .A2(new_n244_), .A3(new_n595_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT102), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT44), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n408_), .A2(G29gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n633_), .B1(new_n652_), .B2(new_n653_), .ZN(G1328gat));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n611_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G36gat), .ZN(new_n656_));
  INV_X1    g455(.A(G36gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n632_), .A2(new_n657_), .A3(new_n611_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n656_), .A2(new_n668_), .A3(KEYINPUT46), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n657_), .B1(new_n652_), .B2(new_n611_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n667_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n672_), .ZN(G1329gat));
  NAND3_X1  g472(.A1(new_n652_), .A2(G43gat), .A3(new_n617_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n632_), .A2(new_n617_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(G43gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT47), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT47), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n674_), .A2(new_n679_), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1330gat));
  INV_X1    g480(.A(G50gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n632_), .A2(new_n682_), .A3(new_n297_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n652_), .A2(new_n297_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(KEYINPUT107), .ZN(new_n685_));
  OAI21_X1  g484(.A(G50gat), .B1(new_n684_), .B2(KEYINPUT107), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(G1331gat));
  NOR2_X1   g486(.A1(new_n549_), .A2(new_n244_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n628_), .A2(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(new_n596_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n408_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT108), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n602_), .A2(new_n629_), .A3(new_n688_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT109), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n408_), .A2(G57gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n692_), .B1(new_n694_), .B2(new_n695_), .ZN(G1332gat));
  INV_X1    g495(.A(G64gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n694_), .B2(new_n611_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT48), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n690_), .A2(new_n697_), .A3(new_n611_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1333gat));
  AOI21_X1  g500(.A(new_n353_), .B1(new_n694_), .B2(new_n617_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT49), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n690_), .A2(new_n353_), .A3(new_n617_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1334gat));
  AOI21_X1  g504(.A(new_n288_), .B1(new_n694_), .B2(new_n297_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT50), .Z(new_n707_));
  NAND3_X1  g506(.A1(new_n690_), .A2(new_n288_), .A3(new_n297_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1335gat));
  NOR3_X1   g508(.A1(new_n549_), .A2(new_n244_), .A3(new_n629_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n648_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n514_), .B1(new_n711_), .B2(new_n408_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n689_), .A2(new_n631_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n713_), .A2(new_n514_), .A3(new_n408_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1336gat));
  NAND3_X1  g514(.A1(new_n713_), .A2(new_n515_), .A3(new_n611_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n711_), .A2(new_n611_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n718_), .B2(new_n515_), .ZN(G1337gat));
  NAND3_X1  g518(.A1(new_n713_), .A2(new_n617_), .A3(new_n518_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n711_), .A2(new_n617_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G99gat), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725_));
  AOI22_X1  g524(.A1(new_n722_), .A2(new_n724_), .B1(KEYINPUT111), .B2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(KEYINPUT111), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1338gat));
  NAND3_X1  g527(.A1(new_n713_), .A2(new_n290_), .A3(new_n297_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n648_), .A2(KEYINPUT112), .A3(new_n297_), .A4(new_n710_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(G106gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n636_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n733_));
  OAI22_X1  g532(.A1(new_n640_), .A2(new_n733_), .B1(new_n646_), .B2(KEYINPUT104), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n643_), .A2(new_n644_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n297_), .B(new_n710_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n730_), .B1(new_n732_), .B2(new_n738_), .ZN(new_n739_));
  AND4_X1   g538(.A1(new_n730_), .A2(new_n738_), .A3(G106gat), .A4(new_n731_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n729_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n729_), .B(new_n742_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1339gat));
  NAND2_X1  g545(.A1(new_n244_), .A2(new_n543_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n535_), .A2(new_n536_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT55), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT115), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n535_), .A2(new_n536_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n748_), .B2(new_n752_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n750_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(KEYINPUT56), .A3(new_n544_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n750_), .A2(new_n753_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n544_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n747_), .B1(new_n755_), .B2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n232_), .A2(new_n233_), .A3(new_n226_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n240_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT116), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n546_), .A3(new_n243_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n766_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT57), .B(new_n630_), .C1(new_n760_), .C2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n764_), .A2(new_n243_), .A3(new_n543_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n755_), .B2(new_n759_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n774_), .A2(KEYINPUT58), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n579_), .B1(new_n774_), .B2(KEYINPUT58), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n630_), .B1(new_n760_), .B2(new_n769_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n595_), .B1(new_n772_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n596_), .A2(new_n549_), .ZN(new_n783_));
  OR3_X1    g582(.A1(new_n783_), .A2(KEYINPUT54), .A3(new_n244_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT54), .B1(new_n783_), .B2(new_n244_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n782_), .A2(new_n786_), .ZN(new_n787_));
  NOR4_X1   g586(.A1(new_n611_), .A2(new_n472_), .A3(new_n297_), .A4(new_n409_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(G113gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n244_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT59), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n544_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n757_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n767_), .B(new_n768_), .C1(new_n796_), .C2(new_n747_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n797_), .A2(new_n771_), .A3(KEYINPUT57), .A4(new_n630_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n770_), .A2(KEYINPUT118), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n775_), .A2(new_n776_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n629_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n786_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n793_), .B(new_n788_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n792_), .A2(KEYINPUT59), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n805_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n787_), .A2(new_n793_), .A3(new_n788_), .A4(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n245_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n791_), .B1(new_n809_), .B2(new_n790_), .ZN(G1340gat));
  INV_X1    g609(.A(G120gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n549_), .B2(KEYINPUT60), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n789_), .B(new_n812_), .C1(KEYINPUT60), .C2(new_n811_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n549_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n811_), .ZN(G1341gat));
  NAND2_X1  g614(.A1(new_n629_), .A2(G127gat), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n629_), .B(new_n788_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n359_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n818_), .B2(new_n359_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n817_), .A2(new_n820_), .A3(new_n821_), .ZN(G1342gat));
  NAND3_X1  g621(.A1(new_n789_), .A2(new_n357_), .A3(new_n573_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n579_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n357_), .ZN(G1343gat));
  NOR2_X1   g624(.A1(new_n802_), .A2(new_n803_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n611_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n827_), .A2(new_n472_), .A3(new_n297_), .A4(new_n408_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT121), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n826_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n244_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n603_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(KEYINPUT122), .B(G148gat), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(G1345gat));
  NAND2_X1  g635(.A1(new_n831_), .A2(new_n629_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1346gat));
  NAND3_X1  g638(.A1(new_n787_), .A2(new_n573_), .A3(new_n829_), .ZN(new_n840_));
  INV_X1    g639(.A(G162gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT123), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n840_), .A2(new_n844_), .A3(new_n841_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n636_), .A2(new_n841_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n843_), .A2(new_n845_), .B1(new_n831_), .B2(new_n846_), .ZN(G1347gat));
  INV_X1    g646(.A(KEYINPUT62), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n410_), .A2(new_n297_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n611_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n787_), .A2(new_n244_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n848_), .B1(new_n853_), .B2(new_n304_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n301_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(G1348gat));
  NAND3_X1  g656(.A1(new_n787_), .A2(new_n603_), .A3(new_n851_), .ZN(new_n858_));
  INV_X1    g657(.A(G176gat), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n303_), .B2(new_n858_), .ZN(G1349gat));
  NAND3_X1  g660(.A1(new_n787_), .A2(new_n629_), .A3(new_n851_), .ZN(new_n862_));
  OR3_X1    g661(.A1(new_n862_), .A2(KEYINPUT124), .A3(new_n329_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT124), .B1(new_n862_), .B2(new_n329_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n826_), .A2(new_n850_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G183gat), .B1(new_n865_), .B2(new_n629_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n863_), .B1(new_n864_), .B2(new_n866_), .ZN(G1350gat));
  NAND4_X1  g666(.A1(new_n865_), .A2(new_n328_), .A3(new_n414_), .A4(new_n573_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n787_), .A2(new_n580_), .A3(new_n851_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n869_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT125), .B1(new_n869_), .B2(G190gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n868_), .B1(new_n870_), .B2(new_n871_), .ZN(G1351gat));
  INV_X1    g671(.A(new_n473_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n827_), .A2(new_n617_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n826_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n244_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n603_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g679(.A(new_n595_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n874_), .B(new_n881_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n882_), .A2(KEYINPUT126), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(KEYINPUT126), .ZN(new_n884_));
  OAI22_X1  g683(.A1(new_n883_), .A2(new_n884_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n882_), .A2(KEYINPUT126), .ZN(new_n886_));
  NOR2_X1   g685(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n882_), .A2(KEYINPUT126), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n885_), .A2(new_n889_), .ZN(G1354gat));
  OAI211_X1 g689(.A(new_n573_), .B(new_n874_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(KEYINPUT127), .ZN(new_n893_));
  AOI21_X1  g692(.A(G218gat), .B1(new_n892_), .B2(KEYINPUT127), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n580_), .A2(G218gat), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n894_), .B1(new_n876_), .B2(new_n895_), .ZN(G1355gat));
endmodule


