//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n918_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT72), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(G43gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT71), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G50gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n210_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G50gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT6), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  OR3_X1    g021(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G85gat), .B(G92gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n225_), .A2(new_n226_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT65), .B(KEYINPUT8), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n231_), .A2(KEYINPUT67), .B1(KEYINPUT8), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(KEYINPUT67), .B2(new_n231_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(new_n225_), .B2(KEYINPUT9), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n237_), .A2(KEYINPUT64), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(KEYINPUT64), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT10), .B(G99gat), .Z(new_n240_));
  INV_X1    g039(.A(G106gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n238_), .A2(new_n221_), .A3(new_n239_), .A4(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n234_), .A2(new_n243_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n219_), .A2(new_n244_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n212_), .A2(new_n216_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n208_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n206_), .A2(new_n207_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n245_), .A2(new_n207_), .A3(new_n248_), .A4(new_n206_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G134gat), .B(G162gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT73), .ZN(new_n255_));
  INV_X1    g054(.A(G190gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G218gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT36), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT74), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n253_), .A2(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n258_), .A2(new_n259_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n251_), .A2(new_n252_), .A3(new_n260_), .A4(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n261_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT37), .B1(new_n267_), .B2(KEYINPUT75), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n266_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT76), .B(G1gat), .ZN(new_n270_));
  INV_X1    g069(.A(G8gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT14), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G15gat), .B(G22gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G1gat), .B(G8gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n274_), .B(KEYINPUT77), .ZN(new_n279_));
  INV_X1    g078(.A(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G231gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G71gat), .B(G78gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G64gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(KEYINPUT11), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n284_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G127gat), .B(G155gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT16), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(G183gat), .ZN(new_n294_));
  INV_X1    g093(.A(G211gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT17), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n296_), .A2(new_n297_), .ZN(new_n299_));
  OR3_X1    g098(.A1(new_n291_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n291_), .A2(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n269_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT78), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G225gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n307_));
  AND2_X1   g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NOR3_X1   g108(.A1(new_n308_), .A2(new_n309_), .A3(KEYINPUT1), .ZN(new_n310_));
  INV_X1    g109(.A(G141gat), .ZN(new_n311_));
  INV_X1    g110(.A(G148gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n307_), .B1(new_n310_), .B2(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n315_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n321_), .A2(new_n324_), .A3(KEYINPUT88), .A4(new_n314_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n311_), .A2(new_n312_), .A3(KEYINPUT89), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT3), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n315_), .A2(KEYINPUT90), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT2), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n323_), .A2(KEYINPUT89), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n315_), .A2(KEYINPUT90), .A3(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n328_), .A2(new_n330_), .A3(new_n332_), .A4(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n308_), .A2(new_n309_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n326_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G127gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(G134gat), .ZN(new_n340_));
  INV_X1    g139(.A(G134gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(G127gat), .ZN(new_n342_));
  INV_X1    g141(.A(G113gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(G120gat), .ZN(new_n344_));
  INV_X1    g143(.A(G120gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n345_), .A2(G113gat), .ZN(new_n346_));
  OAI22_X1  g145(.A1(new_n340_), .A2(new_n342_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G127gat), .B(G134gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT87), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  OR3_X1    g151(.A1(new_n348_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n338_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n306_), .B1(new_n355_), .B2(KEYINPUT4), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT96), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n347_), .A2(new_n350_), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n317_), .A2(new_n325_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n355_), .A2(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n338_), .A2(KEYINPUT96), .A3(new_n354_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n360_), .A2(KEYINPUT97), .A3(KEYINPUT4), .A4(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n352_), .A2(new_n353_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n357_), .B1(new_n363_), .B2(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(new_n358_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n361_), .A4(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT97), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n356_), .B1(new_n362_), .B2(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n364_), .A2(new_n361_), .A3(new_n365_), .A4(new_n305_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT98), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G1gat), .B(G29gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT0), .ZN(new_n373_));
  INV_X1    g172(.A(G57gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G85gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n369_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n356_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n366_), .A2(new_n367_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n366_), .A2(new_n367_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT98), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n370_), .B(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n379_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n378_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G15gat), .B(G43gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT85), .ZN(new_n390_));
  XOR2_X1   g189(.A(G71gat), .B(G99gat), .Z(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n392_), .B(new_n393_), .Z(new_n394_));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT23), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(G169gat), .A2(G176gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G169gat), .A2(G176gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(KEYINPUT24), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT24), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT25), .B(G183gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT26), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G190gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n256_), .A2(KEYINPUT26), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n410_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT83), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n413_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT82), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n411_), .A4(new_n407_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n406_), .B1(new_n415_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G183gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n256_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n397_), .A2(new_n422_), .A3(new_n398_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n402_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT22), .B(G169gat), .ZN(new_n427_));
  INV_X1    g226(.A(G176gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n397_), .A2(new_n422_), .A3(KEYINPUT84), .A4(new_n398_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n425_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n420_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT30), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n394_), .B1(new_n434_), .B2(KEYINPUT86), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(KEYINPUT86), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n354_), .B(KEYINPUT31), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n438_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G211gat), .B(G218gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT21), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT21), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n295_), .A2(G218gat), .ZN(new_n445_));
  INV_X1    g244(.A(G218gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(G211gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n444_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G197gat), .B(G204gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n443_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n442_), .A2(new_n449_), .A3(KEYINPUT21), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(new_n338_), .B2(KEYINPUT29), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G228gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G78gat), .B(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n457_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n338_), .A2(KEYINPUT29), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G22gat), .B(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT28), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n463_), .B(new_n465_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n460_), .A2(new_n462_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n460_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n441_), .A2(new_n470_), .A3(new_n387_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n453_), .B1(new_n420_), .B2(new_n432_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n399_), .A2(new_n405_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n421_), .A2(KEYINPUT25), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT25), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(G183gat), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n409_), .A2(new_n413_), .A3(new_n475_), .A4(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n478_), .A2(new_n403_), .A3(KEYINPUT92), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT92), .B1(new_n478_), .B2(new_n403_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n474_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n402_), .B(KEYINPUT93), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n423_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n427_), .B(KEYINPUT94), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(G176gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n454_), .A2(new_n481_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n472_), .A2(new_n487_), .A3(KEYINPUT20), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G226gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT19), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n481_), .A2(new_n486_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n453_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n490_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n415_), .A2(new_n419_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n431_), .B(new_n454_), .C1(new_n496_), .C2(new_n406_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G8gat), .B(G36gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G64gat), .B(G92gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n499_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n478_), .A2(new_n403_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT92), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n478_), .A2(new_n403_), .A3(KEYINPUT92), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n473_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n427_), .B(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n483_), .B1(new_n513_), .B2(new_n428_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n453_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n497_), .A2(new_n515_), .A3(KEYINPUT20), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n490_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n472_), .A2(new_n487_), .A3(KEYINPUT20), .A4(new_n495_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n504_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n506_), .A2(KEYINPUT27), .A3(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT101), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n495_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n518_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n505_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n519_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT27), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n520_), .A2(KEYINPUT101), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n521_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n471_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n360_), .A2(new_n361_), .A3(new_n306_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n377_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n362_), .A2(new_n368_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n355_), .A2(KEYINPUT4), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(new_n306_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n532_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(new_n525_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n378_), .B2(KEYINPUT33), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n383_), .A2(new_n379_), .A3(new_n385_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT33), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n504_), .A2(KEYINPUT32), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n499_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n517_), .A2(new_n518_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n543_), .B1(new_n544_), .B2(new_n542_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n377_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n539_), .B2(new_n546_), .ZN(new_n547_));
  OAI22_X1  g346(.A1(new_n538_), .A2(new_n541_), .B1(new_n547_), .B2(KEYINPUT99), .ZN(new_n548_));
  INV_X1    g347(.A(new_n545_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n549_), .B1(new_n378_), .B2(new_n386_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT99), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n470_), .B1(new_n548_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT100), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n551_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(KEYINPUT99), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n378_), .A2(KEYINPUT33), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n539_), .A2(new_n540_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(new_n537_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n557_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(KEYINPUT100), .A3(new_n470_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n470_), .A2(new_n388_), .A3(new_n529_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n555_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n441_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n530_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n244_), .A2(new_n289_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n289_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n234_), .B2(new_n243_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(KEYINPUT68), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n568_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT68), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT12), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n572_), .B1(new_n570_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(new_n574_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n574_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n584_));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n580_), .A2(new_n582_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT13), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(KEYINPUT13), .A3(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n247_), .A2(new_n282_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n278_), .A2(new_n281_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n217_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n599_), .A3(KEYINPUT79), .ZN(new_n600_));
  OR3_X1    g399(.A1(new_n247_), .A2(KEYINPUT79), .A3(new_n282_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n600_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT80), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(KEYINPUT80), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n219_), .A2(new_n598_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n602_), .A3(new_n597_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(G169gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(G197gat), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n609_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n613_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT81), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n567_), .A2(new_n596_), .A3(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n304_), .A2(new_n270_), .A3(new_n388_), .A4(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n530_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n561_), .A2(KEYINPUT100), .A3(new_n470_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT100), .B1(new_n561_), .B2(new_n470_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n563_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n628_), .B2(new_n441_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n596_), .A2(new_n302_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n629_), .A2(new_n266_), .A3(new_n619_), .A4(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n387_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n622_), .A2(new_n623_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n624_), .A2(new_n632_), .A3(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(new_n529_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G8gat), .B1(new_n631_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT102), .B(G8gat), .C1(new_n631_), .C2(new_n635_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(KEYINPUT39), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n636_), .A2(new_n637_), .A3(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n304_), .A2(new_n271_), .A3(new_n529_), .A4(new_n621_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT103), .B1(new_n641_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n640_), .A2(new_n647_), .A3(new_n644_), .A4(new_n643_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n646_), .A2(new_n648_), .A3(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n631_), .B2(new_n566_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT41), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n304_), .A2(new_n621_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n656_), .A2(G15gat), .A3(new_n566_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1326gat));
  XOR2_X1   g457(.A(new_n469_), .B(KEYINPUT104), .Z(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G22gat), .B1(new_n631_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n660_), .A2(G22gat), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT106), .Z(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n656_), .B2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n266_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n302_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n621_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n388_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n619_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n302_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n596_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n629_), .B2(new_n269_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n266_), .B(KEYINPUT37), .C1(KEYINPUT75), .C2(new_n267_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n268_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n567_), .A2(KEYINPUT43), .A3(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT44), .B(new_n675_), .C1(new_n677_), .C2(new_n681_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(G29gat), .A3(new_n388_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n675_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n672_), .B1(new_n683_), .B2(new_n686_), .ZN(G1328gat));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688_));
  INV_X1    g487(.A(G36gat), .ZN(new_n689_));
  INV_X1    g488(.A(new_n675_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n567_), .B2(new_n680_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n627_), .A2(new_n563_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n441_), .B1(new_n692_), .B2(new_n562_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n269_), .B(new_n676_), .C1(new_n693_), .C2(new_n530_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n690_), .B1(new_n691_), .B2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n635_), .B1(new_n695_), .B2(KEYINPUT44), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n689_), .B1(new_n696_), .B2(new_n686_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n635_), .A2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT45), .B1(new_n670_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n621_), .A2(new_n701_), .A3(new_n669_), .A4(new_n698_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n688_), .B1(new_n697_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n682_), .A2(new_n529_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n695_), .A2(KEYINPUT44), .ZN(new_n706_));
  OAI21_X1  g505(.A(G36gat), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n700_), .A2(new_n702_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(KEYINPUT107), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n704_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n704_), .A2(new_n709_), .A3(KEYINPUT108), .A4(new_n710_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n707_), .A2(KEYINPUT46), .A3(new_n708_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(new_n714_), .A3(new_n715_), .ZN(G1329gat));
  INV_X1    g515(.A(G43gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(new_n670_), .B2(new_n566_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n682_), .A2(G43gat), .A3(new_n441_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n706_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT109), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n720_), .A2(KEYINPUT109), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n720_), .A2(KEYINPUT109), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(KEYINPUT47), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n671_), .B2(new_n659_), .ZN(new_n728_));
  AOI211_X1 g527(.A(new_n215_), .B(new_n470_), .C1(new_n695_), .C2(KEYINPUT44), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n686_), .ZN(G1331gat));
  NAND2_X1  g529(.A1(new_n596_), .A2(new_n673_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n304_), .A2(new_n629_), .A3(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT110), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n374_), .A3(new_n388_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n596_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(new_n302_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n629_), .A2(new_n266_), .A3(new_n620_), .A4(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G57gat), .B1(new_n738_), .B2(new_n387_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n735_), .A2(new_n739_), .ZN(G1332gat));
  OAI21_X1  g539(.A(G64gat), .B1(new_n738_), .B2(new_n635_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT111), .Z(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT48), .ZN(new_n743_));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n734_), .A2(new_n744_), .A3(new_n529_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n738_), .B2(new_n566_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT112), .Z(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT49), .ZN(new_n749_));
  INV_X1    g548(.A(G71gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n734_), .A2(new_n750_), .A3(new_n441_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1334gat));
  INV_X1    g551(.A(G78gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n734_), .A2(new_n753_), .A3(new_n659_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G78gat), .B1(new_n738_), .B2(new_n660_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT50), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n732_), .A2(new_n302_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n691_), .B2(new_n694_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n376_), .B1(new_n759_), .B2(new_n388_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n567_), .A2(new_n668_), .A3(new_n731_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n761_), .A2(new_n376_), .A3(new_n388_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1336gat));
  AOI21_X1  g562(.A(G92gat), .B1(new_n761_), .B2(new_n529_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT113), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n759_), .A2(G92gat), .A3(new_n529_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1337gat));
  NAND3_X1  g566(.A1(new_n761_), .A2(new_n240_), .A3(new_n441_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT115), .Z(new_n769_));
  INV_X1    g568(.A(G99gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n759_), .B2(new_n441_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(KEYINPUT114), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT114), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT51), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n775_), .A2(KEYINPUT51), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n774_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n774_), .B2(new_n777_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1338gat));
  AOI21_X1  g579(.A(new_n241_), .B1(new_n759_), .B2(new_n469_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n781_), .A2(KEYINPUT52), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(KEYINPUT52), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n761_), .A2(new_n241_), .A3(new_n469_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT117), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n783_), .A3(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g586(.A1(new_n529_), .A2(new_n387_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n441_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n602_), .B1(new_n247_), .B2(new_n282_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n613_), .B1(new_n608_), .B2(new_n792_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n617_), .A2(new_n613_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n592_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n570_), .A2(new_n572_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n289_), .B2(new_n244_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n797_), .A2(new_n581_), .A3(new_n578_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n581_), .B1(new_n797_), .B2(new_n578_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(KEYINPUT55), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(KEYINPUT55), .B2(new_n799_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n588_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  INV_X1    g604(.A(new_n591_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n807_));
  OAI22_X1  g606(.A1(new_n804_), .A2(new_n805_), .B1(new_n807_), .B2(KEYINPUT118), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n619_), .A2(KEYINPUT118), .A3(new_n591_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n799_), .A2(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n580_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n798_), .A2(new_n799_), .A3(KEYINPUT55), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n590_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n805_), .B1(new_n813_), .B2(KEYINPUT119), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n809_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n795_), .B1(new_n808_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n266_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n802_), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n819_));
  NAND2_X1  g618(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n820_));
  OR2_X1    g619(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n813_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n794_), .A2(new_n823_), .A3(new_n591_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n794_), .B2(new_n591_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n819_), .B(new_n822_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n680_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n819_), .A2(new_n822_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n828_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n830_), .B(new_n831_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n817_), .A2(new_n818_), .B1(new_n829_), .B2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n816_), .A2(KEYINPUT57), .A3(new_n266_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n674_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n620_), .A2(new_n680_), .A3(new_n630_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n470_), .B(new_n790_), .C1(new_n835_), .C2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n343_), .A3(new_n619_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  INV_X1    g641(.A(new_n795_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n619_), .A2(new_n591_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n811_), .A2(new_n812_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT119), .B1(new_n846_), .B2(new_n588_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n844_), .A2(new_n845_), .B1(new_n847_), .B2(KEYINPUT56), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n804_), .A2(new_n805_), .B1(new_n807_), .B2(KEYINPUT118), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n843_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n818_), .B1(new_n850_), .B2(new_n667_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n829_), .A2(new_n832_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n834_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n838_), .B1(new_n853_), .B2(new_n302_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n469_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n842_), .B1(new_n855_), .B2(new_n790_), .ZN(new_n856_));
  NOR4_X1   g655(.A1(new_n854_), .A2(KEYINPUT59), .A3(new_n469_), .A4(new_n789_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n856_), .A2(new_n620_), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n841_), .B1(new_n858_), .B2(new_n343_), .ZN(G1340gat));
  NAND2_X1  g658(.A1(new_n839_), .A2(KEYINPUT59), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n853_), .A2(new_n302_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n838_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n863_), .A2(new_n842_), .A3(new_n470_), .A4(new_n790_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n736_), .B2(G120gat), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n863_), .A2(new_n470_), .A3(new_n790_), .A4(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n860_), .A2(new_n596_), .A3(new_n864_), .A4(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G120gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n840_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1341gat));
  NAND3_X1  g670(.A1(new_n840_), .A2(new_n339_), .A3(new_n674_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n856_), .A2(new_n302_), .A3(new_n857_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n339_), .ZN(G1342gat));
  NAND3_X1  g673(.A1(new_n840_), .A2(new_n341_), .A3(new_n667_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n856_), .A2(new_n680_), .A3(new_n857_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n341_), .ZN(G1343gat));
  NOR2_X1   g676(.A1(new_n441_), .A2(new_n470_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n854_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(new_n619_), .A3(new_n788_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n596_), .A3(new_n788_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT123), .B(G148gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1345gat));
  NAND3_X1  g684(.A1(new_n880_), .A2(new_n674_), .A3(new_n788_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G155gat), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT124), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n886_), .B(new_n888_), .ZN(G1346gat));
  NAND2_X1  g688(.A1(new_n880_), .A2(new_n788_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G162gat), .B1(new_n890_), .B2(new_n680_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n266_), .A2(G162gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n890_), .B2(new_n892_), .ZN(G1347gat));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n635_), .A2(new_n388_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n441_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n659_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n863_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n673_), .ZN(new_n899_));
  INV_X1    g698(.A(G169gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n894_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  OAI211_X1 g700(.A(KEYINPUT62), .B(G169gat), .C1(new_n898_), .C2(new_n673_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n513_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(G1348gat));
  INV_X1    g703(.A(new_n898_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G176gat), .B1(new_n905_), .B2(new_n596_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n736_), .A2(new_n428_), .A3(new_n896_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n855_), .B2(new_n907_), .ZN(G1349gat));
  NOR3_X1   g707(.A1(new_n898_), .A2(new_n302_), .A3(new_n407_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n896_), .A2(new_n302_), .ZN(new_n910_));
  AOI21_X1  g709(.A(KEYINPUT125), .B1(new_n855_), .B2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(G183gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n855_), .A2(KEYINPUT125), .A3(new_n910_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n909_), .B1(new_n912_), .B2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n898_), .B2(new_n680_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n266_), .A2(new_n416_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n898_), .B2(new_n916_), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n880_), .A2(new_n619_), .A3(new_n895_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g718(.A1(new_n880_), .A2(new_n596_), .A3(new_n895_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n920_), .B(new_n921_), .Z(G1353gat));
  INV_X1    g721(.A(new_n895_), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n854_), .A2(new_n302_), .A3(new_n879_), .A4(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  AND2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n924_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n924_), .B2(new_n925_), .ZN(G1354gat));
  NOR2_X1   g727(.A1(new_n266_), .A2(G218gat), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n880_), .A2(new_n895_), .A3(new_n929_), .ZN(new_n930_));
  NOR4_X1   g729(.A1(new_n854_), .A2(new_n680_), .A3(new_n879_), .A4(new_n923_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n446_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n930_), .B(KEYINPUT127), .C1(new_n446_), .C2(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1355gat));
endmodule


