//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(KEYINPUT64), .A2(KEYINPUT8), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT64), .A2(KEYINPUT8), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n205_), .B(new_n206_), .C1(new_n207_), .C2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT7), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n209_), .B1(new_n215_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n205_), .A2(new_n206_), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n217_), .A2(new_n219_), .A3(KEYINPUT65), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(new_n214_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n223_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n222_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n223_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT9), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT10), .B(G99gat), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n212_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n233_), .A2(new_n235_), .A3(new_n220_), .A4(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n202_), .B1(new_n231_), .B2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n217_), .A2(new_n219_), .A3(KEYINPUT65), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n228_), .A2(new_n239_), .A3(new_n215_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n230_), .B1(new_n240_), .B2(new_n232_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n202_), .B(new_n237_), .C1(new_n241_), .C2(new_n221_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G57gat), .B(G64gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G71gat), .B(G78gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n244_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n252_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(G230gat), .A2(G233gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT67), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(new_n260_), .A3(new_n257_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n231_), .A2(new_n237_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(KEYINPUT12), .A3(new_n254_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n257_), .B1(new_n244_), .B2(new_n252_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT68), .B1(new_n255_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n239_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT65), .B1(new_n217_), .B2(new_n219_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n232_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n221_), .B1(new_n270_), .B2(KEYINPUT8), .ZN(new_n271_));
  INV_X1    g070(.A(new_n237_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT66), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n252_), .B1(new_n273_), .B2(new_n242_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n274_), .A2(new_n275_), .A3(KEYINPUT12), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n264_), .B(new_n265_), .C1(new_n267_), .C2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G120gat), .B(G148gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT5), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G176gat), .B(G204gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n262_), .A2(KEYINPUT69), .A3(new_n277_), .A4(new_n282_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n259_), .A2(new_n277_), .A3(new_n261_), .A4(new_n282_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n262_), .A2(new_n277_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n281_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT13), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(KEYINPUT70), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT13), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(KEYINPUT13), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n287_), .A2(new_n289_), .A3(new_n294_), .A4(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT71), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n292_), .A2(new_n300_), .A3(new_n297_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT84), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(KEYINPUT23), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n307_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n308_), .B(new_n309_), .C1(G183gat), .C2(G190gat), .ZN(new_n310_));
  INV_X1    g109(.A(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(G176gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT22), .B(G169gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n313_), .B1(new_n314_), .B2(new_n312_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n304_), .B(new_n306_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT25), .B(G183gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT26), .B(G190gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT24), .B1(new_n311_), .B2(new_n312_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321_));
  MUX2_X1   g120(.A(new_n320_), .B(KEYINPUT24), .S(new_n321_), .Z(new_n322_));
  AOI22_X1  g121(.A1(new_n310_), .A2(new_n315_), .B1(new_n319_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G197gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(G204gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT88), .B(G197gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(G204gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT21), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331_));
  INV_X1    g130(.A(G204gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n329_), .B1(G197gat), .B2(G204gat), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n333_), .A2(KEYINPUT89), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT89), .B1(new_n333_), .B2(new_n334_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n330_), .B(new_n331_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n324_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT20), .ZN(new_n341_));
  INV_X1    g140(.A(new_n339_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n308_), .A2(new_n309_), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n318_), .B(KEYINPUT91), .Z(new_n344_));
  INV_X1    g143(.A(new_n317_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n343_), .B(new_n322_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n315_), .B1(new_n316_), .B2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n341_), .B1(new_n342_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT19), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n323_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n359_), .B(KEYINPUT20), .C1(new_n349_), .C2(new_n342_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n352_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n353_), .A2(new_n358_), .A3(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(KEYINPUT100), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n363_), .B2(KEYINPUT100), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n350_), .A2(new_n361_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n358_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n360_), .A2(KEYINPUT92), .A3(new_n352_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT92), .B1(new_n360_), .B2(new_n352_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n367_), .B(new_n368_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n364_), .A2(new_n366_), .A3(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(KEYINPUT94), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n367_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n358_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(KEYINPUT94), .A3(new_n358_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n373_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT102), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n372_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT0), .ZN(new_n383_));
  INV_X1    g182(.A(G57gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(new_n203_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT95), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT86), .ZN(new_n391_));
  INV_X1    g190(.A(G155gat), .ZN(new_n392_));
  INV_X1    g191(.A(G162gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G141gat), .A2(G148gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT2), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G141gat), .A2(G148gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT3), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n397_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT87), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n404_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n395_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n399_), .A2(new_n396_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n391_), .A2(KEYINPUT1), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n391_), .A2(KEYINPUT1), .B1(new_n392_), .B2(new_n393_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G127gat), .B(G134gat), .Z(new_n415_));
  XOR2_X1   g214(.A(G113gat), .B(G120gat), .Z(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n417_), .A2(KEYINPUT85), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(KEYINPUT85), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n416_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n414_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n420_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n408_), .B(new_n413_), .C1(new_n417_), .C2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n421_), .B1(new_n407_), .B2(new_n412_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n389_), .B(new_n423_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n389_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n425_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n387_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n425_), .A2(KEYINPUT4), .A3(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n423_), .A2(new_n389_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n431_), .B(new_n387_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT31), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G71gat), .B(G99gat), .ZN(new_n439_));
  INV_X1    g238(.A(G43gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(G15gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n441_), .B(new_n444_), .Z(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n323_), .A2(KEYINPUT30), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n323_), .A2(KEYINPUT30), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n446_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n449_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(new_n447_), .A3(new_n445_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n438_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n452_), .A3(new_n438_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n454_), .A2(new_n421_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n421_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G228gat), .A2(G233gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT29), .B1(new_n407_), .B2(new_n412_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n460_), .B2(new_n339_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n339_), .A3(new_n459_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G78gat), .B(G106gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n460_), .A2(new_n339_), .A3(new_n459_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n464_), .B1(new_n467_), .B2(new_n461_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT90), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT90), .B1(new_n466_), .B2(new_n468_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G22gat), .B(G50gat), .Z(new_n471_));
  NOR2_X1   g270(.A1(new_n407_), .A2(new_n412_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT28), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n473_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n471_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n477_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n471_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n475_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n469_), .A2(new_n470_), .A3(new_n482_), .ZN(new_n483_));
  AND4_X1   g282(.A1(KEYINPUT90), .A2(new_n482_), .A3(new_n466_), .A4(new_n468_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n458_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n466_), .A2(new_n468_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT90), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n488_), .A2(new_n481_), .A3(new_n478_), .A4(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n456_), .A2(new_n457_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n469_), .B1(new_n470_), .B2(new_n482_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n437_), .B1(new_n485_), .B2(new_n493_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n375_), .A2(KEYINPUT94), .A3(new_n358_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n376_), .B2(new_n374_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT102), .B1(new_n496_), .B2(new_n373_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n381_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n483_), .A2(new_n484_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(new_n458_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n423_), .A2(new_n430_), .ZN(new_n501_));
  OAI221_X1 g300(.A(new_n386_), .B1(new_n427_), .B2(new_n430_), .C1(new_n434_), .C2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT97), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n436_), .B(KEYINPUT33), .ZN(new_n504_));
  AND4_X1   g303(.A1(new_n378_), .A2(new_n503_), .A3(new_n377_), .A4(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT98), .Z(new_n507_));
  OAI211_X1 g306(.A(new_n507_), .B(new_n367_), .C1(new_n370_), .C2(new_n369_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n353_), .A2(new_n362_), .A3(new_n506_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n437_), .A2(KEYINPUT99), .A3(new_n508_), .A4(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT99), .ZN(new_n511_));
  INV_X1    g310(.A(new_n436_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n512_), .B2(new_n432_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n508_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n511_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n500_), .B1(new_n505_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n498_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G29gat), .B(G36gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n244_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n521_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G232gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT34), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n263_), .A2(new_n524_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n522_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n528_), .A2(new_n525_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT73), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n522_), .B(new_n529_), .C1(new_n525_), .C2(new_n528_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT76), .ZN(new_n535_));
  XOR2_X1   g334(.A(G190gat), .B(G218gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT74), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G134gat), .B(G162gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT75), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n533_), .A2(new_n535_), .A3(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n539_), .B(new_n540_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT77), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT78), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT37), .B1(new_n543_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n533_), .A2(new_n535_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n545_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n533_), .A2(new_n535_), .A3(new_n542_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT14), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT79), .B(G1gat), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(G8gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT80), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G15gat), .B(G22gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G1gat), .B(G8gat), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n561_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n252_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT81), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n565_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G127gat), .B(G155gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT16), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G183gat), .B(G211gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT82), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n568_), .A2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n572_), .A2(new_n573_), .ZN(new_n577_));
  OAI22_X1  g376(.A1(new_n576_), .A2(KEYINPUT83), .B1(new_n568_), .B2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n576_), .A2(KEYINPUT83), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n518_), .A2(new_n555_), .A3(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n561_), .B(new_n562_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n521_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n564_), .A2(new_n524_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n521_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n564_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n587_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G169gat), .B(G197gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n591_), .B(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n302_), .A2(new_n581_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n437_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(new_n557_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT38), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT103), .ZN(new_n603_));
  INV_X1    g402(.A(new_n596_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n298_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n580_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n551_), .A2(new_n553_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n605_), .A2(new_n518_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n437_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n600_), .A2(new_n601_), .B1(G1gat), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n603_), .A2(new_n612_), .ZN(G1324gat));
  NAND2_X1  g412(.A1(new_n381_), .A2(new_n497_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n605_), .A2(new_n614_), .A3(new_n518_), .A4(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G8gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT104), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT104), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n618_), .A3(G8gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(G8gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n597_), .A2(new_n623_), .A3(new_n614_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n617_), .A2(KEYINPUT39), .A3(new_n619_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n622_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n622_), .A2(new_n624_), .A3(KEYINPUT40), .A4(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  AOI21_X1  g429(.A(new_n443_), .B1(new_n610_), .B2(new_n458_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n597_), .A2(new_n443_), .A3(new_n458_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n632_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(G1326gat));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n610_), .B2(new_n499_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT42), .Z(new_n639_));
  NAND3_X1  g438(.A1(new_n597_), .A2(new_n637_), .A3(new_n499_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1327gat));
  INV_X1    g440(.A(G29gat), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n580_), .A2(new_n607_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n605_), .A2(new_n518_), .A3(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n644_), .B2(new_n598_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n555_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n518_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n555_), .B1(new_n498_), .B2(new_n517_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n648_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n605_), .A2(new_n606_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n654_), .B1(new_n648_), .B2(new_n652_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(G29gat), .B(new_n437_), .C1(new_n659_), .C2(KEYINPUT44), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT107), .B(new_n645_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n663_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n645_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n664_), .A2(new_n668_), .ZN(G1328gat));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  INV_X1    g469(.A(G36gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n614_), .B1(new_n659_), .B2(KEYINPUT44), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n671_), .B1(new_n661_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n614_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n644_), .A2(G36gat), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n670_), .B1(new_n674_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n676_), .B(KEYINPUT45), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n672_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT46), .B(new_n680_), .C1(new_n681_), .C2(new_n671_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(G1329gat));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n440_), .B1(new_n644_), .B2(new_n491_), .ZN(new_n685_));
  OAI211_X1 g484(.A(G43gat), .B(new_n458_), .C1(new_n659_), .C2(KEYINPUT44), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n684_), .B(new_n685_), .C1(new_n662_), .C2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n685_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT47), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(G1330gat));
  INV_X1    g490(.A(new_n499_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n644_), .A2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(G50gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n659_), .A2(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n499_), .A2(G50gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n694_), .B1(new_n661_), .B2(new_n697_), .ZN(G1331gat));
  INV_X1    g497(.A(new_n301_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n300_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n596_), .B1(new_n498_), .B2(new_n517_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n701_), .A2(new_n702_), .A3(new_n609_), .A4(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n299_), .A2(new_n301_), .A3(new_n609_), .A4(new_n703_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT108), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n704_), .A2(new_n706_), .A3(G57gat), .A4(new_n437_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n581_), .A2(new_n298_), .A3(new_n604_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n384_), .B1(new_n708_), .B2(new_n598_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT109), .ZN(G1332gat));
  OR3_X1    g510(.A1(new_n708_), .A2(G64gat), .A3(new_n675_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n704_), .A2(new_n706_), .A3(new_n614_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G64gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G64gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT110), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n719_), .B(new_n712_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1333gat));
  OR3_X1    g520(.A1(new_n708_), .A2(G71gat), .A3(new_n491_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n704_), .A2(new_n706_), .A3(new_n458_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT49), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G71gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G71gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(G1334gat));
  OR3_X1    g526(.A1(new_n708_), .A2(G78gat), .A3(new_n692_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n704_), .A2(new_n706_), .A3(new_n499_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G78gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G78gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1335gat));
  NAND4_X1  g532(.A1(new_n299_), .A2(new_n301_), .A3(new_n643_), .A4(new_n703_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n735_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n203_), .A3(new_n437_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n648_), .A2(KEYINPUT112), .A3(new_n652_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n298_), .A2(new_n606_), .A3(new_n604_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n653_), .A2(new_n744_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n743_), .A2(new_n437_), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n739_), .B1(new_n746_), .B2(new_n203_), .ZN(G1336gat));
  AOI21_X1  g546(.A(G92gat), .B1(new_n738_), .B2(new_n614_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n750_));
  AND4_X1   g549(.A1(G92gat), .A2(new_n743_), .A3(new_n614_), .A4(new_n745_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(G1337gat));
  NAND4_X1  g551(.A1(new_n745_), .A2(new_n458_), .A3(new_n740_), .A4(new_n742_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G99gat), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n458_), .A2(new_n234_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n738_), .B2(new_n757_), .ZN(new_n758_));
  AOI211_X1 g557(.A(KEYINPUT114), .B(new_n756_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n754_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(new_n763_), .ZN(new_n764_));
  OAI221_X1 g563(.A(new_n754_), .B1(new_n761_), .B2(new_n762_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1338gat));
  NOR2_X1   g565(.A1(new_n741_), .A2(new_n692_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT43), .B1(new_n647_), .B2(KEYINPUT105), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n650_), .A2(new_n651_), .A3(new_n649_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(G106gat), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n770_), .A2(KEYINPUT116), .A3(new_n771_), .A4(G106gat), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(G106gat), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT52), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n738_), .A2(new_n212_), .A3(new_n499_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n778_), .A2(new_n782_), .A3(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1339gat));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n264_), .B(new_n253_), .C1(new_n267_), .C2(new_n276_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n257_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n277_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n255_), .A2(KEYINPUT68), .A3(new_n266_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n275_), .B1(new_n274_), .B2(KEYINPUT12), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n792_), .A2(KEYINPUT55), .A3(new_n264_), .A4(new_n265_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n789_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n788_), .A2(new_n277_), .B1(new_n786_), .B2(new_n257_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(KEYINPUT118), .A3(new_n793_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n282_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n785_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT118), .B1(new_n797_), .B2(new_n793_), .ZN(new_n802_));
  AND4_X1   g601(.A1(KEYINPUT118), .A2(new_n787_), .A3(new_n789_), .A4(new_n793_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n281_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n604_), .B1(new_n286_), .B2(new_n283_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n801_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n591_), .A2(new_n595_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n590_), .A2(new_n586_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n595_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n585_), .A2(new_n586_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n595_), .B1(new_n590_), .B2(new_n586_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(KEYINPUT120), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n290_), .A2(new_n808_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n807_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(KEYINPUT57), .A3(new_n607_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n785_), .B(new_n281_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n808_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n796_), .A2(new_n798_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n785_), .B1(new_n823_), .B2(new_n281_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT58), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n646_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n818_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n608_), .B1(new_n807_), .B2(new_n816_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(KEYINPUT57), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n606_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n555_), .A2(new_n580_), .A3(new_n604_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n298_), .A2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n614_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(G113gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n485_), .A2(new_n598_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n596_), .A4(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n555_), .B1(new_n825_), .B2(KEYINPUT58), .ZN(new_n842_));
  AOI22_X1  g641(.A1(KEYINPUT57), .A2(new_n831_), .B1(new_n842_), .B2(new_n828_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n817_), .A2(new_n607_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n580_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n835_), .B(new_n836_), .Z(new_n848_));
  OAI211_X1 g647(.A(new_n675_), .B(new_n840_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n833_), .A2(new_n837_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n852_), .A2(KEYINPUT59), .A3(new_n675_), .A4(new_n840_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n604_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n841_), .B1(new_n854_), .B2(new_n839_), .ZN(G1340gat));
  INV_X1    g654(.A(KEYINPUT60), .ZN(new_n856_));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n298_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n838_), .A2(new_n840_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n302_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n857_), .ZN(G1341gat));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n838_), .A2(new_n863_), .A3(new_n580_), .A4(new_n840_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n606_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n863_), .ZN(G1342gat));
  INV_X1    g665(.A(G134gat), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n838_), .A2(new_n867_), .A3(new_n608_), .A4(new_n840_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n555_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1343gat));
  NOR2_X1   g669(.A1(new_n493_), .A2(new_n598_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n838_), .A2(new_n596_), .A3(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g672(.A1(new_n838_), .A2(new_n701_), .A3(new_n871_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g674(.A1(new_n838_), .A2(new_n580_), .A3(new_n871_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  NAND2_X1  g677(.A1(new_n838_), .A2(new_n871_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G162gat), .B1(new_n879_), .B2(new_n555_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n608_), .A2(new_n393_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n879_), .B2(new_n881_), .ZN(G1347gat));
  NAND3_X1  g681(.A1(new_n614_), .A2(new_n598_), .A3(new_n458_), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT121), .Z(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n499_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n852_), .A2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G169gat), .B1(new_n886_), .B2(new_n604_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT62), .B(G169gat), .C1(new_n886_), .C2(new_n604_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n886_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n314_), .A3(new_n596_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n890_), .A3(new_n892_), .ZN(G1348gat));
  OAI21_X1  g692(.A(G176gat), .B1(new_n886_), .B2(new_n302_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n298_), .A2(new_n312_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n886_), .B2(new_n895_), .ZN(G1349gat));
  OAI21_X1  g695(.A(G183gat), .B1(new_n886_), .B2(new_n606_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n891_), .A2(new_n580_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n345_), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n886_), .B2(new_n555_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n607_), .A2(new_n344_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n886_), .B2(new_n901_), .ZN(G1351gat));
  NOR2_X1   g701(.A1(new_n493_), .A2(new_n437_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT122), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n675_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n852_), .A2(new_n596_), .A3(new_n905_), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n906_), .A2(KEYINPUT123), .A3(new_n325_), .ZN(new_n907_));
  AOI21_X1  g706(.A(KEYINPUT123), .B1(new_n906_), .B2(new_n325_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n325_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(G1352gat));
  NAND2_X1  g709(.A1(new_n852_), .A2(new_n905_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n302_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1353gat));
  INV_X1    g713(.A(new_n911_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n606_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT125), .Z(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT126), .Z(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n915_), .A2(new_n916_), .A3(new_n920_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1354gat));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n911_), .A2(new_n925_), .A3(new_n555_), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n852_), .A2(new_n608_), .A3(new_n905_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928_));
  AOI21_X1  g727(.A(G218gat), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT127), .B1(new_n911_), .B2(new_n607_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n926_), .B1(new_n929_), .B2(new_n930_), .ZN(G1355gat));
endmodule


