//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT79), .Z(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT22), .B(G169gat), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT81), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n212_), .B1(new_n209_), .B2(KEYINPUT23), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n211_), .B(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n207_), .B1(new_n208_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(KEYINPUT80), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n217_));
  OR3_X1    g016(.A1(new_n209_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n203_), .A2(new_n221_), .ZN(new_n222_));
  OR3_X1    g021(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT25), .B1(new_n225_), .B2(KEYINPUT78), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n225_), .A2(KEYINPUT25), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n224_), .B(new_n226_), .C1(new_n227_), .C2(KEYINPUT78), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n219_), .A2(new_n222_), .A3(new_n223_), .A4(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n215_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G43gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n230_), .B(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234_));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n233_), .B(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G227gat), .A2(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(G15gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n238_), .B(new_n243_), .Z(new_n244_));
  XNOR2_X1  g043(.A(G8gat), .B(G36gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT18), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G64gat), .B(G92gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G211gat), .B(G218gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT84), .B(G197gat), .ZN(new_n251_));
  INV_X1    g050(.A(G204gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT21), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n254_), .B1(G197gat), .B2(G204gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n250_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G197gat), .A2(G204gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(KEYINPUT84), .B(G197gat), .Z(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(G204gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n256_), .B1(KEYINPUT21), .B2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT21), .A3(new_n250_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT85), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT85), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n230_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT19), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n271_));
  INV_X1    g070(.A(new_n202_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n223_), .B1(new_n272_), .B2(new_n220_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n214_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT25), .B(G183gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT88), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n224_), .ZN(new_n277_));
  INV_X1    g076(.A(G190gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n225_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n219_), .A2(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n274_), .A2(new_n277_), .B1(new_n280_), .B2(new_n207_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n271_), .B1(new_n281_), .B2(new_n262_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n267_), .A2(new_n270_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n230_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT20), .B1(new_n281_), .B2(new_n262_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n269_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n283_), .B1(new_n286_), .B2(KEYINPUT89), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n264_), .A2(new_n266_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n230_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n285_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n288_), .B1(new_n293_), .B2(new_n269_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n249_), .B1(new_n287_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  OR2_X1    g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  OR2_X1    g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n304_), .B(new_n305_), .C1(new_n306_), .C2(KEYINPUT3), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n297_), .B(new_n298_), .C1(new_n301_), .C2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(G155gat), .A3(G162gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n297_), .A2(KEYINPUT1), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n310_), .B(new_n298_), .C1(new_n311_), .C2(KEYINPUT82), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(KEYINPUT82), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n306_), .B(new_n302_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n237_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n236_), .A2(new_n308_), .A3(new_n314_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(KEYINPUT4), .A3(new_n317_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n316_), .A2(KEYINPUT90), .A3(KEYINPUT4), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n236_), .B1(new_n314_), .B2(new_n308_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n320_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n296_), .B(new_n318_), .C1(new_n319_), .C2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G1gat), .B(G29gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G85gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT0), .B(G57gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n296_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n316_), .A2(new_n330_), .A3(new_n317_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n324_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n293_), .A2(new_n288_), .A3(new_n269_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n286_), .A2(KEYINPUT89), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n248_), .A4(new_n283_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n295_), .A2(new_n332_), .A3(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n330_), .B(new_n318_), .C1(new_n319_), .C2(new_n323_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n316_), .A2(new_n296_), .A3(new_n317_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT91), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n338_), .A2(KEYINPUT91), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n337_), .A2(new_n328_), .A3(new_n339_), .A4(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT92), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT33), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n337_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n329_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT93), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n341_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(KEYINPUT93), .A3(new_n329_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n291_), .A2(new_n270_), .A3(new_n292_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n267_), .A2(new_n282_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n352_), .B2(new_n270_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(KEYINPUT32), .A3(new_n248_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n248_), .A2(KEYINPUT32), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n333_), .A2(new_n334_), .A3(new_n283_), .A4(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  OAI22_X1  g156(.A1(new_n336_), .A2(new_n344_), .B1(new_n350_), .B2(new_n357_), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n315_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT28), .B1(new_n315_), .B2(KEYINPUT29), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G22gat), .B(G50gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n361_), .B(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G228gat), .A2(G233gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n315_), .A2(KEYINPUT29), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n264_), .A2(new_n266_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT86), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n265_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(G228gat), .A3(G233gat), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n364_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT87), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT87), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n364_), .B(new_n376_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n364_), .A2(new_n372_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n368_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n367_), .A2(new_n371_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n358_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n295_), .A2(new_n335_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n353_), .B2(new_n249_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n386_), .A2(new_n387_), .B1(new_n335_), .B2(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n378_), .A2(new_n382_), .B1(new_n349_), .B2(new_n348_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n244_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n389_), .A2(new_n384_), .A3(new_n350_), .A4(new_n244_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G1gat), .B(G8gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT74), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G22gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n240_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G15gat), .A2(G22gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G1gat), .A2(G8gat), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n400_), .A2(new_n401_), .B1(KEYINPUT14), .B2(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n398_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n398_), .A2(new_n403_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G29gat), .B(G36gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G43gat), .B(G50gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n398_), .B(new_n403_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n409_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G229gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n409_), .B(KEYINPUT15), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n411_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n414_), .A2(new_n416_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n421_), .A2(KEYINPUT76), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G113gat), .B(G141gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G169gat), .B(G197gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n421_), .B2(KEYINPUT76), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT77), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n420_), .A2(new_n427_), .A3(new_n425_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n422_), .A2(new_n426_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n395_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G57gat), .B(G64gat), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n433_), .A2(KEYINPUT11), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(KEYINPUT11), .ZN(new_n435_));
  XOR2_X1   g234(.A(G71gat), .B(G78gat), .Z(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n435_), .A2(new_n436_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(G106gat), .ZN(new_n441_));
  OR2_X1    g240(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n442_), .A2(KEYINPUT64), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT64), .B1(new_n442_), .B2(new_n443_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n441_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT6), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(G99gat), .A3(G106gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n446_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT9), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT65), .B(G85gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT66), .B(G92gat), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G85gat), .A2(G92gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n457_), .A2(new_n453_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT67), .ZN(new_n461_));
  INV_X1    g260(.A(G85gat), .ZN(new_n462_));
  INV_X1    g261(.A(G92gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n458_), .B1(KEYINPUT67), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n452_), .B1(new_n461_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT8), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n468_), .A2(KEYINPUT68), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(KEYINPUT68), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n457_), .A3(new_n464_), .A4(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n472_));
  INV_X1    g271(.A(G99gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n441_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n471_), .B1(new_n476_), .B2(new_n451_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n449_), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n447_), .A2(KEYINPUT6), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT69), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT69), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n448_), .A2(new_n450_), .A3(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n482_), .A3(new_n476_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n464_), .A2(new_n457_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n477_), .B1(new_n486_), .B2(KEYINPUT8), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n440_), .B1(new_n467_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n477_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n474_), .A2(new_n475_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(KEYINPUT69), .B2(new_n451_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n484_), .B1(new_n491_), .B2(new_n482_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n489_), .B1(new_n492_), .B2(new_n468_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n451_), .B(new_n446_), .C1(new_n495_), .C2(new_n465_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n493_), .A2(new_n496_), .A3(new_n439_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n488_), .A2(KEYINPUT12), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n496_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(new_n440_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G230gat), .A2(G233gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT70), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n488_), .A2(new_n497_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n503_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT70), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n506_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G120gat), .B(G148gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT5), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G176gat), .B(G204gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n512_), .A2(new_n517_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT13), .ZN(new_n520_));
  OR3_X1    g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT34), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n493_), .A2(new_n496_), .A3(new_n409_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n409_), .B(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n530_));
  OAI211_X1 g329(.A(KEYINPUT35), .B(new_n525_), .C1(new_n527_), .C2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G190gat), .B(G218gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT71), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G134gat), .B(G162gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(KEYINPUT36), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n499_), .A2(new_n418_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .A4(new_n526_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n531_), .A2(new_n536_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT72), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n531_), .A2(KEYINPUT72), .A3(new_n536_), .A4(new_n540_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n531_), .A2(new_n540_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n535_), .B(KEYINPUT36), .Z(new_n546_));
  AOI22_X1  g345(.A1(new_n543_), .A2(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT37), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n548_), .A2(KEYINPUT37), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n547_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G127gat), .B(G155gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT16), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n439_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n406_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n557_), .B1(new_n560_), .B2(KEYINPUT17), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n561_), .B1(KEYINPUT17), .B2(new_n557_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT75), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n562_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n553_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n523_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n432_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(G1gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n350_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT38), .Z(new_n572_));
  INV_X1    g371(.A(KEYINPUT95), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n547_), .B(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(KEYINPUT96), .B(new_n574_), .C1(new_n392_), .C2(new_n394_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n358_), .A2(new_n384_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n393_), .B1(new_n577_), .B2(new_n244_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT96), .B1(new_n578_), .B2(new_n574_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n431_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n521_), .A2(new_n581_), .A3(new_n522_), .A4(new_n565_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT94), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n569_), .B1(new_n585_), .B2(new_n570_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n572_), .A2(new_n586_), .ZN(G1324gat));
  INV_X1    g386(.A(G8gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n389_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n568_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n584_), .B(new_n589_), .C1(new_n576_), .C2(new_n579_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT97), .B(KEYINPUT39), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n591_), .A2(G8gat), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n591_), .B2(G8gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n590_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT99), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n597_), .B(new_n590_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1325gat));
  NAND2_X1  g401(.A1(new_n585_), .A2(new_n244_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n604_), .A2(KEYINPUT41), .A3(new_n240_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT41), .B1(new_n604_), .B2(new_n240_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n568_), .A2(new_n240_), .A3(new_n244_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT100), .Z(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n606_), .A3(new_n608_), .ZN(G1326gat));
  NAND3_X1  g408(.A1(new_n568_), .A2(new_n399_), .A3(new_n383_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n585_), .A2(new_n383_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n611_), .A2(G22gat), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n611_), .B2(G22gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n610_), .B1(new_n613_), .B2(new_n614_), .ZN(G1327gat));
  INV_X1    g414(.A(new_n565_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n547_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n523_), .A2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n432_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(G29gat), .B1(new_n619_), .B2(new_n570_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n523_), .A2(new_n431_), .A3(new_n565_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT43), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n578_), .A2(KEYINPUT102), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n553_), .B1(new_n578_), .B2(KEYINPUT102), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n622_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n553_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n622_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT103), .B1(new_n395_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n578_), .A2(new_n629_), .A3(new_n622_), .A4(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT44), .B(new_n621_), .C1(new_n625_), .C2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n621_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n623_), .A2(new_n624_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT43), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n628_), .A2(new_n630_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n633_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n638_));
  OAI21_X1  g437(.A(new_n632_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n570_), .A2(G29gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n620_), .B1(new_n640_), .B2(new_n641_), .ZN(G1328gat));
  OR2_X1    g441(.A1(new_n389_), .A2(KEYINPUT105), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n389_), .A2(KEYINPUT105), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(G36gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n432_), .A2(new_n618_), .A3(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT45), .Z(new_n649_));
  OAI211_X1 g448(.A(new_n589_), .B(new_n632_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(G36gat), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT46), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT106), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT107), .Z(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n651_), .B(new_n655_), .ZN(G1329gat));
  NAND2_X1  g455(.A1(new_n244_), .A2(G43gat), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n619_), .A2(new_n244_), .ZN(new_n658_));
  OAI22_X1  g457(.A1(new_n639_), .A2(new_n657_), .B1(G43gat), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g459(.A(G50gat), .B1(new_n619_), .B2(new_n383_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n383_), .A2(G50gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n640_), .B2(new_n662_), .ZN(G1331gat));
  INV_X1    g462(.A(new_n523_), .ZN(new_n664_));
  NOR4_X1   g463(.A1(new_n395_), .A2(new_n581_), .A3(new_n664_), .A4(new_n566_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G57gat), .B1(new_n665_), .B2(new_n570_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n664_), .A2(new_n581_), .A3(new_n616_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n580_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(G57gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n570_), .B2(KEYINPUT108), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(KEYINPUT108), .B2(new_n669_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n666_), .B1(new_n668_), .B2(new_n671_), .ZN(G1332gat));
  INV_X1    g471(.A(G64gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n665_), .A2(new_n673_), .A3(new_n645_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n668_), .A2(new_n645_), .ZN(new_n675_));
  XOR2_X1   g474(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(G64gat), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n675_), .B2(G64gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(G1333gat));
  INV_X1    g478(.A(G71gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n665_), .A2(new_n680_), .A3(new_n244_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n668_), .A2(new_n244_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G71gat), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT49), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(KEYINPUT49), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1334gat));
  INV_X1    g485(.A(G78gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n665_), .A2(new_n687_), .A3(new_n383_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n580_), .A2(new_n383_), .A3(new_n667_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT50), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n689_), .A2(new_n690_), .A3(G78gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n689_), .B2(G78gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1335gat));
  OR4_X1    g494(.A1(new_n395_), .A2(new_n581_), .A3(new_n664_), .A4(new_n617_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n570_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n664_), .A2(new_n581_), .A3(new_n565_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n699_), .B1(new_n625_), .B2(new_n631_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT111), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT111), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n702_), .B(new_n699_), .C1(new_n625_), .C2(new_n631_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n350_), .A2(new_n454_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n698_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(G1336gat));
  AOI21_X1  g507(.A(G92gat), .B1(new_n697_), .B2(new_n589_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n646_), .A2(new_n455_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT113), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n704_), .B2(new_n711_), .ZN(G1337gat));
  OAI211_X1 g511(.A(new_n697_), .B(new_n244_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n244_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n713_), .B1(new_n715_), .B2(new_n473_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n713_), .B(new_n717_), .C1(new_n715_), .C2(new_n473_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1338gat));
  XNOR2_X1  g520(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n383_), .B(new_n699_), .C1(new_n625_), .C2(new_n631_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(G106gat), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n724_), .A2(new_n723_), .A3(G106gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n697_), .A2(new_n441_), .A3(new_n383_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n722_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n727_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n729_), .B(new_n722_), .C1(new_n731_), .C2(new_n725_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1339gat));
  NAND2_X1  g533(.A1(new_n414_), .A2(new_n415_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n425_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n410_), .A2(new_n419_), .A3(new_n416_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n430_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n428_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n512_), .B2(new_n517_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n506_), .A2(new_n742_), .A3(new_n511_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n502_), .A2(new_n503_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(KEYINPUT55), .B2(new_n510_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT56), .B1(new_n746_), .B2(new_n516_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n748_), .B(new_n517_), .C1(new_n743_), .C2(new_n745_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n741_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT58), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n553_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n510_), .A2(KEYINPUT55), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(new_n503_), .B2(new_n502_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n510_), .B(new_n505_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n742_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n748_), .B1(new_n756_), .B2(new_n517_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n746_), .A2(KEYINPUT56), .A3(new_n516_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n759_), .A2(KEYINPUT116), .A3(KEYINPUT58), .A4(new_n741_), .ZN(new_n760_));
  OAI211_X1 g559(.A(KEYINPUT58), .B(new_n741_), .C1(new_n747_), .C2(new_n749_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n752_), .A2(new_n760_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n431_), .B1(new_n512_), .B2(new_n517_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n740_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n547_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n765_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT57), .B(new_n547_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n764_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n764_), .B(KEYINPUT117), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n616_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n567_), .B2(new_n431_), .ZN(new_n780_));
  NOR4_X1   g579(.A1(new_n523_), .A2(new_n566_), .A3(KEYINPUT54), .A4(new_n581_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n778_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n778_), .A2(KEYINPUT118), .A3(new_n783_), .ZN(new_n787_));
  NOR4_X1   g586(.A1(new_n589_), .A2(new_n350_), .A3(new_n714_), .A4(new_n383_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(G113gat), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n786_), .A2(KEYINPUT119), .A3(new_n787_), .A4(new_n788_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n581_), .A4(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n774_), .A2(new_n616_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(new_n782_), .ZN(new_n796_));
  XOR2_X1   g595(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n797_));
  NAND2_X1  g596(.A1(new_n788_), .A2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n431_), .B(new_n799_), .C1(new_n789_), .C2(KEYINPUT59), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n794_), .B1(new_n800_), .B2(new_n792_), .ZN(G1340gat));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n802_), .A2(KEYINPUT60), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n664_), .B2(KEYINPUT60), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n791_), .A2(new_n793_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n664_), .B(new_n799_), .C1(new_n789_), .C2(KEYINPUT59), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n802_), .ZN(G1341gat));
  INV_X1    g606(.A(G127gat), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n791_), .A2(new_n808_), .A3(new_n565_), .A4(new_n793_), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n616_), .B(new_n799_), .C1(new_n789_), .C2(KEYINPUT59), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n808_), .ZN(G1342gat));
  INV_X1    g610(.A(new_n574_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n791_), .A2(new_n812_), .A3(new_n793_), .ZN(new_n813_));
  INV_X1    g612(.A(G134gat), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n799_), .B1(new_n789_), .B2(KEYINPUT59), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n553_), .A2(new_n814_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT121), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n813_), .A2(new_n814_), .B1(new_n815_), .B2(new_n817_), .ZN(G1343gat));
  NOR3_X1   g617(.A1(new_n645_), .A2(new_n350_), .A3(new_n384_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n786_), .A2(new_n714_), .A3(new_n787_), .A4(new_n819_), .ZN(new_n820_));
  OR3_X1    g619(.A1(new_n820_), .A2(G141gat), .A3(new_n431_), .ZN(new_n821_));
  OAI21_X1  g620(.A(G141gat), .B1(new_n820_), .B2(new_n431_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1344gat));
  OR3_X1    g622(.A1(new_n820_), .A2(G148gat), .A3(new_n664_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G148gat), .B1(new_n820_), .B2(new_n664_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1345gat));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G155gat), .ZN(new_n827_));
  OR3_X1    g626(.A1(new_n820_), .A2(new_n616_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n820_), .B2(new_n616_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1346gat));
  OAI21_X1  g629(.A(G162gat), .B1(new_n820_), .B2(new_n553_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n574_), .A2(G162gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n820_), .B2(new_n832_), .ZN(G1347gat));
  NAND3_X1  g632(.A1(new_n645_), .A2(new_n350_), .A3(new_n244_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n383_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n581_), .B(new_n835_), .C1(new_n795_), .C2(new_n782_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(G169gat), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n837_), .A2(KEYINPUT122), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(KEYINPUT122), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(KEYINPUT62), .A3(new_n839_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n835_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n796_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n204_), .A3(new_n581_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n842_), .A2(new_n843_), .A3(new_n846_), .ZN(G1348gat));
  AOI21_X1  g646(.A(G176gat), .B1(new_n845_), .B2(new_n523_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n778_), .A2(KEYINPUT118), .A3(new_n783_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT118), .B1(new_n778_), .B2(new_n783_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n834_), .A2(new_n205_), .A3(new_n664_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n384_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n851_), .A2(KEYINPUT123), .A3(new_n384_), .A4(new_n852_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n848_), .B1(new_n855_), .B2(new_n856_), .ZN(G1349gat));
  NOR4_X1   g656(.A1(new_n796_), .A2(new_n276_), .A3(new_n616_), .A4(new_n844_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n834_), .A2(new_n616_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR4_X1   g659(.A1(new_n849_), .A2(new_n850_), .A3(new_n383_), .A4(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G183gat), .B1(new_n861_), .B2(KEYINPUT124), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n851_), .A2(new_n384_), .A3(new_n859_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n858_), .B1(new_n862_), .B2(new_n865_), .ZN(G1350gat));
  NAND2_X1  g665(.A1(new_n812_), .A2(new_n224_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT125), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n845_), .A2(new_n868_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n796_), .A2(new_n553_), .A3(new_n844_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n278_), .B2(new_n870_), .ZN(G1351gat));
  AND2_X1   g670(.A1(new_n645_), .A2(new_n390_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n786_), .A2(new_n714_), .A3(new_n787_), .A4(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G197gat), .B1(new_n874_), .B2(new_n581_), .ZN(new_n875_));
  INV_X1    g674(.A(G197gat), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n873_), .A2(new_n876_), .A3(new_n431_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1352gat));
  NOR2_X1   g677(.A1(new_n252_), .A2(KEYINPUT126), .ZN(new_n879_));
  OR3_X1    g678(.A1(new_n873_), .A2(new_n664_), .A3(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n873_), .B2(new_n664_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1353gat));
  XOR2_X1   g681(.A(KEYINPUT63), .B(G211gat), .Z(new_n883_));
  NAND3_X1  g682(.A1(new_n874_), .A2(new_n565_), .A3(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n873_), .B2(new_n616_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1354gat));
  NAND2_X1  g686(.A1(new_n874_), .A2(new_n812_), .ZN(new_n888_));
  INV_X1    g687(.A(G218gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n553_), .A2(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT127), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n888_), .A2(new_n889_), .B1(new_n874_), .B2(new_n891_), .ZN(G1355gat));
endmodule


