//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_;
  XOR2_X1   g000(.A(G120gat), .B(G148gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G176gat), .B(G204gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G230gat), .A2(G233gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT7), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  OAI22_X1  g014(.A1(new_n211_), .A2(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(G99gat), .A4(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n209_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(KEYINPUT8), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n220_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT67), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n224_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT8), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n220_), .A2(new_n230_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n216_), .B(new_n219_), .C1(G106gat), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT9), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n223_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n223_), .B2(new_n238_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n222_), .B1(new_n238_), .B2(new_n223_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n236_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n232_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n247_));
  INV_X1    g046(.A(G57gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(G64gat), .ZN(new_n249_));
  INV_X1    g048(.A(G64gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(G57gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n247_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(G57gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(G64gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(KEYINPUT68), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(new_n253_), .A3(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G71gat), .B(G78gat), .Z(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(new_n256_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(KEYINPUT11), .ZN(new_n262_));
  AOI211_X1 g061(.A(KEYINPUT69), .B(new_n253_), .C1(new_n252_), .C2(new_n256_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n259_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n254_), .A2(new_n255_), .A3(KEYINPUT68), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT68), .B1(new_n254_), .B2(new_n255_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT11), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT69), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n261_), .A2(new_n260_), .A3(KEYINPUT11), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n246_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n232_), .A3(new_n245_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n207_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT70), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n271_), .B1(new_n232_), .B2(new_n245_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(KEYINPUT12), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT12), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n273_), .A2(KEYINPUT72), .A3(new_n280_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n220_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n282_), .A2(new_n230_), .B1(KEYINPUT8), .B2(new_n228_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n244_), .B1(new_n283_), .B2(new_n227_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n264_), .A2(new_n270_), .A3(KEYINPUT12), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(new_n236_), .B2(new_n243_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n216_), .A2(new_n219_), .ZN(new_n289_));
  OAI221_X1 g088(.A(new_n222_), .B1(new_n238_), .B2(new_n223_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n235_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n215_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n289_), .A2(new_n290_), .A3(KEYINPUT71), .A4(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n232_), .A2(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n271_), .A2(new_n284_), .B1(new_n286_), .B2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n279_), .A2(new_n281_), .A3(new_n296_), .A4(new_n207_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n206_), .B1(new_n276_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n207_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n274_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n299_), .B1(new_n300_), .B2(new_n278_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT70), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n275_), .A2(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n297_), .A2(new_n302_), .A3(new_n304_), .A4(new_n206_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT13), .B1(new_n298_), .B2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n297_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n206_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT13), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(new_n305_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G29gat), .B(G36gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G43gat), .B(G50gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT15), .Z(new_n317_));
  XNOR2_X1  g116(.A(G15gat), .B(G22gat), .ZN(new_n318_));
  INV_X1    g117(.A(G1gat), .ZN(new_n319_));
  INV_X1    g118(.A(G8gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT14), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G8gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  OR2_X1    g123(.A1(new_n317_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G229gat), .A2(G233gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(new_n324_), .B2(new_n316_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n324_), .B(new_n316_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n325_), .A2(new_n328_), .B1(new_n329_), .B2(new_n327_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G113gat), .B(G141gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(G169gat), .B(G197gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n330_), .A2(new_n333_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n313_), .A2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n339_));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT83), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n342_), .A2(new_n343_), .A3(KEYINPUT83), .A4(new_n344_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(G169gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT25), .B(G183gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT26), .B(G190gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n352_), .A2(new_n353_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT24), .ZN(new_n358_));
  INV_X1    g157(.A(G169gat), .ZN(new_n359_));
  INV_X1    g158(.A(G176gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n351_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G71gat), .B(G99gat), .ZN(new_n366_));
  INV_X1    g165(.A(G43gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n365_), .A2(new_n368_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n339_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n339_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n369_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G134gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G127gat), .ZN(new_n378_));
  INV_X1    g177(.A(G127gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G134gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G120gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G113gat), .ZN(new_n383_));
  INV_X1    g182(.A(G113gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(G120gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n381_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G127gat), .B(G134gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G113gat), .B(G120gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n387_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n389_), .A3(KEYINPUT84), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G15gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT30), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n394_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n376_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n372_), .A2(new_n375_), .A3(new_n398_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G141gat), .A2(G148gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT88), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT2), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT2), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(KEYINPUT88), .A3(new_n406_), .ZN(new_n407_));
  OAI22_X1  g206(.A1(KEYINPUT87), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n405_), .A2(new_n407_), .A3(new_n408_), .A4(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n413_));
  INV_X1    g212(.A(G155gat), .ZN(new_n414_));
  INV_X1    g213(.A(G162gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n412_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(KEYINPUT1), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT1), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(G155gat), .A3(G162gat), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n416_), .A2(new_n421_), .A3(new_n423_), .A4(new_n417_), .ZN(new_n424_));
  XOR2_X1   g223(.A(G141gat), .B(G148gat), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n420_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n394_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT95), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n381_), .A2(new_n386_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n378_), .A2(new_n380_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n387_), .A2(new_n390_), .A3(KEYINPUT95), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n432_), .A2(new_n420_), .A3(new_n426_), .A4(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n428_), .A2(KEYINPUT4), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT4), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n427_), .A2(new_n438_), .A3(new_n394_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n428_), .A2(new_n436_), .A3(new_n434_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G1gat), .B(G29gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G57gat), .B(G85gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT99), .ZN(new_n449_));
  INV_X1    g248(.A(new_n447_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n440_), .A2(new_n450_), .A3(new_n441_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n442_), .A2(KEYINPUT99), .A3(new_n447_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G22gat), .B(G50gat), .Z(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n412_), .A2(new_n419_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT29), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n455_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n458_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n427_), .B2(KEYINPUT29), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n454_), .A3(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G78gat), .B(G106gat), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n461_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n467_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G228gat), .A2(G233gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n470_), .B(KEYINPUT90), .Z(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(G197gat), .A2(G204gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G197gat), .A2(G204gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(KEYINPUT21), .A3(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G211gat), .B(G218gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT91), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G218gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(G211gat), .ZN(new_n479_));
  INV_X1    g278(.A(G211gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G218gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  AND2_X1   g281(.A1(G197gat), .A2(G204gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G197gat), .A2(G204gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n482_), .A2(new_n485_), .A3(new_n486_), .A4(KEYINPUT21), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n477_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT92), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT21), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n475_), .A2(new_n491_), .A3(new_n476_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n488_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n489_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n427_), .A2(KEYINPUT29), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n472_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n488_), .A2(new_n492_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n496_), .A2(new_n498_), .A3(new_n472_), .ZN(new_n499_));
  OAI22_X1  g298(.A1(new_n468_), .A2(new_n469_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n461_), .A2(new_n465_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n466_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n497_), .A2(new_n499_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n461_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n452_), .A2(new_n453_), .B1(new_n500_), .B2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G8gat), .B(G36gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT18), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G64gat), .B(G92gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G226gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT19), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n365_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n362_), .A2(KEYINPUT93), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n361_), .A2(new_n342_), .A3(new_n519_), .A4(new_n344_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n357_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n350_), .A2(new_n345_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n517_), .B1(new_n523_), .B2(new_n498_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n514_), .B1(new_n516_), .B2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n513_), .A2(new_n517_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n523_), .B2(new_n498_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n495_), .B2(new_n365_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n511_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n498_), .A2(KEYINPUT92), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n488_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n365_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n523_), .A2(new_n498_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT20), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n513_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n527_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n365_), .A3(new_n531_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n510_), .A3(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n529_), .A2(new_n539_), .A3(KEYINPUT94), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT27), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n542_), .B(new_n511_), .C1(new_n525_), .C2(new_n528_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n540_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n539_), .A2(KEYINPUT101), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n510_), .B(KEYINPUT100), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n532_), .A2(new_n534_), .A3(new_n513_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n523_), .A2(new_n498_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n514_), .B1(new_n550_), .B2(new_n537_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n546_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT101), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n535_), .A2(new_n538_), .A3(new_n553_), .A4(new_n510_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n545_), .A2(KEYINPUT27), .A3(new_n552_), .A4(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n506_), .A2(new_n544_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n500_), .A2(new_n505_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n540_), .A2(new_n543_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n451_), .A2(KEYINPUT33), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT33), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n440_), .A2(new_n560_), .A3(new_n450_), .A4(new_n441_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n428_), .A2(new_n437_), .A3(new_n434_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n447_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT97), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n435_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n562_), .A2(new_n566_), .A3(new_n447_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n559_), .A2(new_n561_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n558_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n510_), .A2(KEYINPUT32), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n525_), .A2(new_n528_), .A3(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n571_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n452_), .A2(new_n453_), .A3(new_n572_), .A4(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n557_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n402_), .B1(new_n556_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n557_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n402_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n578_));
  AND4_X1   g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n544_), .A4(new_n555_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n338_), .B1(new_n576_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT37), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT74), .B(KEYINPUT35), .Z(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n586_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n232_), .A2(new_n316_), .A3(new_n245_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n317_), .B1(new_n232_), .B2(new_n294_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n588_), .B(new_n589_), .C1(new_n590_), .C2(KEYINPUT75), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n288_), .A2(new_n293_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n283_), .B2(new_n227_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT75), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n317_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n587_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n594_), .B1(new_n593_), .B2(new_n317_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n589_), .A2(new_n588_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n590_), .A2(KEYINPUT75), .ZN(new_n599_));
  INV_X1    g398(.A(new_n587_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .A4(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT76), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT36), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT77), .Z(new_n608_));
  NAND3_X1  g407(.A1(new_n596_), .A2(new_n601_), .A3(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n605_), .B(new_n606_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n596_), .B2(new_n601_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT79), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  AOI211_X1 g412(.A(KEYINPUT79), .B(new_n610_), .C1(new_n596_), .C2(new_n601_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n582_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT78), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n609_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n611_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n596_), .A2(new_n601_), .A3(KEYINPUT78), .A4(new_n608_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n617_), .A2(new_n618_), .A3(KEYINPUT37), .A4(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n615_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n324_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n264_), .A2(new_n623_), .A3(new_n270_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n264_), .B2(new_n270_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n622_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n271_), .A2(new_n324_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n628_), .A2(G231gat), .A3(G233gat), .A4(new_n624_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT17), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n635_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n627_), .A2(new_n629_), .A3(new_n637_), .A4(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT81), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n627_), .A2(new_n629_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(new_n636_), .ZN(new_n642_));
  AOI211_X1 g441(.A(KEYINPUT81), .B(new_n637_), .C1(new_n627_), .C2(new_n629_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT82), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT82), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n639_), .B(new_n646_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n621_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n581_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n451_), .A2(new_n449_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n450_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n453_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n651_), .A2(new_n319_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n657_), .A2(new_n658_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n644_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n338_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n576_), .A2(new_n580_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n613_), .A2(new_n614_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT102), .ZN(new_n665_));
  AND4_X1   g464(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .A4(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n319_), .B1(new_n666_), .B2(new_n656_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n659_), .A2(new_n660_), .A3(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT103), .Z(G1324gat));
  NAND2_X1  g468(.A1(new_n544_), .A2(new_n555_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n651_), .A2(new_n320_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n666_), .A2(new_n670_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n320_), .B1(KEYINPUT104), .B2(KEYINPUT39), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n673_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n671_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g477(.A(new_n402_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n666_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G15gat), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT105), .Z(new_n682_));
  OR2_X1    g481(.A1(new_n682_), .A2(KEYINPUT41), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(KEYINPUT41), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n650_), .A2(G15gat), .A3(new_n402_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(G1326gat));
  INV_X1    g485(.A(G22gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n557_), .B(KEYINPUT106), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n666_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT42), .Z(new_n691_));
  NAND3_X1  g490(.A1(new_n651_), .A2(new_n687_), .A3(new_n689_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1327gat));
  INV_X1    g492(.A(new_n664_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n648_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n581_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n656_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n663_), .A2(new_n701_), .A3(new_n621_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n570_), .A2(new_n574_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n577_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n506_), .A2(new_n544_), .A3(new_n555_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n679_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT108), .B1(new_n706_), .B2(new_n579_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n621_), .A2(KEYINPUT109), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n615_), .A2(new_n709_), .A3(new_n620_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n576_), .A2(new_n711_), .A3(new_n580_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n707_), .A2(new_n708_), .A3(new_n710_), .A4(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n714_));
  AOI21_X1  g513(.A(new_n702_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n338_), .A2(new_n695_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n700_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n714_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n572_), .A2(new_n573_), .ZN(new_n720_));
  AOI22_X1  g519(.A1(new_n656_), .A2(new_n720_), .B1(new_n558_), .B2(new_n569_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n705_), .B1(new_n721_), .B2(new_n557_), .ZN(new_n722_));
  AOI211_X1 g521(.A(KEYINPUT108), .B(new_n579_), .C1(new_n722_), .C2(new_n402_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n711_), .B1(new_n576_), .B2(new_n580_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n615_), .A2(new_n709_), .A3(new_n620_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n709_), .B1(new_n615_), .B2(new_n620_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n719_), .B1(new_n725_), .B2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT44), .B(new_n716_), .C1(new_n729_), .C2(new_n702_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n718_), .A2(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n656_), .A2(G29gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n699_), .B1(new_n731_), .B2(new_n732_), .ZN(G1328gat));
  XNOR2_X1  g532(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n718_), .A2(new_n730_), .A3(new_n670_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G36gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT110), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n735_), .A2(new_n738_), .A3(G36gat), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n670_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n697_), .A2(G36gat), .A3(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT45), .Z(new_n743_));
  AOI21_X1  g542(.A(new_n734_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n735_), .A2(new_n738_), .A3(G36gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n738_), .B1(new_n735_), .B2(G36gat), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n743_), .B(new_n734_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n744_), .A2(new_n748_), .ZN(G1329gat));
  NAND3_X1  g548(.A1(new_n731_), .A2(G43gat), .A3(new_n679_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n367_), .B1(new_n697_), .B2(new_n402_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g552(.A1(new_n697_), .A2(G50gat), .A3(new_n688_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n731_), .A2(new_n557_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n755_), .A2(KEYINPUT112), .A3(G50gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT112), .B1(new_n755_), .B2(G50gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n756_), .B2(new_n757_), .ZN(G1331gat));
  NAND3_X1  g557(.A1(new_n645_), .A2(new_n647_), .A3(new_n336_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n313_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n665_), .A2(new_n663_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n656_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G57gat), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n313_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n764_), .A2(new_n663_), .A3(new_n336_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n649_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n656_), .A2(new_n248_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1332gat));
  OAI21_X1  g567(.A(G64gat), .B1(new_n761_), .B2(new_n741_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT48), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n670_), .A2(new_n250_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n766_), .B2(new_n771_), .ZN(G1333gat));
  OAI21_X1  g571(.A(G71gat), .B1(new_n761_), .B2(new_n402_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT49), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n402_), .A2(G71gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n766_), .B2(new_n775_), .ZN(G1334gat));
  OAI21_X1  g575(.A(G78gat), .B1(new_n761_), .B2(new_n688_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT50), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n688_), .A2(G78gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n766_), .B2(new_n779_), .ZN(G1335gat));
  NAND2_X1  g579(.A1(new_n765_), .A2(new_n696_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(G85gat), .B1(new_n782_), .B2(new_n656_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n715_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n313_), .A2(new_n695_), .A3(new_n337_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n656_), .A2(G85gat), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT113), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n783_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT114), .ZN(G1336gat));
  INV_X1    g589(.A(G92gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n782_), .A2(new_n791_), .A3(new_n670_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n786_), .A2(new_n670_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n791_), .ZN(G1337gat));
  AND2_X1   g593(.A1(new_n786_), .A2(new_n679_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(new_n214_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n679_), .A2(new_n291_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n781_), .A2(new_n797_), .ZN(new_n798_));
  OR3_X1    g597(.A1(new_n796_), .A2(KEYINPUT51), .A3(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT51), .B1(new_n796_), .B2(new_n798_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1338gat));
  NAND3_X1  g600(.A1(new_n782_), .A2(new_n215_), .A3(new_n557_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n784_), .A2(new_n557_), .A3(new_n785_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805_));
  AND4_X1   g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n805_), .A4(G106gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n215_), .B1(KEYINPUT115), .B2(KEYINPUT52), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n804_), .A2(new_n807_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n802_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g609(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n759_), .A2(KEYINPUT116), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n645_), .A2(new_n813_), .A3(new_n647_), .A4(new_n336_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n812_), .A2(new_n313_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n621_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n811_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n812_), .A2(new_n313_), .A3(new_n814_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n811_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n818_), .A2(new_n621_), .A3(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n329_), .A2(new_n326_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n326_), .B1(new_n324_), .B2(new_n316_), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n333_), .B(new_n822_), .C1(new_n325_), .C2(new_n823_), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n334_), .B(new_n824_), .C1(new_n310_), .C2(new_n305_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n337_), .A2(new_n305_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n274_), .B1(new_n593_), .B2(new_n285_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n273_), .A2(new_n280_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n277_), .B2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(KEYINPUT55), .A3(new_n207_), .A4(new_n281_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n831_));
  NAND2_X1  g630(.A1(new_n297_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n279_), .A2(new_n281_), .A3(new_n296_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n299_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n309_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n826_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n835_), .A2(new_n309_), .A3(new_n837_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n825_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT57), .B1(new_n841_), .B2(new_n664_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n835_), .A2(new_n309_), .A3(new_n837_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n837_), .B1(new_n835_), .B2(new_n309_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n826_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n843_), .B(new_n694_), .C1(new_n846_), .C2(new_n825_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n836_), .A2(KEYINPUT56), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n835_), .A2(new_n849_), .A3(new_n309_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n306_), .A2(new_n334_), .A3(new_n824_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n852_), .A2(new_n853_), .B1(new_n615_), .B2(new_n620_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n842_), .A2(new_n847_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n821_), .B1(new_n856_), .B2(new_n661_), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n670_), .A2(new_n762_), .A3(new_n557_), .A4(new_n402_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(new_n384_), .A3(new_n337_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n821_), .B1(new_n856_), .B2(new_n695_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n858_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n859_), .A2(KEYINPUT59), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n866_), .A2(new_n337_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n861_), .B1(new_n867_), .B2(new_n384_), .ZN(G1340gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n764_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n866_), .A2(KEYINPUT120), .A3(new_n764_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(G120gat), .A3(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n382_), .B1(new_n313_), .B2(KEYINPUT60), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n860_), .B(new_n874_), .C1(KEYINPUT60), .C2(new_n382_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1341gat));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n859_), .A2(G127gat), .A3(new_n648_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n866_), .A2(new_n661_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n877_), .B(new_n879_), .C1(new_n880_), .C2(new_n379_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n379_), .B1(new_n866_), .B2(new_n661_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT121), .B1(new_n882_), .B2(new_n878_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1342gat));
  INV_X1    g683(.A(new_n665_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G134gat), .B1(new_n860_), .B2(new_n885_), .ZN(new_n886_));
  XOR2_X1   g685(.A(KEYINPUT122), .B(G134gat), .Z(new_n887_));
  NOR2_X1   g686(.A1(new_n816_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n866_), .B2(new_n888_), .ZN(G1343gat));
  NOR4_X1   g688(.A1(new_n670_), .A2(new_n679_), .A3(new_n762_), .A4(new_n577_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n857_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n337_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n764_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g694(.A1(new_n891_), .A2(new_n695_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT123), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n891_), .A2(new_n898_), .A3(new_n695_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n897_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n897_), .B2(new_n899_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1346gat));
  AOI21_X1  g702(.A(G162gat), .B1(new_n891_), .B2(new_n885_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n726_), .A2(new_n727_), .A3(new_n415_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n891_), .B2(new_n905_), .ZN(G1347gat));
  NAND2_X1  g705(.A1(new_n670_), .A2(new_n578_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n689_), .A2(new_n907_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n862_), .A2(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(KEYINPUT124), .A3(new_n337_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n862_), .A2(new_n337_), .A3(new_n908_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n359_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n910_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n910_), .B2(new_n913_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT22), .B(G169gat), .Z(new_n917_));
  OAI22_X1  g716(.A1(new_n915_), .A2(new_n916_), .B1(new_n911_), .B2(new_n917_), .ZN(G1348gat));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n313_), .A2(new_n907_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n857_), .A2(new_n921_), .A3(new_n577_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n857_), .B2(new_n577_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n920_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G176gat), .ZN(new_n925_));
  AND4_X1   g724(.A1(new_n360_), .A2(new_n862_), .A3(new_n764_), .A4(new_n908_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n919_), .B1(new_n925_), .B2(new_n927_), .ZN(new_n928_));
  AOI211_X1 g727(.A(KEYINPUT126), .B(new_n926_), .C1(new_n924_), .C2(G176gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1349gat));
  NOR2_X1   g729(.A1(new_n648_), .A2(new_n907_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n931_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n932_));
  INV_X1    g731(.A(G183gat), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n644_), .A2(new_n352_), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n932_), .A2(new_n933_), .B1(new_n909_), .B2(new_n934_), .ZN(G1350gat));
  NAND2_X1  g734(.A1(new_n909_), .A2(new_n621_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(G190gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n909_), .A2(new_n353_), .A3(new_n885_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1351gat));
  INV_X1    g738(.A(new_n857_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n670_), .A2(new_n506_), .A3(new_n402_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n337_), .ZN(new_n943_));
  INV_X1    g742(.A(G197gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(KEYINPUT127), .B1(new_n943_), .B2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n944_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n942_), .A2(new_n947_), .A3(G197gat), .A4(new_n337_), .ZN(new_n948_));
  AND3_X1   g747(.A1(new_n945_), .A2(new_n946_), .A3(new_n948_), .ZN(G1352gat));
  NAND2_X1  g748(.A1(new_n942_), .A2(new_n764_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g750(.A1(new_n940_), .A2(new_n644_), .A3(new_n941_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n952_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953_));
  XOR2_X1   g752(.A(KEYINPUT63), .B(G211gat), .Z(new_n954_));
  AOI21_X1  g753(.A(new_n953_), .B1(new_n952_), .B2(new_n954_), .ZN(G1354gat));
  NAND3_X1  g754(.A1(new_n942_), .A2(new_n478_), .A3(new_n885_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n940_), .A2(new_n816_), .A3(new_n941_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n478_), .B2(new_n957_), .ZN(G1355gat));
endmodule


