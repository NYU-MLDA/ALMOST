//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n969_, new_n970_, new_n971_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n982_, new_n983_, new_n985_, new_n986_,
    new_n988_, new_n989_, new_n990_, new_n992_, new_n993_, new_n994_,
    new_n995_;
  XOR2_X1   g000(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G155gat), .ZN(new_n204_));
  INV_X1    g003(.A(G162gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT88), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT88), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(G155gat), .B2(G162gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT90), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT90), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n213_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n212_), .A2(new_n214_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n220_), .A2(KEYINPUT91), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT91), .B1(new_n220_), .B2(new_n221_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n210_), .B1(new_n219_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n215_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n226_), .A2(new_n220_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT89), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n209_), .B2(KEYINPUT1), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n230_), .A2(KEYINPUT89), .A3(G155gat), .A4(G162gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n206_), .A2(new_n233_), .A3(new_n208_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n227_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n225_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G134gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G127gat), .ZN(new_n238_));
  INV_X1    g037(.A(G127gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G134gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G120gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G113gat), .ZN(new_n243_));
  INV_X1    g042(.A(G113gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G120gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n238_), .A2(new_n240_), .A3(new_n243_), .A4(new_n245_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(KEYINPUT87), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n241_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT87), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(new_n243_), .A4(new_n245_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n236_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n248_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n225_), .A2(new_n235_), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(KEYINPUT4), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n260_));
  AND4_X1   g059(.A1(KEYINPUT97), .A2(new_n236_), .A3(new_n260_), .A4(new_n253_), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n225_), .A2(new_n235_), .B1(new_n252_), .B2(new_n249_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT97), .B1(new_n262_), .B2(new_n260_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n257_), .B(new_n259_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n220_), .A2(new_n221_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT91), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n220_), .A2(KEYINPUT91), .A3(new_n221_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n216_), .B2(new_n215_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n269_), .A2(new_n214_), .A3(new_n212_), .A4(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n229_), .A2(new_n231_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n206_), .A2(new_n233_), .A3(new_n208_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n272_), .A2(new_n210_), .B1(new_n275_), .B2(new_n227_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n249_), .A2(new_n252_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n256_), .B(new_n258_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G1gat), .B(G29gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G57gat), .B(G85gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n203_), .B1(new_n264_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n254_), .A2(new_n256_), .A3(new_n259_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n283_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n225_), .A2(new_n235_), .A3(new_n255_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(new_n262_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n259_), .B1(new_n291_), .B2(KEYINPUT4), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n236_), .A2(new_n260_), .A3(new_n253_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT97), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n262_), .A2(KEYINPUT97), .A3(new_n260_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n289_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n278_), .A2(KEYINPUT33), .A3(new_n283_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n258_), .B1(new_n291_), .B2(KEYINPUT4), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n300_), .B2(new_n297_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n286_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT93), .ZN(new_n304_));
  XOR2_X1   g103(.A(G197gat), .B(G204gat), .Z(new_n305_));
  AND3_X1   g104(.A1(new_n304_), .A2(KEYINPUT21), .A3(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n303_), .A2(KEYINPUT93), .ZN(new_n307_));
  XOR2_X1   g106(.A(G211gat), .B(G218gat), .Z(new_n308_));
  INV_X1    g107(.A(KEYINPUT21), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT92), .ZN(new_n312_));
  INV_X1    g111(.A(G197gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(G204gat), .ZN(new_n314_));
  OAI211_X1 g113(.A(KEYINPUT21), .B(new_n314_), .C1(new_n305_), .C2(new_n312_), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n306_), .A2(new_n307_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G169gat), .ZN(new_n317_));
  INV_X1    g116(.A(G176gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(KEYINPUT82), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT82), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(G169gat), .B2(G176gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n319_), .A2(new_n321_), .A3(KEYINPUT24), .A4(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G183gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT78), .B1(new_n325_), .B2(KEYINPUT25), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(G183gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(KEYINPUT80), .A2(KEYINPUT26), .ZN(new_n331_));
  NOR2_X1   g130(.A1(KEYINPUT80), .A2(KEYINPUT26), .ZN(new_n332_));
  OAI21_X1  g131(.A(G190gat), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT79), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G190gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n337_), .A3(KEYINPUT26), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n328_), .A2(G183gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n330_), .A2(new_n333_), .A3(new_n338_), .A4(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n324_), .B1(new_n341_), .B2(KEYINPUT81), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT24), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n320_), .A2(G169gat), .A3(G176gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT82), .B1(new_n317_), .B2(new_n318_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n343_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n346_), .A2(KEYINPUT83), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT24), .B1(new_n319_), .B2(new_n321_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n354_), .B1(new_n355_), .B2(new_n351_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT79), .B(G190gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n339_), .B1(new_n358_), .B2(KEYINPUT26), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT81), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n333_), .A4(new_n330_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n342_), .A2(new_n357_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT22), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(G169gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G169gat), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n318_), .B(new_n365_), .C1(new_n366_), .C2(new_n363_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n358_), .A2(new_n325_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n367_), .B(new_n322_), .C1(new_n368_), .C2(new_n351_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n316_), .B1(new_n362_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT19), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n311_), .A2(new_n315_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n307_), .A2(KEYINPUT21), .A3(new_n305_), .A4(new_n304_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT25), .B(G183gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT26), .B(G190gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n346_), .A2(new_n378_), .A3(new_n352_), .A4(new_n323_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n366_), .A2(new_n318_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n380_), .B(new_n322_), .C1(new_n351_), .C2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT20), .B1(new_n375_), .B2(new_n383_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n370_), .A2(new_n372_), .A3(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n372_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n341_), .A2(KEYINPUT81), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(new_n361_), .A3(new_n323_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT83), .B1(new_n346_), .B2(new_n352_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n355_), .A2(new_n354_), .A3(new_n351_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n316_), .B(new_n369_), .C1(new_n393_), .C2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT20), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(new_n375_), .B2(new_n383_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n391_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n385_), .A2(new_n390_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n390_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n362_), .A2(new_n369_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n375_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n384_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n391_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n397_), .A2(new_n399_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n372_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n402_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n401_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT100), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n302_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n402_), .A2(KEYINPUT32), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n372_), .B1(new_n370_), .B2(new_n384_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n397_), .A2(new_n391_), .A3(new_n399_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n385_), .A2(new_n400_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(new_n413_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n264_), .A2(new_n278_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n288_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n264_), .A2(new_n285_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n257_), .B(new_n258_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n289_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n278_), .A2(KEYINPUT33), .A3(new_n283_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n264_), .A2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n284_), .B1(new_n300_), .B2(new_n297_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n426_), .B(new_n428_), .C1(new_n429_), .C2(new_n203_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n390_), .B1(new_n385_), .B2(new_n400_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n406_), .A2(new_n408_), .A3(new_n402_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT100), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n412_), .A2(new_n423_), .A3(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G22gat), .B(G50gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT28), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n436_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G78gat), .B(G106gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT94), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G228gat), .A2(G233gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n375_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT29), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n225_), .B2(new_n235_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n447_), .B2(new_n316_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n441_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT95), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n439_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n441_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n443_), .B1(new_n442_), .B2(new_n375_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n447_), .A2(new_n316_), .A3(new_n445_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n444_), .A2(new_n448_), .A3(new_n441_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n455_), .A2(new_n439_), .A3(new_n450_), .A4(new_n456_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n435_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT27), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n433_), .A2(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n414_), .A2(new_n415_), .ZN(new_n464_));
  OAI211_X1 g263(.A(KEYINPUT27), .B(new_n432_), .C1(new_n464_), .C2(new_n402_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n429_), .B1(new_n288_), .B2(new_n419_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(new_n459_), .A3(new_n458_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT101), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n460_), .A2(new_n422_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT101), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n463_), .A4(new_n465_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n461_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n403_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n362_), .A2(new_n369_), .A3(new_n474_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G71gat), .B(G99gat), .ZN(new_n480_));
  INV_X1    g279(.A(G43gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G227gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(G15gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n482_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n277_), .B(KEYINPUT31), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n476_), .A2(new_n478_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT86), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n490_), .A2(new_n479_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n487_), .B(new_n488_), .C1(new_n491_), .C2(new_n486_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n488_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n486_), .B1(new_n490_), .B2(new_n479_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n487_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n492_), .A2(new_n496_), .A3(new_n467_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n463_), .A2(new_n460_), .A3(new_n465_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT102), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n500_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT102), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n497_), .A2(new_n502_), .A3(new_n503_), .A4(new_n467_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n473_), .A2(new_n498_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT15), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G29gat), .B(G36gat), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(KEYINPUT69), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(KEYINPUT69), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n506_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n508_), .A2(new_n509_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n510_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT15), .A3(new_n511_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520_));
  INV_X1    g319(.A(G1gat), .ZN(new_n521_));
  INV_X1    g320(.A(G8gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G8gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n517_), .A2(new_n511_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(new_n526_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n528_), .A3(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n532_), .A2(KEYINPUT76), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n529_), .B(new_n526_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n532_), .B(KEYINPUT76), .C1(new_n528_), .C2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G113gat), .B(G141gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G169gat), .B(G197gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  OR2_X1    g337(.A1(new_n538_), .A2(KEYINPUT77), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n533_), .A2(new_n535_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n539_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n505_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT37), .ZN(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT10), .B(G99gat), .Z(new_n546_));
  INV_X1    g345(.A(G106gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G85gat), .B(G92gat), .Z(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT9), .ZN(new_n550_));
  INV_X1    g349(.A(G85gat), .ZN(new_n551_));
  INV_X1    g350(.A(G92gat), .ZN(new_n552_));
  OR3_X1    g351(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT9), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n548_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT64), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(KEYINPUT6), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(KEYINPUT6), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT6), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(KEYINPUT64), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n558_), .B1(new_n556_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n554_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT65), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT66), .ZN(new_n570_));
  INV_X1    g369(.A(G99gat), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n547_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n573_));
  OR2_X1    g372(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n574_));
  NAND2_X1  g373(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n569_), .A2(new_n561_), .A3(new_n564_), .A4(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT8), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n549_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n577_), .B2(new_n549_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n567_), .B(new_n529_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT70), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT34), .Z(new_n584_));
  INV_X1    g383(.A(KEYINPUT35), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n585_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n580_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n577_), .A2(new_n578_), .A3(new_n549_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n566_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n514_), .A2(new_n518_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n581_), .B(new_n588_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n587_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT74), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n567_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n519_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n597_), .A2(new_n582_), .A3(new_n581_), .A4(new_n586_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n594_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n595_), .B1(new_n594_), .B2(new_n598_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT71), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT36), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n599_), .A2(new_n600_), .A3(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n594_), .B2(new_n598_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n545_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT72), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n612_), .B(new_n608_), .C1(new_n594_), .C2(new_n598_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n594_), .A2(new_n598_), .A3(new_n605_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n545_), .B1(new_n616_), .B2(KEYINPUT73), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT73), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n594_), .A2(new_n618_), .A3(new_n598_), .A4(new_n605_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n613_), .A2(new_n615_), .A3(new_n617_), .A4(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n610_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT13), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G57gat), .B(G64gat), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT11), .ZN(new_n624_));
  XOR2_X1   g423(.A(G71gat), .B(G78gat), .Z(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n624_), .A2(new_n625_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n623_), .A2(KEYINPUT11), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n596_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT12), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n596_), .A2(new_n629_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n596_), .A2(KEYINPUT68), .A3(KEYINPUT12), .A4(new_n629_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n596_), .A2(KEYINPUT12), .A3(new_n629_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT68), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .A4(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n630_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n632_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n634_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT5), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n645_), .B(new_n646_), .Z(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n639_), .A2(new_n643_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n648_), .B1(new_n639_), .B2(new_n643_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n622_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n651_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(KEYINPUT13), .A3(new_n649_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(G231gat), .A2(G233gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n526_), .B(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(new_n629_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT75), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(G127gat), .B(G155gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT16), .ZN(new_n662_));
  XNOR2_X1  g461(.A(G183gat), .B(G211gat), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT17), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n660_), .B(new_n665_), .ZN(new_n666_));
  OR3_X1    g465(.A1(new_n658_), .A2(KEYINPUT17), .A3(new_n664_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n621_), .A2(new_n655_), .A3(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n544_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n521_), .A3(new_n422_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT38), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n607_), .A2(new_n609_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n505_), .A2(new_n675_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n655_), .A2(new_n543_), .A3(new_n669_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n521_), .B1(new_n678_), .B2(new_n422_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n674_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n680_), .B1(new_n673_), .B2(new_n672_), .ZN(G1324gat));
  AOI21_X1  g480(.A(new_n522_), .B1(new_n678_), .B2(new_n466_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT39), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n671_), .A2(new_n522_), .A3(new_n466_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(G1325gat));
  AOI21_X1  g486(.A(new_n484_), .B1(new_n678_), .B2(new_n497_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT41), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n671_), .A2(new_n484_), .A3(new_n497_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1326gat));
  INV_X1    g490(.A(G22gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n460_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n678_), .B2(new_n693_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT42), .Z(new_n695_));
  NAND3_X1  g494(.A1(new_n671_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1327gat));
  INV_X1    g496(.A(new_n675_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n655_), .A2(new_n698_), .A3(new_n668_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n544_), .A2(new_n699_), .ZN(new_n700_));
  OR3_X1    g499(.A1(new_n700_), .A2(G29gat), .A3(new_n467_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n655_), .A2(new_n543_), .A3(new_n668_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n616_), .A2(KEYINPUT73), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT37), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n619_), .B1(new_n609_), .B2(KEYINPUT72), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n705_), .A2(new_n706_), .A3(new_n614_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n594_), .A2(new_n598_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT74), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n594_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n605_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT37), .B1(new_n711_), .B2(new_n611_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT103), .B1(new_n707_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n610_), .A2(new_n714_), .A3(new_n620_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n505_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n469_), .A2(new_n472_), .ZN(new_n718_));
  AOI22_X1  g517(.A1(new_n424_), .A2(new_n425_), .B1(new_n264_), .B2(new_n427_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n421_), .A2(new_n202_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n432_), .A4(new_n431_), .ZN(new_n721_));
  AOI22_X1  g520(.A1(new_n721_), .A2(KEYINPUT100), .B1(new_n422_), .B2(new_n418_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n693_), .B1(new_n722_), .B2(new_n412_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n498_), .B1(new_n718_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n504_), .A2(new_n501_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n621_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n703_), .B1(new_n717_), .B2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT104), .B1(new_n729_), .B2(KEYINPUT44), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n707_), .A2(new_n712_), .A3(KEYINPUT103), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n714_), .B1(new_n610_), .B2(new_n620_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n727_), .B1(new_n726_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n621_), .A2(new_n727_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n702_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n730_), .A2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT44), .B(new_n702_), .C1(new_n734_), .C2(new_n736_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n422_), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(G29gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(G29gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n701_), .B1(new_n745_), .B2(new_n746_), .ZN(G1328gat));
  INV_X1    g546(.A(new_n466_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n700_), .A2(G36gat), .A3(new_n748_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT45), .Z(new_n750_));
  NAND2_X1  g549(.A1(new_n742_), .A2(new_n466_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n729_), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n738_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT106), .B1(new_n755_), .B2(G36gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n751_), .B1(new_n730_), .B2(new_n740_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n758_));
  INV_X1    g557(.A(G36gat), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n750_), .B1(new_n756_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(KEYINPUT46), .B(new_n750_), .C1(new_n756_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1329gat));
  XNOR2_X1  g564(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n741_), .A2(G43gat), .A3(new_n497_), .A4(new_n742_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n481_), .B1(new_n700_), .B2(new_n498_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n767_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n768_), .A2(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT108), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n766_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n773_), .A2(new_n777_), .ZN(G1330gat));
  AND3_X1   g577(.A1(new_n741_), .A2(new_n693_), .A3(new_n742_), .ZN(new_n779_));
  INV_X1    g578(.A(G50gat), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n693_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT109), .ZN(new_n782_));
  OAI22_X1  g581(.A1(new_n779_), .A2(new_n780_), .B1(new_n700_), .B2(new_n782_), .ZN(G1331gat));
  NAND4_X1  g582(.A1(new_n676_), .A2(new_n543_), .A3(new_n655_), .A4(new_n668_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT111), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G57gat), .B1(new_n786_), .B2(new_n467_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n726_), .A2(new_n543_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT110), .ZN(new_n789_));
  INV_X1    g588(.A(new_n621_), .ZN(new_n790_));
  AND4_X1   g589(.A1(new_n655_), .A2(new_n789_), .A3(new_n668_), .A4(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(G57gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n422_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n787_), .A2(new_n793_), .ZN(G1332gat));
  INV_X1    g593(.A(G64gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n785_), .B2(new_n466_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT48), .Z(new_n797_));
  NAND3_X1  g596(.A1(new_n791_), .A2(new_n795_), .A3(new_n466_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1333gat));
  INV_X1    g598(.A(G71gat), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n791_), .A2(new_n800_), .A3(new_n497_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n785_), .A2(new_n497_), .ZN(new_n802_));
  XOR2_X1   g601(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n803_));
  AND3_X1   g602(.A1(new_n802_), .A2(G71gat), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n802_), .B2(G71gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(G1334gat));
  INV_X1    g605(.A(G78gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n791_), .A2(new_n807_), .A3(new_n693_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n785_), .A2(new_n693_), .ZN(new_n809_));
  XOR2_X1   g608(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(G78gat), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n809_), .B2(G78gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(G1335gat));
  AND4_X1   g612(.A1(new_n655_), .A2(new_n789_), .A3(new_n669_), .A4(new_n675_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n551_), .A3(new_n422_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n717_), .A2(new_n728_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n655_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n817_), .A2(new_n542_), .A3(new_n668_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G85gat), .B1(new_n819_), .B2(new_n467_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n820_), .ZN(G1336gat));
  NAND3_X1  g620(.A1(new_n814_), .A2(new_n552_), .A3(new_n466_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G92gat), .B1(new_n819_), .B2(new_n748_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1337gat));
  NAND3_X1  g623(.A1(new_n814_), .A2(new_n497_), .A3(new_n546_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n819_), .A2(new_n498_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n571_), .B2(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n816_), .A2(new_n693_), .A3(new_n818_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(G106gat), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n831_), .B1(new_n830_), .B2(G106gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n829_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n834_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(KEYINPUT52), .A3(new_n832_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n814_), .A2(new_n547_), .A3(new_n693_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1339gat));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n670_), .B2(new_n543_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n790_), .A2(new_n817_), .A3(new_n543_), .A4(new_n668_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(KEYINPUT54), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n845_), .B2(KEYINPUT116), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n844_), .B2(KEYINPUT54), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n538_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n528_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n534_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT117), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n527_), .A2(new_n852_), .A3(new_n531_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(new_n850_), .C1(new_n534_), .C2(new_n852_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n854_), .A2(KEYINPUT118), .A3(new_n855_), .A4(new_n857_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n851_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n862_), .A2(new_n649_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT55), .ZN(new_n864_));
  INV_X1    g663(.A(new_n629_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n631_), .B1(new_n591_), .B2(new_n865_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n638_), .A2(new_n640_), .A3(new_n866_), .A4(new_n635_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n864_), .B1(new_n867_), .B2(new_n642_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n642_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT56), .B1(new_n870_), .B2(new_n647_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n868_), .A2(new_n869_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n867_), .A2(new_n864_), .A3(new_n642_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT56), .B(new_n647_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n863_), .B1(new_n871_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n863_), .B(KEYINPUT58), .C1(new_n871_), .C2(new_n875_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n879_), .A3(new_n621_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n542_), .A2(new_n649_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n647_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n881_), .B1(new_n884_), .B2(new_n874_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n653_), .A2(new_n649_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n862_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n698_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  OAI211_X1 g689(.A(KEYINPUT57), .B(new_n698_), .C1(new_n885_), .C2(new_n887_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n880_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n669_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n849_), .A2(new_n893_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n498_), .A2(new_n500_), .A3(new_n467_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n244_), .B1(new_n896_), .B2(new_n543_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n848_), .A2(new_n846_), .B1(new_n892_), .B2(new_n669_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT59), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n846_), .A2(new_n848_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n893_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n892_), .A2(KEYINPUT120), .A3(new_n669_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n901_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(KEYINPUT59), .B1(new_n895_), .B2(KEYINPUT119), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(KEYINPUT119), .B2(new_n895_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n900_), .B1(new_n905_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n542_), .A2(G113gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n897_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  OAI211_X1 g711(.A(KEYINPUT121), .B(new_n897_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1340gat));
  XNOR2_X1  g713(.A(KEYINPUT122), .B(G120gat), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n896_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n817_), .B2(new_n916_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n655_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n916_), .B1(new_n921_), .B2(new_n908_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1341gat));
  OAI21_X1  g723(.A(G127gat), .B1(new_n908_), .B2(new_n669_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n917_), .A2(new_n239_), .A3(new_n668_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1342gat));
  OAI21_X1  g726(.A(G134gat), .B1(new_n908_), .B2(new_n790_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n917_), .A2(new_n237_), .A3(new_n675_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1343gat));
  NOR2_X1   g729(.A1(new_n497_), .A2(new_n460_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n466_), .A2(new_n467_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n894_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n542_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n655_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n934_), .A2(new_n939_), .A3(new_n668_), .ZN(new_n940_));
  OAI21_X1  g739(.A(KEYINPUT123), .B1(new_n933_), .B2(new_n669_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT61), .B(G155gat), .ZN(new_n942_));
  AND3_X1   g741(.A1(new_n940_), .A2(new_n941_), .A3(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1346gat));
  NOR3_X1   g744(.A1(new_n933_), .A2(new_n205_), .A3(new_n716_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n934_), .A2(new_n675_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n205_), .ZN(G1347gat));
  INV_X1    g747(.A(new_n904_), .ZN(new_n949_));
  AOI21_X1  g748(.A(KEYINPUT120), .B1(new_n892_), .B2(new_n669_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n849_), .B1(new_n949_), .B2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n499_), .A2(new_n748_), .ZN(new_n952_));
  XOR2_X1   g751(.A(new_n952_), .B(KEYINPUT124), .Z(new_n953_));
  NOR2_X1   g752(.A1(new_n953_), .A2(new_n693_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n951_), .A2(new_n954_), .ZN(new_n955_));
  OAI21_X1  g754(.A(G169gat), .B1(new_n955_), .B2(new_n543_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n954_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n903_), .A2(new_n904_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n959_), .B1(new_n960_), .B2(new_n849_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n961_), .A2(new_n366_), .A3(new_n542_), .ZN(new_n962_));
  OAI211_X1 g761(.A(KEYINPUT62), .B(G169gat), .C1(new_n955_), .C2(new_n543_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n958_), .A2(new_n962_), .A3(new_n963_), .ZN(G1348gat));
  AOI21_X1  g763(.A(G176gat), .B1(new_n961_), .B2(new_n655_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n898_), .A2(new_n693_), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n953_), .A2(new_n318_), .A3(new_n817_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(G1349gat));
  NOR2_X1   g767(.A1(new_n953_), .A2(new_n669_), .ZN(new_n969_));
  AOI21_X1  g768(.A(G183gat), .B1(new_n966_), .B2(new_n969_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n669_), .A2(new_n376_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n970_), .B1(new_n961_), .B2(new_n971_), .ZN(G1350gat));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n334_), .B1(new_n961_), .B2(new_n621_), .ZN(new_n974_));
  AND2_X1   g773(.A1(new_n675_), .A2(new_n377_), .ZN(new_n975_));
  AND3_X1   g774(.A1(new_n951_), .A2(new_n954_), .A3(new_n975_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n973_), .B1(new_n974_), .B2(new_n976_), .ZN(new_n977_));
  OAI21_X1  g776(.A(G190gat), .B1(new_n955_), .B2(new_n790_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n961_), .A2(new_n975_), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n978_), .A2(KEYINPUT125), .A3(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n977_), .A2(new_n980_), .ZN(G1351gat));
  NAND4_X1  g780(.A1(new_n894_), .A2(new_n467_), .A3(new_n466_), .A4(new_n931_), .ZN(new_n982_));
  NOR2_X1   g781(.A1(new_n982_), .A2(new_n543_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(new_n983_), .B(new_n313_), .ZN(G1352gat));
  INV_X1    g783(.A(new_n982_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n985_), .A2(new_n655_), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n986_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g786(.A(new_n669_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n988_));
  AND2_X1   g787(.A1(new_n985_), .A2(new_n988_), .ZN(new_n989_));
  NOR2_X1   g788(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n990_));
  XNOR2_X1  g789(.A(new_n989_), .B(new_n990_), .ZN(G1354gat));
  NAND2_X1  g790(.A1(new_n985_), .A2(new_n675_), .ZN(new_n992_));
  XOR2_X1   g791(.A(KEYINPUT126), .B(G218gat), .Z(new_n993_));
  NOR2_X1   g792(.A1(new_n790_), .A2(new_n993_), .ZN(new_n994_));
  XOR2_X1   g793(.A(new_n994_), .B(KEYINPUT127), .Z(new_n995_));
  AOI22_X1  g794(.A1(new_n992_), .A2(new_n993_), .B1(new_n985_), .B2(new_n995_), .ZN(G1355gat));
endmodule


