//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_, new_n960_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G1gat), .A2(G8gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(new_n207_), .A3(KEYINPUT14), .ZN(new_n208_));
  INV_X1    g007(.A(G15gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G22gat), .ZN(new_n210_));
  INV_X1    g009(.A(G22gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G15gat), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n208_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  AND2_X1   g012(.A1(G1gat), .A2(G8gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G1gat), .A2(G8gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT74), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G1gat), .ZN(new_n217_));
  INV_X1    g016(.A(G8gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(new_n206_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT14), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT73), .B1(new_n214_), .B2(new_n222_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n213_), .A2(new_n216_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n208_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n216_), .A2(new_n221_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G36gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G29gat), .ZN(new_n231_));
  INV_X1    g030(.A(G29gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G36gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G50gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G43gat), .ZN(new_n236_));
  INV_X1    g035(.A(G43gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G50gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n231_), .A2(new_n233_), .A3(new_n236_), .A4(new_n238_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n229_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT15), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT15), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n245_), .A2(new_n224_), .A3(new_n228_), .A4(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n243_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT77), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n240_), .A2(new_n241_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n224_), .A2(new_n251_), .A3(new_n228_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n251_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n250_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n224_), .A2(new_n251_), .A3(new_n228_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n243_), .A2(KEYINPUT77), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n248_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n249_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n205_), .B1(new_n259_), .B2(KEYINPUT78), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT78), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n248_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n261_), .B(new_n204_), .C1(new_n262_), .C2(new_n249_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n267_), .B1(G155gat), .B2(G162gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(G155gat), .A3(G162gat), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n266_), .A2(new_n268_), .B1(new_n269_), .B2(KEYINPUT85), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n269_), .A2(KEYINPUT85), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G141gat), .ZN(new_n273_));
  INV_X1    g072(.A(G148gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n266_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(KEYINPUT86), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n282_), .B1(KEYINPUT2), .B2(new_n275_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(KEYINPUT3), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT3), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(G141gat), .B2(G148gat), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n284_), .A2(new_n286_), .B1(new_n281_), .B2(KEYINPUT86), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n280_), .B1(new_n283_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n265_), .B1(new_n278_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n287_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n275_), .A2(KEYINPUT2), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n281_), .B2(KEYINPUT86), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n266_), .B(new_n279_), .C1(new_n290_), .C2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n272_), .A2(new_n277_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT87), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(KEYINPUT29), .A3(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT90), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT21), .ZN(new_n300_));
  XOR2_X1   g099(.A(G197gat), .B(G204gat), .Z(new_n301_));
  INV_X1    g100(.A(KEYINPUT91), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n299_), .B(new_n303_), .C1(new_n302_), .C2(new_n301_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n301_), .A2(KEYINPUT89), .ZN(new_n305_));
  INV_X1    g104(.A(G204gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT21), .ZN(new_n308_));
  OAI221_X1 g107(.A(new_n297_), .B1(KEYINPUT21), .B2(new_n301_), .C1(new_n305_), .C2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G228gat), .A2(G233gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n296_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G78gat), .B(G106gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT93), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT94), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(KEYINPUT92), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT92), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n304_), .A2(new_n309_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n293_), .A2(new_n294_), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n316_), .A2(new_n318_), .B1(KEYINPUT29), .B2(new_n319_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n312_), .B(new_n315_), .C1(new_n320_), .C2(new_n311_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT95), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n318_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n317_), .B1(new_n304_), .B2(new_n309_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n278_), .A2(new_n288_), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n324_), .A2(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n311_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n330_), .A2(KEYINPUT95), .A3(new_n312_), .A4(new_n315_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n323_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n289_), .A2(new_n295_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n326_), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G22gat), .B(G50gat), .Z(new_n337_));
  INV_X1    g136(.A(new_n335_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n326_), .A3(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n337_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n338_), .B1(new_n333_), .B2(new_n326_), .ZN(new_n342_));
  AOI211_X1 g141(.A(KEYINPUT29), .B(new_n335_), .C1(new_n289_), .C2(new_n295_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n304_), .A2(new_n309_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n345_), .A2(new_n329_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n328_), .A2(new_n329_), .B1(new_n296_), .B2(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n340_), .B(new_n344_), .C1(new_n347_), .C2(new_n314_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n332_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n330_), .A2(new_n312_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n315_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n352_), .A2(new_n321_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT84), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G113gat), .B(G120gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n355_), .B(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT23), .ZN(new_n360_));
  OR2_X1    g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(KEYINPUT24), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT82), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n360_), .B(new_n364_), .C1(KEYINPUT24), .C2(new_n361_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G183gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT79), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n367_), .A2(KEYINPUT79), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n370_));
  OAI211_X1 g169(.A(KEYINPUT25), .B(new_n368_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n372_));
  OR3_X1    g171(.A1(new_n370_), .A2(new_n367_), .A3(KEYINPUT25), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT26), .B(G190gat), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n361_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT24), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n371_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT81), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n366_), .A2(new_n375_), .A3(new_n378_), .A4(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n369_), .A2(new_n368_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n360_), .B1(new_n382_), .B2(G190gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G169gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G71gat), .B(G99gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT83), .B(G43gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n381_), .A2(new_n386_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n381_), .B2(new_n386_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n358_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n355_), .B(new_n356_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n390_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(new_n209_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT30), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT31), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n393_), .A2(new_n396_), .A3(new_n401_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n349_), .A2(new_n353_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n345_), .A2(new_n381_), .A3(new_n386_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n360_), .B1(G183gat), .B2(G190gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT22), .B(G169gat), .ZN(new_n409_));
  INV_X1    g208(.A(G176gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n376_), .B(KEYINPUT97), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n408_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT98), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n408_), .A2(KEYINPUT98), .A3(new_n411_), .A4(new_n412_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT96), .B(KEYINPUT24), .Z(new_n417_));
  OR2_X1    g216(.A1(new_n417_), .A2(new_n361_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n418_), .A2(new_n360_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT25), .B(G183gat), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n377_), .A2(new_n417_), .B1(new_n374_), .B2(new_n420_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n415_), .A2(new_n416_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n407_), .B(KEYINPUT20), .C1(new_n345_), .C2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT19), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT20), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n381_), .A2(new_n386_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n310_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n425_), .B1(new_n422_), .B2(new_n345_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n423_), .A2(new_n425_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT18), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G64gat), .B(G92gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n432_), .B(new_n433_), .Z(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT32), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT100), .B1(new_n430_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n407_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT20), .B1(new_n422_), .B2(new_n345_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n425_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n428_), .A2(new_n429_), .ZN(new_n440_));
  AND4_X1   g239(.A1(KEYINPUT100), .A2(new_n439_), .A3(new_n440_), .A4(new_n435_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n423_), .A2(new_n425_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n425_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n419_), .A2(new_n421_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n316_), .A2(new_n444_), .A3(new_n413_), .A4(new_n318_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n443_), .B1(new_n428_), .B2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  OAI22_X1  g246(.A1(new_n436_), .A2(new_n441_), .B1(new_n447_), .B2(new_n435_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n289_), .A2(new_n395_), .A3(new_n295_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n358_), .A2(new_n327_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G225gat), .A2(G233gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G1gat), .B(G29gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(G85gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT0), .B(G57gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n455_), .B(new_n456_), .Z(new_n457_));
  INV_X1    g256(.A(KEYINPUT4), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n289_), .A2(new_n395_), .A3(new_n295_), .A4(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT99), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n449_), .A2(KEYINPUT4), .A3(new_n450_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n452_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n453_), .B(new_n457_), .C1(new_n460_), .C2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT101), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT99), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n459_), .B(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n461_), .A2(new_n462_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT101), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n453_), .A4(new_n457_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n465_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT102), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n467_), .A2(new_n468_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n473_), .B1(new_n474_), .B2(new_n457_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n453_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n457_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(KEYINPUT102), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n448_), .B1(new_n472_), .B2(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n439_), .A2(new_n440_), .A3(new_n434_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n434_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n474_), .A2(KEYINPUT33), .A3(new_n457_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT33), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n464_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n457_), .B1(new_n451_), .B2(new_n462_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n461_), .A2(new_n452_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n487_), .B1(new_n460_), .B2(new_n488_), .ZN(new_n489_));
  AND4_X1   g288(.A1(new_n483_), .A2(new_n484_), .A3(new_n486_), .A4(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n406_), .B1(new_n480_), .B2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n403_), .A2(new_n404_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n340_), .A2(new_n344_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n347_), .A2(new_n315_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n321_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n405_), .B(new_n497_), .C1(new_n348_), .C2(new_n332_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n439_), .A2(new_n440_), .A3(new_n434_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT27), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n442_), .A2(new_n446_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n434_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT27), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT103), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  OAI211_X1 g307(.A(KEYINPUT103), .B(new_n505_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n504_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n465_), .A2(new_n471_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n499_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n264_), .B1(new_n491_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G230gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT64), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT10), .B(G99gat), .Z(new_n517_));
  INV_X1    g316(.A(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G85gat), .B(G92gat), .Z(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT9), .ZN(new_n521_));
  INV_X1    g320(.A(G85gat), .ZN(new_n522_));
  INV_X1    g321(.A(G92gat), .ZN(new_n523_));
  OR3_X1    g322(.A1(new_n522_), .A2(new_n523_), .A3(KEYINPUT9), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT6), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(G99gat), .A3(G106gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n519_), .A2(new_n521_), .A3(new_n524_), .A4(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(G99gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(new_n518_), .A3(KEYINPUT65), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT7), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT7), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n534_), .A2(new_n531_), .A3(new_n518_), .A4(KEYINPUT65), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n529_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT8), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n536_), .A2(new_n520_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n538_), .B1(new_n536_), .B2(new_n520_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n530_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542_));
  NOR2_X1   g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n545_), .B2(KEYINPUT11), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT67), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n545_), .B2(KEYINPUT11), .ZN(new_n548_));
  INV_X1    g347(.A(G64gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(G57gat), .ZN(new_n550_));
  INV_X1    g349(.A(G57gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(G64gat), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n550_), .A2(new_n552_), .A3(new_n547_), .A4(KEYINPUT11), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n546_), .B1(new_n548_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n550_), .A2(new_n552_), .A3(KEYINPUT11), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT67), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(new_n552_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT11), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n557_), .A2(new_n560_), .A3(new_n544_), .A4(new_n553_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n541_), .A2(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n562_), .B(new_n530_), .C1(new_n540_), .C2(new_n539_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(KEYINPUT12), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT12), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n541_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n516_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n516_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G120gat), .B(G148gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n569_), .A2(new_n571_), .A3(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n577_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT13), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT70), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT34), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n245_), .A2(new_n246_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n541_), .A2(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n242_), .B(new_n530_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n592_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n593_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n541_), .A2(new_n246_), .A3(new_n245_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n593_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n597_), .A4(new_n596_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n588_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT71), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT37), .B1(new_n603_), .B2(new_n604_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n599_), .A2(new_n586_), .A3(new_n602_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT69), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT69), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n599_), .A2(new_n610_), .A3(new_n602_), .A4(new_n586_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n599_), .A2(new_n602_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT72), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n599_), .A2(KEYINPUT72), .A3(new_n602_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n588_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n612_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT37), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n607_), .A2(new_n612_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(G231gat), .ZN(new_n622_));
  INV_X1    g421(.A(G233gat), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n229_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n229_), .A2(new_n624_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n562_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n563_), .A3(new_n626_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(G127gat), .B(G155gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT16), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT17), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n630_), .A2(KEYINPUT75), .A3(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n628_), .A2(new_n636_), .A3(new_n629_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT75), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n634_), .B(new_n635_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n630_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n641_), .A2(KEYINPUT76), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT76), .B1(new_n641_), .B2(new_n644_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n581_), .A2(new_n621_), .A3(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n514_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n512_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n217_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n647_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n619_), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n654_), .B(new_n655_), .C1(new_n491_), .C2(new_n513_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n581_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n264_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n512_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n651_), .A2(new_n652_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n653_), .A2(new_n660_), .A3(new_n661_), .ZN(G1324gat));
  INV_X1    g461(.A(new_n510_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n649_), .A2(new_n218_), .A3(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G8gat), .B1(new_n659_), .B2(new_n510_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n664_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT40), .B(new_n664_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n659_), .B2(new_n492_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT41), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n649_), .A2(new_n209_), .A3(new_n405_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n349_), .A2(new_n353_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G22gat), .B1(new_n659_), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT42), .ZN(new_n679_));
  INV_X1    g478(.A(new_n677_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n649_), .A2(new_n211_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1327gat));
  NOR3_X1   g481(.A1(new_n657_), .A2(new_n264_), .A3(new_n647_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n491_), .A2(new_n513_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n621_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT43), .B(new_n621_), .C1(new_n491_), .C2(new_n513_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n683_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT44), .B(new_n683_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n650_), .A3(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(KEYINPUT104), .ZN(new_n694_));
  OAI21_X1  g493(.A(G29gat), .B1(new_n693_), .B2(KEYINPUT104), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n654_), .A2(new_n655_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(new_n657_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n514_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT105), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n514_), .A2(new_n700_), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n650_), .A2(new_n232_), .ZN(new_n703_));
  OAI22_X1  g502(.A1(new_n694_), .A2(new_n695_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  NAND3_X1  g503(.A1(new_n691_), .A2(new_n663_), .A3(new_n692_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n510_), .A2(G36gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n699_), .A2(new_n701_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT45), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n699_), .A2(new_n710_), .A3(new_n701_), .A4(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n706_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n706_), .A2(KEYINPUT46), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND3_X1  g516(.A1(new_n691_), .A2(new_n405_), .A3(new_n692_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G43gat), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n699_), .A2(new_n237_), .A3(new_n405_), .A4(new_n701_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1330gat));
  NAND4_X1  g525(.A1(new_n691_), .A2(G50gat), .A3(new_n680_), .A4(new_n692_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n235_), .B1(new_n702_), .B2(new_n677_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1331gat));
  INV_X1    g528(.A(new_n264_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n581_), .A2(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n685_), .A2(new_n731_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n732_), .A2(new_n647_), .A3(new_n621_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n551_), .A3(new_n650_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n656_), .A2(new_n731_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(new_n650_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n736_), .B2(new_n551_), .ZN(G1332gat));
  AOI21_X1  g536(.A(new_n549_), .B1(new_n735_), .B2(new_n663_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT48), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n733_), .A2(new_n549_), .A3(new_n663_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1333gat));
  INV_X1    g540(.A(G71gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n735_), .B2(new_n405_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT49), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n733_), .A2(new_n742_), .A3(new_n405_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1334gat));
  INV_X1    g545(.A(G78gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n735_), .B2(new_n680_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n733_), .A2(new_n747_), .A3(new_n680_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1335gat));
  INV_X1    g551(.A(new_n696_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n732_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n522_), .A3(new_n650_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n581_), .A2(new_n647_), .A3(new_n730_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n756_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT108), .B(new_n756_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n512_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n755_), .B1(new_n761_), .B2(new_n522_), .ZN(G1336gat));
  NAND3_X1  g561(.A1(new_n754_), .A2(new_n523_), .A3(new_n663_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n510_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n523_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT109), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n763_), .C1(new_n764_), .C2(new_n523_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1337gat));
  NAND3_X1  g568(.A1(new_n754_), .A2(new_n405_), .A3(new_n517_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n492_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n531_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT51), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n770_), .C1(new_n771_), .C2(new_n531_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1338gat));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n518_), .B1(new_n777_), .B2(KEYINPUT52), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n757_), .B2(new_n677_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(KEYINPUT111), .A3(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n732_), .A2(new_n518_), .A3(new_n680_), .A4(new_n753_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT110), .ZN(new_n783_));
  OAI221_X1 g582(.A(new_n778_), .B1(new_n777_), .B2(KEYINPUT52), .C1(new_n757_), .C2(new_n677_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n781_), .A2(new_n783_), .A3(new_n784_), .A4(new_n786_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1339gat));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n648_), .A2(KEYINPUT113), .A3(new_n791_), .A4(new_n264_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n621_), .A2(new_n581_), .A3(new_n647_), .A4(new_n264_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(KEYINPUT54), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(KEYINPUT54), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n792_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n569_), .A2(new_n571_), .A3(new_n577_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n264_), .B2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n578_), .A2(KEYINPUT114), .A3(new_n263_), .A4(new_n260_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n566_), .A2(new_n568_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n570_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n569_), .A2(KEYINPUT55), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT115), .B1(new_n803_), .B2(new_n570_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n566_), .A2(new_n809_), .A3(new_n516_), .A4(new_n568_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .A4(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n577_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n577_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n802_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n258_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n243_), .A2(new_n247_), .A3(new_n258_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n205_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n204_), .B1(new_n262_), .B2(new_n249_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n580_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n619_), .B1(new_n816_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n799_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n577_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n577_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n621_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT58), .B(new_n826_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n824_), .A2(new_n825_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n827_), .A2(new_n828_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n822_), .B1(new_n834_), .B2(new_n802_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(KEYINPUT57), .A3(new_n619_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n797_), .B1(new_n654_), .B2(new_n837_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n663_), .A2(new_n512_), .A3(new_n498_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n829_), .A2(new_n830_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n843_), .A2(new_n832_), .A3(new_n686_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT57), .B1(new_n835_), .B2(new_n619_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT117), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n824_), .A2(new_n825_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n831_), .A2(new_n832_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n846_), .A2(new_n836_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n797_), .B1(new_n851_), .B2(new_n654_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n839_), .A2(KEYINPUT116), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n839_), .A2(KEYINPUT116), .ZN(new_n854_));
  OR3_X1    g653(.A1(new_n853_), .A2(new_n854_), .A3(KEYINPUT59), .ZN(new_n855_));
  OAI22_X1  g654(.A1(new_n841_), .A2(new_n842_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n264_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n841_), .ZN(new_n858_));
  OR3_X1    g657(.A1(new_n858_), .A2(G113gat), .A3(new_n264_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1340gat));
  XOR2_X1   g659(.A(KEYINPUT118), .B(G120gat), .Z(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n856_), .B2(new_n581_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n657_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT119), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n841_), .B(new_n865_), .C1(new_n864_), .C2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n862_), .A2(new_n868_), .ZN(G1341gat));
  OAI21_X1  g668(.A(G127gat), .B1(new_n856_), .B2(new_n654_), .ZN(new_n870_));
  OR3_X1    g669(.A1(new_n858_), .A2(G127gat), .A3(new_n654_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1342gat));
  AOI21_X1  g671(.A(G134gat), .B1(new_n841_), .B2(new_n655_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n856_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n686_), .A2(G134gat), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT120), .Z(new_n876_));
  AOI21_X1  g675(.A(new_n873_), .B1(new_n874_), .B2(new_n876_), .ZN(G1343gat));
  NAND2_X1  g676(.A1(new_n837_), .A2(new_n654_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n797_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n493_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n880_), .A2(new_n510_), .A3(new_n650_), .A4(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n264_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n273_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n581_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n274_), .ZN(G1345gat));
  NOR2_X1   g685(.A1(new_n882_), .A2(new_n654_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT61), .B(G155gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n882_), .B2(new_n621_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n619_), .A2(G162gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n882_), .B2(new_n891_), .ZN(G1347gat));
  NOR3_X1   g691(.A1(new_n650_), .A2(new_n510_), .A3(new_n492_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n677_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT121), .B1(new_n852_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896_));
  INV_X1    g695(.A(new_n894_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n836_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n847_), .A2(new_n849_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(KEYINPUT117), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n647_), .B1(new_n900_), .B2(new_n850_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n896_), .B(new_n897_), .C1(new_n901_), .C2(new_n797_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n895_), .A2(new_n902_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n730_), .A2(new_n409_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n836_), .B1(new_n833_), .B2(new_n848_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n844_), .A2(new_n845_), .A3(KEYINPUT117), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n654_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n879_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n730_), .A3(new_n897_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n910_), .A2(new_n911_), .A3(G169gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n910_), .B2(G169gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n905_), .B1(new_n912_), .B2(new_n913_), .ZN(G1348gat));
  NOR2_X1   g713(.A1(new_n838_), .A2(new_n680_), .ZN(new_n915_));
  AND4_X1   g714(.A1(G176gat), .A2(new_n915_), .A3(new_n657_), .A4(new_n893_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n896_), .B1(new_n909_), .B2(new_n897_), .ZN(new_n917_));
  AOI211_X1 g716(.A(KEYINPUT121), .B(new_n894_), .C1(new_n908_), .C2(new_n879_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n657_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n916_), .B1(new_n919_), .B2(new_n410_), .ZN(G1349gat));
  AND2_X1   g719(.A1(new_n893_), .A2(new_n647_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n382_), .B1(new_n915_), .B2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n654_), .A2(new_n420_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n903_), .B2(new_n923_), .ZN(G1350gat));
  AND2_X1   g723(.A1(new_n655_), .A2(new_n374_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n903_), .A2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(G190gat), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n621_), .B1(new_n895_), .B2(new_n902_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(G1351gat));
  XNOR2_X1  g728(.A(KEYINPUT123), .B(G197gat), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n650_), .A2(new_n510_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n881_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n838_), .B2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n933_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n880_), .A2(KEYINPUT122), .A3(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n930_), .B1(new_n937_), .B2(new_n730_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(G197gat), .ZN(new_n940_));
  AOI211_X1 g739(.A(new_n264_), .B(new_n940_), .C1(new_n934_), .C2(new_n936_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n938_), .A2(new_n941_), .ZN(G1352gat));
  AND2_X1   g741(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n943_));
  NOR2_X1   g742(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n944_));
  OAI211_X1 g743(.A(new_n937_), .B(new_n657_), .C1(new_n943_), .C2(new_n944_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n581_), .B1(new_n934_), .B2(new_n936_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(new_n944_), .ZN(G1353gat));
  NOR2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n948_), .A2(KEYINPUT125), .ZN(new_n949_));
  AOI211_X1 g748(.A(new_n949_), .B(new_n654_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(new_n934_), .B2(new_n936_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n948_), .A2(KEYINPUT125), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(KEYINPUT126), .ZN(new_n954_));
  INV_X1    g753(.A(new_n954_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n952_), .B(new_n955_), .ZN(G1354gat));
  NAND2_X1  g755(.A1(new_n937_), .A2(new_n655_), .ZN(new_n957_));
  INV_X1    g756(.A(G218gat), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n621_), .A2(new_n958_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(KEYINPUT127), .ZN(new_n960_));
  AOI22_X1  g759(.A1(new_n957_), .A2(new_n958_), .B1(new_n937_), .B2(new_n960_), .ZN(G1355gat));
endmodule


