//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT81), .B1(new_n203_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT81), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(new_n202_), .B2(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT76), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G183gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OAI22_X1  g012(.A1(new_n206_), .A2(new_n208_), .B1(G190gat), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT22), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n217_));
  AOI21_X1  g016(.A(G176gat), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT22), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G169gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n218_), .B1(new_n222_), .B2(new_n217_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n214_), .A2(new_n223_), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n232_));
  INV_X1    g031(.A(G190gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT77), .B1(new_n233_), .B2(KEYINPUT26), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT77), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(G190gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(KEYINPUT26), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G183gat), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n234_), .A2(new_n237_), .A3(new_n238_), .A4(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n210_), .A2(new_n212_), .A3(KEYINPUT25), .ZN(new_n242_));
  OAI211_X1 g041(.A(KEYINPUT79), .B(new_n232_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n204_), .B1(G183gat), .B2(G190gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NOR3_X1   g045(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n210_), .A2(new_n212_), .A3(KEYINPUT25), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n239_), .A2(G183gat), .B1(new_n233_), .B2(KEYINPUT26), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n250_), .A2(new_n237_), .A3(new_n234_), .A4(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT79), .B1(new_n252_), .B2(new_n232_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n229_), .B1(new_n249_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT30), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT82), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G71gat), .B(G99gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(G43gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260_));
  INV_X1    g059(.A(G15gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n259_), .B(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n256_), .A2(KEYINPUT82), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n263_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G113gat), .B(G120gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT31), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n265_), .A2(new_n267_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT27), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G226gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G218gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(G211gat), .ZN(new_n280_));
  INV_X1    g079(.A(G211gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G218gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n284_));
  INV_X1    g083(.A(G204gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT21), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(G197gat), .B2(G204gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n283_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G197gat), .A2(G204gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT85), .B(G197gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(G204gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n290_), .B1(new_n293_), .B2(KEYINPUT21), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n288_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT86), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(KEYINPUT85), .A2(G197gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(G204gat), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n291_), .ZN(new_n300_));
  AND4_X1   g099(.A1(KEYINPUT86), .A2(new_n295_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n294_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n254_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n247_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n224_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n304_), .B1(new_n230_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n206_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n208_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n209_), .A2(KEYINPUT25), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n240_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n236_), .A2(G190gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT88), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n238_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n313_), .B2(new_n238_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n312_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n246_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G176gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n216_), .A2(new_n220_), .A3(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n228_), .A2(new_n322_), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n309_), .A2(new_n318_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n295_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n293_), .A2(KEYINPUT86), .A3(new_n295_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n299_), .A2(new_n300_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n288_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n327_), .A2(new_n328_), .B1(new_n330_), .B2(new_n290_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT20), .B1(new_n324_), .B2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n278_), .B1(new_n303_), .B2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G8gat), .B(G36gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n254_), .A2(new_n302_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT20), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n324_), .B2(new_n331_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n278_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n333_), .A2(new_n338_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n338_), .B1(new_n333_), .B2(new_n343_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n344_), .B1(new_n345_), .B2(KEYINPUT90), .ZN(new_n346_));
  INV_X1    g145(.A(new_n338_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n232_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n331_), .B1(new_n351_), .B2(new_n229_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n228_), .B(new_n322_), .C1(new_n246_), .C2(new_n319_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n313_), .A2(new_n238_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT88), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n311_), .B1(new_n355_), .B2(new_n315_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n247_), .B1(new_n231_), .B2(new_n224_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n353_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT20), .B1(new_n302_), .B2(new_n359_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n352_), .A2(new_n360_), .A3(new_n278_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n351_), .A2(new_n331_), .A3(new_n229_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n340_), .B1(new_n302_), .B2(new_n359_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n342_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(KEYINPUT90), .B(new_n347_), .C1(new_n361_), .C2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n275_), .B1(new_n346_), .B2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n361_), .A2(new_n364_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n275_), .B1(new_n368_), .B2(new_n338_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT94), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n278_), .B1(new_n352_), .B2(new_n360_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n363_), .A3(new_n342_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n370_), .B1(new_n373_), .B2(new_n347_), .ZN(new_n374_));
  AOI211_X1 g173(.A(KEYINPUT94), .B(new_n338_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n369_), .B(KEYINPUT95), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n367_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(new_n347_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT94), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n373_), .A2(new_n370_), .A3(new_n347_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT95), .B1(new_n381_), .B2(new_n369_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT83), .B1(new_n384_), .B2(KEYINPUT1), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT1), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(G155gat), .A4(G162gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(KEYINPUT1), .ZN(new_n389_));
  OR2_X1    g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n385_), .A2(new_n388_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G141gat), .B(G148gat), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394_));
  INV_X1    g193(.A(G141gat), .ZN(new_n395_));
  INV_X1    g194(.A(G148gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n397_), .A2(new_n399_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n390_), .A2(new_n384_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n393_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n270_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n268_), .B(new_n269_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n393_), .A3(new_n404_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(KEYINPUT4), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n405_), .A2(new_n270_), .A3(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n409_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n406_), .A2(new_n410_), .A3(new_n408_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT92), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n406_), .A2(new_n417_), .A3(new_n410_), .A4(new_n408_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n419_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n414_), .A2(new_n416_), .A3(new_n424_), .A4(new_n418_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G106gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n405_), .A2(KEYINPUT29), .ZN(new_n431_));
  INV_X1    g230(.A(G78gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n302_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n432_), .B1(new_n302_), .B2(new_n431_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n430_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n435_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(G106gat), .A3(new_n433_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G22gat), .B(G50gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n405_), .A2(KEYINPUT29), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT28), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n302_), .A2(new_n444_), .B1(G228gat), .B2(G233gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n443_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n440_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n436_), .A2(new_n438_), .A3(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n441_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n446_), .B1(new_n441_), .B2(new_n448_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n274_), .A2(new_n383_), .A3(new_n429_), .A4(new_n451_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n449_), .A2(new_n450_), .A3(new_n428_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n347_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT90), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(new_n344_), .A3(new_n365_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n409_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n406_), .A2(new_n411_), .A3(new_n408_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n425_), .A2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT33), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n427_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(new_n427_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT93), .B1(new_n457_), .B2(new_n464_), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n361_), .A2(new_n364_), .A3(new_n347_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n466_), .B1(new_n455_), .B2(new_n454_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n427_), .A2(new_n463_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n427_), .B2(new_n461_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n470_), .A4(new_n365_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n338_), .A2(KEYINPUT32), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n373_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n368_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n428_), .B(new_n473_), .C1(new_n474_), .C2(new_n472_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n465_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n453_), .A2(new_n383_), .B1(new_n476_), .B2(new_n451_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n452_), .B1(new_n477_), .B2(new_n274_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G8gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT74), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G22gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n261_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G15gat), .A2(G22gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G1gat), .A2(G8gat), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n483_), .A2(new_n484_), .B1(KEYINPUT14), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n481_), .B(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G29gat), .B(G36gat), .Z(new_n488_));
  XOR2_X1   g287(.A(G43gat), .B(G50gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n487_), .B(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n487_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n490_), .B(KEYINPUT15), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n493_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n491_), .A2(new_n493_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G113gat), .B(G141gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(G169gat), .B(G197gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n498_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n501_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n502_), .A2(KEYINPUT75), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT75), .B1(new_n502_), .B2(new_n503_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n478_), .A2(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n508_), .A2(KEYINPUT96), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G85gat), .B(G92gat), .Z(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT10), .B(G99gat), .Z(new_n514_));
  AOI22_X1  g313(.A1(KEYINPUT9), .A2(new_n513_), .B1(new_n514_), .B2(new_n430_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT64), .B(G92gat), .Z(new_n516_));
  INV_X1    g315(.A(KEYINPUT9), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(G85gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n512_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT70), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n512_), .A2(new_n515_), .A3(KEYINPUT70), .A4(new_n518_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT66), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n524_), .A2(G99gat), .A3(G106gat), .ZN(new_n525_));
  INV_X1    g324(.A(G99gat), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(new_n430_), .C1(new_n523_), .C2(KEYINPUT66), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n512_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT8), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n513_), .A2(KEYINPUT67), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n530_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n521_), .B(new_n522_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n495_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n519_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n529_), .A2(new_n531_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT8), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n539_), .B2(new_n532_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n490_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT34), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n536_), .A2(new_n541_), .A3(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n544_), .A2(new_n545_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(new_n548_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G134gat), .B(G162gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT36), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n554_), .B(KEYINPUT36), .Z(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(KEYINPUT73), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT37), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n559_), .A2(new_n561_), .A3(KEYINPUT37), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G71gat), .B(G78gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT68), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n567_), .B1(new_n570_), .B2(KEYINPUT11), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n571_), .B1(KEYINPUT11), .B2(new_n570_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(KEYINPUT11), .A3(new_n567_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n494_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578_));
  XOR2_X1   g377(.A(G127gat), .B(G155gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT16), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  OR3_X1    g381(.A1(new_n577_), .A2(new_n578_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(KEYINPUT17), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n566_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n519_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n572_), .A2(new_n573_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n540_), .A2(new_n574_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n588_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT69), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n572_), .A2(KEYINPUT12), .A3(new_n573_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n535_), .A2(new_n596_), .B1(new_n540_), .B2(new_n574_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT12), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n540_), .B2(new_n574_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n588_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n593_), .A2(new_n594_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n595_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(G120gat), .B(G148gat), .Z(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT72), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n602_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT13), .ZN(new_n611_));
  INV_X1    g410(.A(new_n607_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n595_), .A2(new_n612_), .A3(new_n600_), .A4(new_n601_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n610_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n611_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n508_), .B2(KEYINPUT96), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n509_), .A2(new_n587_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n429_), .A2(G1gat), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n623_), .A2(KEYINPUT38), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n621_), .A2(KEYINPUT38), .A3(new_n622_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n586_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n626_), .B(new_n507_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT98), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n476_), .A2(new_n451_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n382_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n630_), .A2(new_n453_), .A3(new_n367_), .A4(new_n376_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n272_), .A2(new_n273_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n630_), .A2(new_n451_), .A3(new_n367_), .A4(new_n376_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(new_n428_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n632_), .A2(new_n633_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n560_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n628_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n639_), .B2(new_n429_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n624_), .A2(new_n625_), .A3(new_n640_), .ZN(G1324gat));
  INV_X1    g440(.A(G8gat), .ZN(new_n642_));
  INV_X1    g441(.A(new_n383_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n621_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n628_), .A2(new_n643_), .A3(new_n638_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n645_), .A2(new_n646_), .A3(G8gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n645_), .B2(G8gat), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n644_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(G1325gat));
  NAND3_X1  g453(.A1(new_n621_), .A2(new_n261_), .A3(new_n274_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G15gat), .B1(new_n639_), .B2(new_n633_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT41), .Z(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1326gat));
  INV_X1    g457(.A(new_n451_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n621_), .A2(new_n482_), .A3(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G22gat), .B1(new_n639_), .B2(new_n451_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT42), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1327gat));
  NOR2_X1   g462(.A1(new_n626_), .A2(new_n559_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n509_), .A2(new_n618_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n666_), .B2(new_n428_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n616_), .A2(new_n586_), .A3(new_n507_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n565_), .B1(new_n478_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n637_), .A2(KEYINPUT101), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n563_), .A2(new_n670_), .A3(new_n564_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n637_), .B2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n478_), .A2(new_n566_), .A3(KEYINPUT102), .A4(new_n670_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n669_), .B1(new_n674_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT44), .B(new_n669_), .C1(new_n674_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n428_), .A2(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n667_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  OR2_X1    g486(.A1(new_n383_), .A2(G36gat), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n665_), .A2(new_n688_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT45), .Z(new_n690_));
  NAND3_X1  g489(.A1(new_n682_), .A2(new_n643_), .A3(new_n683_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n691_), .A2(new_n692_), .A3(G36gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n691_), .B2(G36gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT46), .B(new_n690_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1329gat));
  AOI21_X1  g498(.A(G43gat), .B1(new_n666_), .B2(new_n274_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT104), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n685_), .A2(G43gat), .A3(new_n274_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT47), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n701_), .A2(new_n705_), .A3(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1330gat));
  AOI21_X1  g506(.A(G50gat), .B1(new_n666_), .B2(new_n659_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n659_), .A2(G50gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n685_), .B2(new_n709_), .ZN(G1331gat));
  NOR3_X1   g509(.A1(new_n637_), .A2(new_n507_), .A3(new_n616_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n587_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT105), .Z(new_n713_));
  AOI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n428_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n616_), .A2(new_n586_), .A3(new_n507_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n638_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(G57gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n428_), .B2(KEYINPUT106), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(KEYINPUT106), .B2(new_n718_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n714_), .B1(new_n717_), .B2(new_n720_), .ZN(G1332gat));
  INV_X1    g520(.A(G64gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n713_), .A2(new_n722_), .A3(new_n643_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G64gat), .B1(new_n716_), .B2(new_n383_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT48), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1333gat));
  INV_X1    g525(.A(G71gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n713_), .A2(new_n727_), .A3(new_n274_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G71gat), .B1(new_n716_), .B2(new_n633_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT49), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1334gat));
  NAND3_X1  g530(.A1(new_n713_), .A2(new_n432_), .A3(new_n659_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G78gat), .B1(new_n716_), .B2(new_n451_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT50), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1335gat));
  INV_X1    g534(.A(G85gat), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n616_), .A2(new_n626_), .A3(new_n507_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n672_), .A2(new_n673_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT43), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n677_), .A2(new_n678_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(KEYINPUT108), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n674_), .B2(new_n679_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n738_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n736_), .B1(new_n745_), .B2(new_n428_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n711_), .A2(new_n664_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT107), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n748_), .A2(G85gat), .A3(new_n429_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n746_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(G1336gat));
  INV_X1    g551(.A(new_n748_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G92gat), .B1(new_n753_), .B2(new_n643_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n643_), .A2(new_n516_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n745_), .B2(new_n755_), .ZN(G1337gat));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT51), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n274_), .A2(new_n514_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n748_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n745_), .A2(new_n274_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(G99gat), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n757_), .A2(KEYINPUT51), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(G1338gat));
  NAND2_X1  g563(.A1(new_n737_), .A2(new_n659_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n766_));
  OR3_X1    g565(.A1(new_n766_), .A2(KEYINPUT111), .A3(new_n430_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT111), .B1(new_n766_), .B2(new_n430_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(KEYINPUT52), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n451_), .A2(G106gat), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n753_), .A2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n768_), .B2(KEYINPUT52), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT53), .B1(new_n770_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n773_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n769_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(G1339gat));
  AND2_X1   g577(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n779_));
  NOR2_X1   g578(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n507_), .A2(new_n586_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT112), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n565_), .B1(new_n783_), .B2(KEYINPUT112), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n781_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n783_), .A2(KEYINPUT112), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n788_), .A2(new_n784_), .A3(new_n565_), .A4(new_n779_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n588_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n600_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n597_), .A2(KEYINPUT55), .A3(new_n588_), .A4(new_n599_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n609_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT56), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n501_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n492_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n496_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n503_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n608_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n797_), .A2(new_n613_), .A3(new_n803_), .A4(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT58), .B1(new_n807_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n613_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n812_));
  AOI211_X1 g611(.A(KEYINPUT56), .B(new_n608_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n812_), .A2(new_n802_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT114), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n565_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n809_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n808_), .B1(new_n814_), .B2(KEYINPUT114), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n807_), .A2(new_n810_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n566_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT115), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n822_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n812_), .A2(new_n506_), .A3(new_n813_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n802_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n559_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT57), .B(new_n559_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n823_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n790_), .B1(new_n832_), .B2(new_n586_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n635_), .A2(new_n428_), .A3(new_n274_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT116), .Z(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(G113gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n507_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n790_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n830_), .B1(new_n818_), .B2(new_n822_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n626_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(KEYINPUT59), .A3(new_n835_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n506_), .B1(new_n841_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n839_), .B1(new_n846_), .B2(new_n838_), .ZN(G1340gat));
  NOR2_X1   g646(.A1(new_n616_), .A2(KEYINPUT60), .ZN(new_n848_));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  MUX2_X1   g648(.A(KEYINPUT60), .B(new_n848_), .S(new_n849_), .Z(new_n850_));
  NAND2_X1  g649(.A1(new_n837_), .A2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n851_), .A2(KEYINPUT117), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(KEYINPUT117), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n616_), .B1(new_n841_), .B2(new_n845_), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n852_), .A2(new_n853_), .B1(new_n849_), .B2(new_n854_), .ZN(G1341gat));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n626_), .A2(G127gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT118), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n841_), .B2(new_n845_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n844_), .A2(new_n626_), .A3(new_n835_), .ZN(new_n861_));
  INV_X1    g660(.A(G127gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n856_), .B1(new_n860_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n845_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT59), .B1(new_n844_), .B2(new_n835_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n858_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n868_), .A2(KEYINPUT119), .A3(new_n863_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n865_), .A2(new_n869_), .ZN(G1342gat));
  NAND2_X1  g669(.A1(new_n566_), .A2(G134gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT121), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n841_), .B2(new_n845_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n833_), .A2(new_n559_), .A3(new_n836_), .ZN(new_n874_));
  OR3_X1    g673(.A1(new_n874_), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT120), .B1(new_n874_), .B2(G134gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n873_), .B1(new_n875_), .B2(new_n876_), .ZN(G1343gat));
  NAND3_X1  g676(.A1(new_n633_), .A2(new_n659_), .A3(new_n428_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n833_), .A2(new_n643_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n507_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n617_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n626_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  INV_X1    g685(.A(G162gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n879_), .A2(new_n887_), .A3(new_n560_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n879_), .A2(new_n566_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n887_), .ZN(G1347gat));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n636_), .A2(new_n451_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n844_), .A2(new_n507_), .A3(new_n643_), .A4(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n894_), .A2(new_n895_), .A3(G169gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n894_), .B2(G169gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n891_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n894_), .A2(G169gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT122), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n894_), .A2(new_n895_), .A3(G169gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n900_), .A2(KEYINPUT62), .A3(new_n901_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n894_), .A2(new_n221_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n898_), .A2(new_n902_), .A3(new_n903_), .ZN(G1348gat));
  NOR3_X1   g703(.A1(new_n833_), .A2(new_n383_), .A3(new_n892_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n617_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g706(.A1(new_n844_), .A2(new_n626_), .A3(new_n643_), .A4(new_n893_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n909_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n910_), .A2(new_n911_), .A3(new_n213_), .ZN(new_n912_));
  OR3_X1    g711(.A1(new_n908_), .A2(KEYINPUT123), .A3(new_n312_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT123), .B1(new_n908_), .B2(new_n312_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n912_), .A2(new_n915_), .ZN(G1350gat));
  INV_X1    g715(.A(new_n905_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G190gat), .B1(new_n917_), .B2(new_n565_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n560_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n917_), .B2(new_n919_), .ZN(G1351gat));
  NAND2_X1  g719(.A1(new_n633_), .A2(new_n453_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n833_), .A2(new_n383_), .A3(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n507_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n617_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g725(.A(new_n921_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n844_), .A2(new_n626_), .A3(new_n643_), .A4(new_n927_), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT63), .B(G211gat), .Z(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(KEYINPUT125), .B1(new_n928_), .B2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n928_), .A2(new_n932_), .A3(new_n281_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n928_), .A2(KEYINPUT125), .A3(new_n930_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1354gat));
  XNOR2_X1  g735(.A(KEYINPUT127), .B(G218gat), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n565_), .A2(new_n937_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n922_), .A2(new_n938_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n844_), .A2(new_n560_), .A3(new_n643_), .A4(new_n927_), .ZN(new_n940_));
  XOR2_X1   g739(.A(new_n940_), .B(KEYINPUT126), .Z(new_n941_));
  AOI21_X1  g740(.A(new_n939_), .B1(new_n941_), .B2(new_n937_), .ZN(G1355gat));
endmodule


