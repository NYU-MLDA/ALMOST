//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n913_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT96), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT21), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n203_), .A2(KEYINPUT96), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n208_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n207_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n206_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT95), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n209_), .B1(new_n212_), .B2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT90), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT24), .A3(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n217_), .B(KEYINPUT90), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT23), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT26), .B(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT25), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT89), .B1(new_n228_), .B2(G183gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT25), .B(G183gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n227_), .B(new_n229_), .C1(new_n230_), .C2(KEYINPUT89), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n221_), .A2(new_n224_), .A3(new_n226_), .A4(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n226_), .B1(G183gat), .B2(G190gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT22), .B(G169gat), .Z(new_n234_));
  INV_X1    g033(.A(KEYINPUT91), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G169gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(KEYINPUT22), .B2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n238_), .A2(G176gat), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n233_), .B(new_n220_), .C1(new_n236_), .C2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n216_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT20), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G226gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT19), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n233_), .B(new_n220_), .C1(G176gat), .C2(new_n234_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n227_), .B(KEYINPUT100), .ZN(new_n248_));
  INV_X1    g047(.A(new_n230_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n221_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n247_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n246_), .B1(new_n252_), .B2(new_n216_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n243_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n216_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n213_), .B(KEYINPUT95), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n211_), .A3(new_n210_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n257_), .A2(new_n209_), .A3(new_n232_), .A4(new_n240_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n258_), .A3(KEYINPUT20), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n245_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT101), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n259_), .A2(KEYINPUT101), .A3(new_n245_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n254_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G8gat), .B(G36gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n264_), .A2(new_n270_), .ZN(new_n271_));
  AOI211_X1 g070(.A(new_n269_), .B(new_n254_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n202_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT105), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n252_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n216_), .A2(KEYINPUT97), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT97), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n257_), .A2(new_n277_), .A3(new_n209_), .ZN(new_n278_));
  OAI211_X1 g077(.A(KEYINPUT105), .B(new_n247_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n275_), .A2(new_n276_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n242_), .A2(KEYINPUT20), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n246_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n259_), .A2(new_n245_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n269_), .B(KEYINPUT107), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n202_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n264_), .A2(new_n270_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n273_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n276_), .A2(new_n278_), .ZN(new_n290_));
  INV_X1    g089(.A(G155gat), .ZN(new_n291_));
  INV_X1    g090(.A(G162gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT3), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT92), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301_));
  INV_X1    g100(.A(G141gat), .ZN(new_n302_));
  INV_X1    g101(.A(G148gat), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n300_), .B(new_n301_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n302_), .A2(new_n303_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT2), .B1(new_n305_), .B2(KEYINPUT92), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n299_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT93), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT93), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n299_), .A2(new_n309_), .A3(new_n306_), .A4(new_n304_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n297_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n296_), .B1(new_n294_), .B2(KEYINPUT1), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n293_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n315_), .A2(new_n305_), .A3(new_n298_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT29), .B1(new_n311_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n290_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G228gat), .ZN(new_n319_));
  INV_X1    g118(.A(G233gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT98), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT98), .ZN(new_n323_));
  INV_X1    g122(.A(new_n321_), .ZN(new_n324_));
  AOI211_X1 g123(.A(new_n323_), .B(new_n324_), .C1(new_n290_), .C2(new_n317_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n317_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n216_), .A2(new_n324_), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n322_), .A2(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G22gat), .B(G50gat), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n311_), .A2(new_n316_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR4_X1   g135(.A1(new_n311_), .A2(new_n316_), .A3(KEYINPUT29), .A4(new_n329_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G78gat), .B(G106gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT99), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n335_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n339_), .A2(new_n342_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n340_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n328_), .B(new_n343_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n326_), .A2(new_n327_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n318_), .A2(new_n321_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n323_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n318_), .A2(KEYINPUT98), .A3(new_n321_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n347_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n339_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n345_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n346_), .A2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n289_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G127gat), .B(G134gat), .Z(new_n357_));
  XOR2_X1   g156(.A(G113gat), .B(G120gat), .Z(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n331_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n359_), .B1(new_n311_), .B2(new_n316_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(KEYINPUT4), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n362_), .A2(KEYINPUT4), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(G85gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT0), .B(G57gat), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n370_), .B(new_n371_), .Z(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n367_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n368_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n366_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n372_), .B1(new_n377_), .B2(new_n374_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G43gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n241_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(new_n359_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(G15gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT30), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT31), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n384_), .A2(new_n389_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n380_), .A2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n356_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n254_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n263_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT101), .B1(new_n259_), .B2(new_n245_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n269_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n287_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n401_), .A2(new_n202_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n402_), .A2(new_n355_), .A3(KEYINPUT108), .A4(new_n379_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT108), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n379_), .A2(new_n346_), .A3(new_n354_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n404_), .B1(new_n289_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT103), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n378_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n378_), .B2(new_n408_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n361_), .A2(new_n362_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT104), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n361_), .A2(new_n362_), .A3(KEYINPUT104), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n367_), .A3(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n416_), .B(new_n373_), .C1(new_n367_), .C2(new_n365_), .ZN(new_n417_));
  OAI211_X1 g216(.A(KEYINPUT33), .B(new_n372_), .C1(new_n377_), .C2(new_n374_), .ZN(new_n418_));
  AND4_X1   g217(.A1(new_n287_), .A2(new_n400_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n421_), .B(KEYINPUT106), .Z(new_n422_));
  INV_X1    g221(.A(new_n420_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n376_), .A2(new_n378_), .B1(new_n264_), .B2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n411_), .A2(new_n419_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n403_), .B(new_n406_), .C1(new_n425_), .C2(new_n355_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n395_), .B1(new_n426_), .B2(new_n393_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT36), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT68), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT8), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT64), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(KEYINPUT6), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(KEYINPUT64), .ZN(new_n436_));
  INV_X1    g235(.A(G99gat), .ZN(new_n437_));
  INV_X1    g236(.A(G106gat), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n434_), .A2(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(KEYINPUT64), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n433_), .A2(KEYINPUT6), .ZN(new_n441_));
  AND2_X1   g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT66), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n444_), .A2(new_n437_), .A3(new_n438_), .A4(KEYINPUT7), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n437_), .A2(new_n438_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(KEYINPUT7), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT7), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT66), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n439_), .A2(new_n443_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(G85gat), .ZN(new_n452_));
  INV_X1    g251(.A(G92gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G85gat), .A2(G92gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n432_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n457_));
  OAI22_X1  g256(.A1(new_n448_), .A2(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n444_), .A2(KEYINPUT7), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n445_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n442_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n460_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n456_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n430_), .A2(KEYINPUT67), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n432_), .B2(KEYINPUT67), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n463_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n438_), .A3(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n454_), .A2(KEYINPUT9), .A3(new_n455_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n455_), .A2(KEYINPUT9), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n439_), .A2(new_n443_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT65), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n461_), .A2(new_n462_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT65), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n457_), .B(new_n467_), .C1(new_n475_), .C2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G29gat), .B(G36gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT35), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT77), .B(KEYINPUT34), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G232gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n481_), .A2(new_n484_), .B1(new_n485_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT78), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n484_), .B(KEYINPUT15), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n480_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n480_), .A2(new_n491_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT78), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n489_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n488_), .A2(new_n485_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n489_), .A2(new_n494_), .A3(new_n498_), .A4(new_n492_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G190gat), .B(G218gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT79), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G134gat), .B(G162gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n497_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n497_), .A2(KEYINPUT80), .A3(new_n499_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n428_), .A2(new_n505_), .B1(new_n506_), .B2(new_n503_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n428_), .A3(new_n503_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n427_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT13), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT11), .ZN(new_n514_));
  INV_X1    g313(.A(G71gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT69), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT69), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G71gat), .ZN(new_n518_));
  INV_X1    g317(.A(G78gat), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n514_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n516_), .A2(new_n518_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(G78gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(KEYINPUT11), .A3(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G57gat), .B(G64gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n522_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n524_), .A2(KEYINPUT11), .A3(new_n529_), .A4(new_n525_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n479_), .A2(new_n475_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n456_), .B1(new_n474_), .B2(new_n460_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n467_), .B1(new_n533_), .B2(new_n431_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n531_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT71), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n528_), .A2(new_n530_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n478_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n473_), .A2(KEYINPUT65), .A3(new_n474_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n538_), .A2(new_n541_), .A3(new_n467_), .A4(new_n457_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT70), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n431_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n533_), .B2(new_n466_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n546_), .A2(KEYINPUT70), .A3(new_n538_), .A4(new_n541_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n480_), .A2(KEYINPUT71), .A3(new_n531_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n537_), .A2(new_n544_), .A3(new_n547_), .A4(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT12), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT72), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n480_), .A2(new_n531_), .A3(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n480_), .B2(new_n531_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n542_), .A2(new_n550_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G120gat), .B(G148gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n552_), .A2(new_n561_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT75), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n549_), .A2(new_n551_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(KEYINPUT75), .A3(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT76), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n544_), .A2(new_n547_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n480_), .A2(KEYINPUT71), .A3(new_n531_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT71), .B1(new_n480_), .B2(new_n531_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n550_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n480_), .A2(new_n531_), .A3(new_n554_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n538_), .B1(new_n546_), .B2(new_n541_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(new_n556_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(new_n559_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT73), .B1(new_n579_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT73), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n552_), .A2(new_n585_), .A3(new_n561_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n566_), .A3(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n573_), .A2(new_n574_), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n574_), .B1(new_n573_), .B2(new_n587_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n513_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n568_), .A2(new_n569_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT75), .B1(new_n571_), .B2(new_n567_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n566_), .B1(new_n571_), .B2(new_n585_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n579_), .A2(KEYINPUT73), .A3(new_n583_), .ZN(new_n594_));
  OAI22_X1  g393(.A1(new_n591_), .A2(new_n592_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT76), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n573_), .A2(new_n587_), .A3(new_n574_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(KEYINPUT13), .A3(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n590_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G15gat), .B(G22gat), .ZN(new_n601_));
  INV_X1    g400(.A(G1gat), .ZN(new_n602_));
  INV_X1    g401(.A(G8gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT14), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G1gat), .B(G8gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(new_n484_), .Z(new_n608_));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n491_), .A2(new_n607_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n607_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n484_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n614_), .A3(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G169gat), .B(G197gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT86), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n611_), .A2(new_n615_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT87), .B1(new_n622_), .B2(new_n619_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT87), .ZN(new_n624_));
  INV_X1    g423(.A(new_n619_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n616_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n621_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT88), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(KEYINPUT88), .B(new_n621_), .C1(new_n623_), .C2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n607_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(new_n531_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G127gat), .B(G155gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G183gat), .B(G211gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(KEYINPUT17), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(KEYINPUT17), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n635_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT85), .Z(new_n644_));
  NAND2_X1  g443(.A1(new_n635_), .A2(new_n641_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT84), .Z(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n600_), .A2(new_n632_), .A3(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n512_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(new_n380_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(new_n602_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n427_), .A2(new_n632_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(KEYINPUT81), .A2(KEYINPUT37), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n654_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(KEYINPUT81), .A2(KEYINPUT37), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT82), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n654_), .B(new_n657_), .C1(new_n507_), .C2(new_n509_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n647_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n653_), .A2(new_n599_), .A3(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n602_), .A3(new_n380_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n651_), .B1(new_n652_), .B2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n664_), .B1(new_n652_), .B2(new_n663_), .ZN(G1324gat));
  NAND3_X1  g464(.A1(new_n662_), .A2(new_n603_), .A3(new_n289_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n649_), .A2(new_n289_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(G8gat), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT39), .B(new_n603_), .C1(new_n649_), .C2(new_n289_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(G1325gat));
  NAND3_X1  g472(.A1(new_n662_), .A2(new_n386_), .A3(new_n392_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n649_), .A2(new_n392_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n675_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT41), .B1(new_n675_), .B2(G15gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n674_), .B1(new_n676_), .B2(new_n677_), .ZN(G1326gat));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n662_), .A2(new_n679_), .A3(new_n355_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n649_), .A2(new_n355_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(G22gat), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT42), .B(new_n679_), .C1(new_n649_), .C2(new_n355_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT109), .ZN(G1327gat));
  INV_X1    g485(.A(new_n647_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(new_n510_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n599_), .A2(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n653_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n380_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT112), .B1(KEYINPUT111), .B2(KEYINPUT44), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n403_), .A2(new_n406_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n411_), .A2(new_n419_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n422_), .A2(new_n424_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n355_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n393_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n395_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n659_), .A2(new_n660_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n700_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n427_), .B2(new_n702_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n599_), .A2(new_n631_), .A3(new_n647_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n693_), .B1(new_n706_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n704_), .A2(new_n705_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n708_), .B(KEYINPUT110), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n692_), .A4(new_n707_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n380_), .A2(G29gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n691_), .B1(new_n716_), .B2(new_n717_), .ZN(G1328gat));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n653_), .A2(new_n719_), .A3(new_n289_), .A4(new_n689_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT45), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n402_), .B1(new_n712_), .B2(new_n715_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n719_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT46), .B(new_n721_), .C1(new_n722_), .C2(new_n719_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1329gat));
  INV_X1    g526(.A(G43gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n690_), .A2(new_n728_), .A3(new_n392_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n393_), .B1(new_n712_), .B2(new_n715_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(new_n728_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OAI211_X1 g532(.A(KEYINPUT47), .B(new_n729_), .C1(new_n730_), .C2(new_n728_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1330gat));
  AOI21_X1  g534(.A(G50gat), .B1(new_n690_), .B2(new_n355_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n355_), .A2(G50gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n716_), .B2(new_n737_), .ZN(G1331gat));
  NOR2_X1   g537(.A1(new_n427_), .A2(new_n631_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n739_), .A2(new_n600_), .A3(new_n661_), .ZN(new_n740_));
  INV_X1    g539(.A(G57gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n380_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n599_), .A2(new_n631_), .A3(new_n647_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n512_), .A2(new_n380_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G57gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n742_), .A2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(G64gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n740_), .A2(new_n747_), .A3(new_n289_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n512_), .A2(new_n289_), .A3(new_n743_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G64gat), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT48), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT48), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1333gat));
  NAND3_X1  g552(.A1(new_n740_), .A2(new_n515_), .A3(new_n392_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n512_), .A2(new_n392_), .A3(new_n743_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(G71gat), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G71gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1334gat));
  NAND3_X1  g558(.A1(new_n740_), .A2(new_n519_), .A3(new_n355_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n512_), .A2(new_n355_), .A3(new_n743_), .ZN(new_n761_));
  XOR2_X1   g560(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(G78gat), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(G78gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(G1335gat));
  NOR3_X1   g564(.A1(new_n599_), .A2(new_n631_), .A3(new_n687_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n713_), .A2(new_n766_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n767_), .A2(new_n452_), .A3(new_n379_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n739_), .A2(new_n600_), .A3(new_n688_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT115), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n452_), .B1(new_n770_), .B2(new_n379_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT116), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n452_), .C1(new_n770_), .C2(new_n379_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n768_), .B1(new_n772_), .B2(new_n774_), .ZN(G1336gat));
  OAI21_X1  g574(.A(G92gat), .B1(new_n767_), .B2(new_n402_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n289_), .A2(new_n453_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n770_), .B2(new_n777_), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n767_), .B2(new_n393_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n392_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n770_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n713_), .A2(new_n355_), .A3(new_n766_), .ZN(new_n783_));
  XOR2_X1   g582(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n784_));
  AND3_X1   g583(.A1(new_n783_), .A2(G106gat), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n783_), .B2(G106gat), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n355_), .A2(new_n438_), .ZN(new_n787_));
  OAI22_X1  g586(.A1(new_n785_), .A2(new_n786_), .B1(new_n770_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  OAI221_X1 g590(.A(new_n789_), .B1(new_n770_), .B2(new_n787_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1339gat));
  OR2_X1    g592(.A1(new_n623_), .A2(new_n626_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n608_), .A2(new_n609_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n612_), .A2(new_n614_), .A3(new_n610_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n625_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n794_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n575_), .A2(new_n558_), .A3(KEYINPUT119), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n544_), .A2(new_n547_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n582_), .B2(new_n802_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n800_), .A2(new_n803_), .A3(new_n551_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n582_), .B2(new_n559_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n557_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n560_), .A2(new_n807_), .A3(KEYINPUT55), .A4(new_n580_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n566_), .B1(new_n804_), .B2(new_n809_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n810_), .A2(KEYINPUT56), .B1(new_n570_), .B2(new_n572_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n812_), .B(new_n566_), .C1(new_n804_), .C2(new_n809_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n631_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n511_), .B1(new_n799_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT57), .B1(new_n815_), .B2(KEYINPUT120), .ZN(new_n816_));
  INV_X1    g615(.A(new_n798_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n807_), .A2(new_n544_), .A3(new_n547_), .A4(new_n580_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n550_), .B1(new_n819_), .B2(new_n801_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n809_), .B1(new_n800_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n567_), .ZN(new_n822_));
  AND4_X1   g621(.A1(new_n631_), .A2(new_n822_), .A3(new_n573_), .A4(new_n813_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n510_), .B1(new_n818_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n811_), .A2(KEYINPUT58), .A3(new_n798_), .A4(new_n813_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n822_), .A2(new_n798_), .A3(new_n573_), .A4(new_n813_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n703_), .A2(new_n828_), .A3(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n816_), .A2(new_n827_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n647_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n661_), .A2(new_n632_), .A3(new_n598_), .A4(new_n590_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT54), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n599_), .A2(new_n837_), .A3(new_n632_), .A4(new_n661_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n356_), .A2(new_n380_), .A3(new_n392_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT59), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n833_), .A2(new_n647_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n841_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(G113gat), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n632_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n840_), .A2(new_n842_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n850_), .B2(new_n632_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n851_), .A2(new_n852_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n849_), .B1(new_n853_), .B2(new_n854_), .ZN(G1340gat));
  OAI21_X1  g654(.A(G120gat), .B1(new_n847_), .B2(new_n599_), .ZN(new_n856_));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n599_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(KEYINPUT60), .B2(new_n857_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n850_), .B2(new_n859_), .ZN(G1341gat));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n847_), .A2(new_n861_), .A3(new_n647_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n850_), .B2(new_n647_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n863_), .A2(new_n864_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n862_), .B1(new_n865_), .B2(new_n866_), .ZN(G1342gat));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n702_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n870_));
  AND4_X1   g669(.A1(new_n660_), .A2(new_n831_), .A3(new_n828_), .A4(new_n659_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n824_), .A2(new_n825_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(KEYINPUT57), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n687_), .B1(new_n873_), .B2(new_n827_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n836_), .A2(new_n838_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n511_), .B(new_n842_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n868_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n876_), .B2(new_n868_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n870_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT124), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n870_), .B(new_n882_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1343gat));
  NAND2_X1  g683(.A1(new_n355_), .A2(new_n393_), .ZN(new_n885_));
  NOR4_X1   g684(.A1(new_n844_), .A2(new_n289_), .A3(new_n379_), .A4(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n631_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n600_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n687_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1346gat));
  NAND3_X1  g692(.A1(new_n886_), .A2(new_n292_), .A3(new_n511_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n886_), .A2(new_n703_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n292_), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n402_), .A2(new_n380_), .ZN(new_n897_));
  AOI21_X1  g696(.A(KEYINPUT125), .B1(new_n897_), .B2(new_n392_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n355_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n392_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n844_), .A2(new_n898_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n631_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G169gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n906_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n904_), .A2(G169gat), .A3(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n907_), .B(new_n909_), .C1(new_n234_), .C2(new_n904_), .ZN(G1348gat));
  NAND2_X1  g709(.A1(new_n903_), .A2(new_n600_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g711(.A1(new_n903_), .A2(new_n687_), .ZN(new_n913_));
  MUX2_X1   g712(.A(new_n230_), .B(G183gat), .S(new_n913_), .Z(G1350gat));
  INV_X1    g713(.A(new_n248_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n903_), .A2(new_n915_), .A3(new_n511_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n903_), .A2(new_n703_), .ZN(new_n917_));
  INV_X1    g716(.A(G190gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(G1351gat));
  NOR4_X1   g718(.A1(new_n844_), .A2(new_n402_), .A3(new_n380_), .A4(new_n885_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n631_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n600_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n925_));
  INV_X1    g724(.A(G211gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n687_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT127), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n920_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n926_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1354gat));
  INV_X1    g730(.A(G218gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n920_), .A2(new_n932_), .A3(new_n511_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n920_), .A2(new_n703_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n934_), .B2(new_n932_), .ZN(G1355gat));
endmodule


