//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n604_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G85gat), .B(G92gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR3_X1   g004(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n203_), .B1(new_n207_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n202_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n203_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n209_), .A2(new_n211_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n204_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n216_), .B1(new_n217_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT64), .B1(new_n217_), .B2(new_n222_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n207_), .A2(new_n226_), .A3(new_n212_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n203_), .A2(KEYINPUT8), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n215_), .A2(new_n224_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT10), .B(G99gat), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n220_), .ZN(new_n233_));
  INV_X1    g032(.A(G85gat), .ZN(new_n234_));
  INV_X1    g033(.A(G92gat), .ZN(new_n235_));
  OR3_X1    g034(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT9), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n231_), .A2(new_n233_), .A3(new_n236_), .A4(new_n212_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n230_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G57gat), .B(G64gat), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n241_));
  XOR2_X1   g040(.A(G71gat), .B(G78gat), .Z(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n241_), .A2(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n238_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT66), .B(KEYINPUT12), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(KEYINPUT67), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n245_), .B1(new_n230_), .B2(new_n237_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n252_), .B2(new_n248_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(KEYINPUT12), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n230_), .A2(new_n245_), .A3(new_n237_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G230gat), .A2(G233gat), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n250_), .A2(new_n253_), .A3(new_n254_), .A4(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n247_), .A2(new_n255_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT69), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G176gat), .B(G204gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n262_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n258_), .A2(new_n261_), .A3(new_n268_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n262_), .A2(KEYINPUT70), .A3(new_n269_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n274_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT13), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(KEYINPUT71), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT72), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n277_), .A2(new_n283_), .A3(new_n280_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G15gat), .B(G22gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G1gat), .A2(G8gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT14), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G1gat), .ZN(new_n290_));
  INV_X1    g089(.A(G8gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n287_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n286_), .A2(new_n287_), .A3(new_n292_), .A4(new_n288_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G43gat), .B(G50gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G36gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G29gat), .ZN(new_n300_));
  INV_X1    g099(.A(G29gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G36gat), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n300_), .A2(new_n302_), .A3(KEYINPUT75), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT75), .B1(new_n300_), .B2(new_n302_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n298_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n301_), .A2(G36gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n299_), .A2(G29gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n300_), .A2(new_n302_), .A3(KEYINPUT75), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n297_), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n305_), .A2(KEYINPUT15), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT15), .B1(new_n305_), .B2(new_n311_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n296_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n305_), .A2(new_n311_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT82), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n305_), .A2(new_n311_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n296_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n315_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n316_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT81), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT81), .ZN(new_n324_));
  AOI211_X1 g123(.A(new_n324_), .B(new_n316_), .C1(new_n320_), .C2(new_n315_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n318_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G113gat), .B(G141gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT83), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G169gat), .B(G197gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n326_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT84), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n318_), .B(new_n330_), .C1(new_n323_), .C2(new_n325_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(KEYINPUT84), .A3(new_n331_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n285_), .A2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n238_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n230_), .A2(new_n311_), .A3(new_n305_), .A4(new_n237_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G232gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n343_), .A2(KEYINPUT35), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n339_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(KEYINPUT35), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT74), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n339_), .A2(new_n340_), .A3(new_n344_), .A4(new_n347_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT36), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G190gat), .B(G218gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G134gat), .B(G162gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n352_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n349_), .A2(new_n356_), .A3(new_n351_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n353_), .B1(new_n352_), .B2(new_n357_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n362_), .B(KEYINPUT100), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT23), .ZN(new_n366_));
  OR2_X1    g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(KEYINPUT24), .A3(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  NOR3_X1   g169(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT25), .B(G183gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT26), .B(G190gat), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G204gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(G197gat), .ZN(new_n377_));
  INV_X1    g176(.A(G197gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(G204gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT21), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G211gat), .B(G218gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n376_), .B2(G197gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n378_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n383_), .B(new_n384_), .C1(new_n378_), .C2(G204gat), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n380_), .B(new_n381_), .C1(new_n385_), .C2(KEYINPUT21), .ZN(new_n386_));
  INV_X1    g185(.A(new_n381_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(KEYINPUT21), .A3(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n366_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G169gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n375_), .A2(new_n386_), .A3(new_n388_), .A4(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT22), .B(G169gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT94), .ZN(new_n396_));
  INV_X1    g195(.A(G176gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n390_), .A2(new_n368_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n398_), .A2(new_n399_), .B1(new_n374_), .B2(new_n370_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n386_), .A2(new_n388_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT20), .B(new_n394_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT19), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n400_), .A2(new_n401_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT20), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n375_), .A2(new_n393_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n386_), .A2(new_n388_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n404_), .B1(new_n407_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n406_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT95), .ZN(new_n415_));
  XOR2_X1   g214(.A(G8gat), .B(G36gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT18), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(new_n415_), .A3(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n402_), .A2(new_n405_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n421_), .B2(new_n412_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT95), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G127gat), .B(G134gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G113gat), .B(G120gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n426_), .B(KEYINPUT86), .Z(new_n427_));
  NAND2_X1  g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT89), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT89), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(G155gat), .A3(G162gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  OR3_X1    g231(.A1(new_n432_), .A2(KEYINPUT90), .A3(KEYINPUT1), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT90), .B1(new_n432_), .B2(KEYINPUT1), .ZN(new_n434_));
  INV_X1    g233(.A(G155gat), .ZN(new_n435_));
  INV_X1    g234(.A(G162gat), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n432_), .A2(KEYINPUT1), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n433_), .A2(new_n434_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G141gat), .A2(G148gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT88), .ZN(new_n440_));
  INV_X1    g239(.A(G141gat), .ZN(new_n441_));
  INV_X1    g240(.A(G148gat), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n439_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n442_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n445_), .A2(KEYINPUT2), .B1(new_n446_), .B2(KEYINPUT3), .ZN(new_n447_));
  OAI221_X1 g246(.A(new_n447_), .B1(KEYINPUT3), .B2(new_n446_), .C1(new_n440_), .C2(KEYINPUT2), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n429_), .A2(new_n431_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n444_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n427_), .A2(new_n451_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n438_), .A2(new_n443_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n426_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(KEYINPUT4), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G225gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n427_), .A2(new_n451_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G1gat), .B(G29gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G57gat), .B(G85gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n462_), .B(new_n463_), .Z(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n456_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n452_), .A2(new_n454_), .A3(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n459_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n421_), .A2(new_n412_), .A3(new_n419_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AND4_X1   g269(.A1(new_n420_), .A2(new_n423_), .A3(new_n468_), .A4(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n455_), .A2(new_n466_), .A3(new_n458_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n452_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n464_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT98), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n472_), .A2(KEYINPUT33), .A3(new_n473_), .A4(new_n464_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n471_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n476_), .A2(KEYINPUT98), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n472_), .A2(new_n473_), .A3(new_n464_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n464_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n419_), .A2(KEYINPUT32), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n406_), .B2(new_n413_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n402_), .A2(new_n404_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n410_), .B(KEYINPUT92), .ZN(new_n490_));
  INV_X1    g289(.A(new_n400_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT20), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT99), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n409_), .A2(new_n410_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT99), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n495_), .B(KEYINPUT20), .C1(new_n490_), .C2(new_n491_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n493_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n489_), .B1(new_n497_), .B2(new_n404_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(new_n484_), .ZN(new_n499_));
  OAI22_X1  g298(.A1(new_n479_), .A2(new_n480_), .B1(new_n488_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G71gat), .B(G99gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(G43gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n409_), .B(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G227gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(G15gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT30), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n427_), .B(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n509_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G78gat), .B(G106gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(G228gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n401_), .B(KEYINPUT92), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT29), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n453_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n516_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n451_), .A2(KEYINPUT29), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n401_), .A2(new_n516_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n515_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n490_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n526_), .A2(new_n516_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n515_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT93), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n453_), .A2(new_n518_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G22gat), .B(G50gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT28), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n530_), .B(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n525_), .A2(new_n528_), .A3(new_n529_), .A4(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n525_), .A2(new_n528_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n513_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n534_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT93), .B1(new_n527_), .B2(new_n515_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n540_), .A2(new_n533_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n513_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n534_), .A3(new_n512_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT27), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n423_), .A2(new_n470_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n420_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  OAI211_X1 g347(.A(KEYINPUT27), .B(new_n422_), .C1(new_n498_), .C2(new_n419_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n481_), .A2(new_n482_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n500_), .A2(new_n538_), .B1(new_n544_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n296_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(new_n246_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT79), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G127gat), .B(G155gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G183gat), .B(G211gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT17), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n556_), .B(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n561_), .A2(KEYINPUT17), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n563_), .B1(new_n555_), .B2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT80), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n364_), .A2(new_n552_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n338_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(G1gat), .B1(new_n568_), .B2(new_n550_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT101), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n337_), .B(KEYINPUT85), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n361_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(new_n359_), .A3(new_n358_), .A4(new_n573_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(new_n566_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR4_X1   g379(.A1(new_n285_), .A2(new_n552_), .A3(new_n572_), .A4(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n290_), .A3(new_n483_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT38), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n570_), .A2(new_n583_), .ZN(G1324gat));
  AND2_X1   g383(.A1(new_n548_), .A2(new_n549_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G8gat), .B1(new_n568_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT102), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n586_), .A2(new_n587_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n590_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n585_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n581_), .A2(new_n291_), .A3(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n592_), .A2(KEYINPUT40), .A3(new_n593_), .A4(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT40), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n595_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n591_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(G1325gat));
  OAI21_X1  g399(.A(G15gat), .B1(new_n568_), .B2(new_n512_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT41), .Z(new_n602_));
  INV_X1    g401(.A(G15gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n581_), .A2(new_n603_), .A3(new_n513_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(G1326gat));
  NOR2_X1   g404(.A1(new_n539_), .A2(new_n541_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G22gat), .B1(new_n568_), .B2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT42), .ZN(new_n609_));
  INV_X1    g408(.A(G22gat), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n581_), .A2(new_n610_), .A3(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(G1327gat));
  INV_X1    g411(.A(new_n362_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n566_), .A2(new_n613_), .ZN(new_n614_));
  NOR4_X1   g413(.A1(new_n285_), .A2(new_n552_), .A3(new_n572_), .A4(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n301_), .A3(new_n483_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT43), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n575_), .A2(new_n577_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n552_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n566_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n544_), .A2(new_n551_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n469_), .B1(KEYINPUT95), .B2(new_n422_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n622_), .A2(new_n478_), .A3(new_n420_), .A4(new_n468_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n624_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n623_), .A2(new_n480_), .A3(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n499_), .A2(new_n550_), .A3(new_n486_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n538_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n618_), .B1(new_n621_), .B2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n620_), .B1(new_n629_), .B2(KEYINPUT43), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n338_), .A2(new_n619_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n632_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n483_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(KEYINPUT103), .ZN(new_n637_));
  OAI21_X1  g436(.A(G29gat), .B1(new_n636_), .B2(KEYINPUT103), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n616_), .B1(new_n637_), .B2(new_n638_), .ZN(G1328gat));
  NAND2_X1  g438(.A1(new_n633_), .A2(new_n634_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G36gat), .B1(new_n640_), .B2(new_n585_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n615_), .A2(new_n299_), .A3(new_n594_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT45), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(G1329gat));
  NAND3_X1  g445(.A1(new_n635_), .A2(G43gat), .A3(new_n513_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n615_), .A2(new_n513_), .ZN(new_n648_));
  INV_X1    g447(.A(G43gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n647_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT47), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT47), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n647_), .A2(new_n655_), .A3(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1330gat));
  AOI21_X1  g456(.A(G50gat), .B1(new_n615_), .B2(new_n606_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n606_), .A2(G50gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n635_), .B2(new_n659_), .ZN(G1331gat));
  AND3_X1   g459(.A1(new_n282_), .A2(new_n337_), .A3(new_n284_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n621_), .A2(new_n628_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n580_), .ZN(new_n664_));
  INV_X1    g463(.A(G57gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n665_), .A3(new_n483_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n662_), .A2(new_n620_), .A3(new_n363_), .A4(new_n572_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n282_), .A2(new_n284_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n667_), .A2(new_n550_), .A3(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n666_), .B1(new_n669_), .B2(new_n665_), .ZN(G1332gat));
  INV_X1    g469(.A(G64gat), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n667_), .A2(new_n668_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n594_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT48), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n664_), .A2(new_n671_), .A3(new_n594_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1333gat));
  INV_X1    g475(.A(G71gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n664_), .A2(new_n677_), .A3(new_n513_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n672_), .A2(new_n513_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G71gat), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(KEYINPUT49), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(KEYINPUT49), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT106), .ZN(G1334gat));
  INV_X1    g483(.A(G78gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n664_), .A2(new_n685_), .A3(new_n606_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n672_), .A2(new_n606_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G78gat), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT50), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT50), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT107), .Z(G1335gat));
  NAND3_X1  g491(.A1(new_n662_), .A2(KEYINPUT43), .A3(new_n578_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n619_), .A2(new_n693_), .A3(new_n566_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n282_), .A2(new_n337_), .A3(new_n284_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT108), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n630_), .A2(new_n661_), .A3(new_n697_), .A4(new_n619_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G85gat), .B1(new_n700_), .B2(new_n550_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n663_), .A2(new_n614_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n234_), .A3(new_n483_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1336gat));
  OAI21_X1  g503(.A(G92gat), .B1(new_n700_), .B2(new_n585_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n702_), .A2(new_n235_), .A3(new_n594_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1337gat));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n702_), .A2(new_n232_), .A3(new_n513_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n699_), .A2(new_n513_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(G99gat), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT51), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n702_), .A2(new_n232_), .A3(new_n513_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n512_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n714_), .B(new_n715_), .C1(new_n716_), .C2(new_n219_), .ZN(new_n717_));
  AOI22_X1  g516(.A1(new_n711_), .A2(new_n713_), .B1(new_n717_), .B2(new_n712_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n708_), .B1(new_n718_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n717_), .A2(new_n712_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n715_), .B(new_n713_), .C1(new_n716_), .C2(new_n219_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(KEYINPUT111), .A3(new_n720_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n722_), .A2(new_n726_), .ZN(G1338gat));
  NOR2_X1   g526(.A1(new_n694_), .A2(new_n695_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n220_), .B1(new_n728_), .B2(new_n606_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT52), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n702_), .A2(new_n220_), .A3(new_n606_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT53), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n730_), .A2(new_n734_), .A3(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1339gat));
  INV_X1    g535(.A(KEYINPUT54), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n571_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n579_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n579_), .B2(new_n738_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n742_));
  INV_X1    g541(.A(new_n334_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n317_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n314_), .A2(new_n315_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n330_), .B1(new_n321_), .B2(new_n317_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n743_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n273_), .A2(new_n274_), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n250_), .A2(new_n253_), .A3(new_n255_), .A4(new_n254_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n260_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n258_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n248_), .B1(new_n238_), .B2(new_n246_), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n754_), .A2(KEYINPUT67), .B1(KEYINPUT12), .B2(new_n252_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n755_), .A2(KEYINPUT55), .A3(new_n253_), .A4(new_n257_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n751_), .A2(new_n753_), .A3(new_n756_), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n749_), .B(KEYINPUT56), .C1(new_n757_), .C2(new_n269_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759_));
  INV_X1    g558(.A(new_n272_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n337_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n272_), .A2(KEYINPUT112), .A3(new_n336_), .A4(new_n335_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n758_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n757_), .A2(new_n269_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n269_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n749_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n748_), .B1(new_n764_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n742_), .B1(new_n770_), .B2(new_n613_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n748_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n269_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT56), .B1(new_n757_), .B2(new_n269_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(KEYINPUT113), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n765_), .A2(KEYINPUT113), .A3(new_n766_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n762_), .A3(new_n761_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n772_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n362_), .A2(KEYINPUT57), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n747_), .A2(new_n272_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n747_), .A2(new_n272_), .A3(KEYINPUT115), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n786_), .B(KEYINPUT58), .C1(new_n773_), .C2(new_n774_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n578_), .A3(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n771_), .A2(new_n781_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n620_), .B1(new_n792_), .B2(KEYINPUT116), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n771_), .A2(new_n794_), .A3(new_n781_), .A4(new_n791_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n741_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n585_), .A2(new_n483_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n796_), .A2(new_n542_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n337_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G113gat), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n797_), .A2(KEYINPUT59), .A3(new_n542_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n792_), .A2(new_n566_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT117), .ZN(new_n803_));
  INV_X1    g602(.A(new_n741_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n802_), .A2(KEYINPUT117), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n801_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n798_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n571_), .A2(G113gat), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT118), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n800_), .B1(new_n810_), .B2(new_n812_), .ZN(G1340gat));
  OAI21_X1  g612(.A(G120gat), .B1(new_n809_), .B2(new_n668_), .ZN(new_n814_));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n668_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n798_), .B(new_n816_), .C1(KEYINPUT60), .C2(new_n815_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(G1341gat));
  OAI21_X1  g617(.A(G127gat), .B1(new_n809_), .B2(new_n566_), .ZN(new_n819_));
  INV_X1    g618(.A(G127gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n798_), .A2(new_n820_), .A3(new_n620_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1342gat));
  AOI21_X1  g621(.A(G134gat), .B1(new_n798_), .B2(new_n364_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n578_), .A2(G134gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT119), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n810_), .B2(new_n825_), .ZN(G1343gat));
  OAI21_X1  g625(.A(new_n791_), .B1(new_n770_), .B2(new_n779_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n742_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n778_), .B2(new_n362_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT116), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(new_n566_), .A3(new_n795_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n804_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n797_), .A2(new_n543_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n337_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(new_n441_), .ZN(G1344gat));
  NOR2_X1   g635(.A1(new_n834_), .A2(new_n668_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT120), .B(G148gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1345gat));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n840_));
  INV_X1    g639(.A(new_n834_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n620_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n834_), .A2(KEYINPUT121), .A3(new_n566_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT61), .B(G155gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n846_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1346gat));
  NAND3_X1  g649(.A1(new_n841_), .A2(new_n436_), .A3(new_n364_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n834_), .A2(new_n618_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n436_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT122), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n851_), .B(new_n855_), .C1(new_n436_), .C2(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1347gat));
  NOR2_X1   g656(.A1(new_n585_), .A2(new_n483_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n513_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n606_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n799_), .B(new_n860_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n861_), .A2(new_n862_), .A3(G169gat), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n805_), .A2(new_n806_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n860_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n799_), .A3(new_n396_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n862_), .B1(new_n861_), .B2(G169gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n863_), .B1(new_n867_), .B2(new_n868_), .ZN(G1348gat));
  NAND2_X1  g668(.A1(new_n866_), .A2(new_n285_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n796_), .A2(new_n606_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n668_), .A2(new_n397_), .A3(new_n859_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n870_), .A2(new_n397_), .B1(new_n871_), .B2(new_n872_), .ZN(G1349gat));
  NOR3_X1   g672(.A1(new_n865_), .A2(new_n566_), .A3(new_n372_), .ZN(new_n874_));
  INV_X1    g673(.A(G183gat), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n871_), .A2(new_n620_), .A3(new_n513_), .A4(new_n858_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(G1350gat));
  OAI21_X1  g676(.A(G190gat), .B1(new_n865_), .B2(new_n618_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n364_), .A2(new_n373_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT123), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n865_), .B2(new_n880_), .ZN(G1351gat));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n585_), .A2(new_n483_), .A3(new_n543_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n796_), .B2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n832_), .A2(KEYINPUT124), .A3(new_n883_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n799_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n668_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n376_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT124), .B1(new_n832_), .B2(new_n883_), .ZN(new_n893_));
  AOI211_X1 g692(.A(new_n882_), .B(new_n884_), .C1(new_n831_), .C2(new_n804_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n285_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(KEYINPUT125), .A3(G204gat), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n892_), .A2(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n376_), .B(new_n285_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n887_), .A2(KEYINPUT126), .A3(new_n376_), .A4(new_n285_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n897_), .A2(new_n902_), .ZN(G1353gat));
  AOI21_X1  g702(.A(new_n566_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n887_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT127), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n905_), .B(new_n908_), .ZN(G1354gat));
  INV_X1    g708(.A(new_n887_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G218gat), .B1(new_n910_), .B2(new_n618_), .ZN(new_n911_));
  INV_X1    g710(.A(G218gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n887_), .A2(new_n912_), .A3(new_n364_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1355gat));
endmodule


