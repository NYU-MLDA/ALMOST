//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n956_, new_n957_, new_n958_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_, new_n980_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT105), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT98), .ZN(new_n208_));
  INV_X1    g007(.A(G211gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G218gat), .ZN(new_n210_));
  INV_X1    g009(.A(G218gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(G211gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n208_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(G211gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(G218gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT98), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217_));
  INV_X1    g016(.A(G197gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G204gat), .ZN(new_n219_));
  INV_X1    g018(.A(G204gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G197gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n217_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n213_), .A2(new_n216_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT99), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n213_), .A2(KEYINPUT99), .A3(new_n222_), .A4(new_n216_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n219_), .A2(new_n221_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n229_));
  AOI22_X1  g028(.A1(new_n213_), .A2(new_n216_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n218_), .A2(KEYINPUT96), .A3(G204gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n219_), .A2(new_n221_), .ZN(new_n232_));
  OAI211_X1 g031(.A(KEYINPUT21), .B(new_n231_), .C1(new_n232_), .C2(KEYINPUT96), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n227_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G169gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT22), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT22), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G169gat), .ZN(new_n239_));
  INV_X1    g038(.A(G176gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT23), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(G183gat), .A3(G190gat), .ZN(new_n247_));
  INV_X1    g046(.A(G183gat), .ZN(new_n248_));
  INV_X1    g047(.A(G190gat), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n245_), .A2(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT104), .B1(new_n243_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n247_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(G183gat), .B2(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n242_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT22), .B(G169gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(new_n240_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT104), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n244_), .A2(new_n246_), .ZN(new_n259_));
  NOR3_X1   g058(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT25), .B(G183gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G190gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT24), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n265_), .B1(G169gat), .B2(G176gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n236_), .A2(new_n240_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n263_), .A2(new_n264_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n262_), .B1(new_n268_), .B2(KEYINPUT103), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(new_n264_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(KEYINPUT24), .A3(new_n242_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n270_), .A2(KEYINPUT103), .A3(new_n271_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n251_), .B(new_n258_), .C1(new_n269_), .C2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n207_), .B1(new_n235_), .B2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n244_), .B(new_n246_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n249_), .A2(KEYINPUT80), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT80), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G190gat), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n276_), .A2(new_n278_), .A3(new_n248_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n242_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n238_), .A2(KEYINPUT84), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT84), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT22), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(G169gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n237_), .A2(new_n240_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(G169gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(KEYINPUT85), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n280_), .B1(new_n286_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n271_), .A2(KEYINPUT83), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT83), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n266_), .A2(new_n292_), .A3(new_n267_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n262_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT81), .B1(new_n249_), .B2(KEYINPUT26), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT81), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT26), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(G190gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n276_), .A2(new_n278_), .A3(KEYINPUT26), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n263_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT82), .A4(new_n263_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n294_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n235_), .B1(new_n290_), .B2(new_n305_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n225_), .A2(new_n226_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n268_), .A2(KEYINPUT103), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n268_), .A2(KEYINPUT103), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n262_), .A3(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n258_), .A2(new_n251_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n307_), .A2(new_n310_), .A3(KEYINPUT105), .A4(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n274_), .A2(new_n306_), .A3(new_n312_), .A4(KEYINPUT20), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT19), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n303_), .A2(new_n304_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n294_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n289_), .A2(new_n286_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n280_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n307_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n235_), .A2(new_n273_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(KEYINPUT20), .A4(new_n315_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n206_), .B1(new_n317_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n326_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n316_), .B2(new_n313_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n206_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT27), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G1gat), .B(G29gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G85gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT0), .B(G57gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n334_), .B(new_n335_), .Z(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT89), .ZN(new_n338_));
  INV_X1    g137(.A(G127gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(G134gat), .ZN(new_n340_));
  INV_X1    g139(.A(G134gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(G127gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n338_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(G127gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(G134gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(KEYINPUT89), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G113gat), .B(G120gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n346_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G113gat), .B(G120gat), .Z(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G141gat), .A2(G148gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n357_), .A2(KEYINPUT94), .A3(KEYINPUT1), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT94), .B1(new_n357_), .B2(KEYINPUT1), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT93), .ZN(new_n361_));
  INV_X1    g160(.A(G155gat), .ZN(new_n362_));
  INV_X1    g161(.A(G162gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT93), .B1(G155gat), .B2(G162gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT1), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(G155gat), .A3(G162gat), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n356_), .B1(new_n360_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(new_n365_), .A3(new_n357_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT2), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n352_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n370_), .B1(new_n374_), .B2(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n348_), .B(new_n351_), .C1(new_n369_), .C2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n357_), .A2(KEYINPUT1), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT94), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n357_), .A2(KEYINPUT94), .A3(KEYINPUT1), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n355_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n354_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n389_), .A2(new_n376_), .A3(new_n377_), .A4(new_n371_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n390_), .A2(new_n364_), .A3(new_n365_), .A4(new_n357_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n343_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n347_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n387_), .B(new_n391_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n380_), .A2(new_n394_), .A3(KEYINPUT4), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT106), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n380_), .A2(new_n394_), .A3(KEYINPUT106), .A4(KEYINPUT4), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT107), .ZN(new_n400_));
  OAI211_X1 g199(.A(G225gat), .B(G233gat), .C1(new_n380_), .C2(KEYINPUT4), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n380_), .A2(new_n394_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n401_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(new_n400_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n337_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n408_), .A2(new_n400_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n408_), .A2(new_n400_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n336_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n306_), .A2(KEYINPUT20), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n253_), .A2(new_n256_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n307_), .A2(new_n310_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n315_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n324_), .A2(new_n325_), .A3(KEYINPUT20), .A4(new_n316_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n205_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n327_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n332_), .A2(new_n414_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT87), .Z(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G99gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n320_), .A2(new_n323_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT30), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n320_), .A2(new_n323_), .A3(KEYINPUT30), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G15gat), .B(G43gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT86), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G71gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n431_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n436_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n428_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n431_), .A2(new_n432_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n435_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(new_n427_), .A3(new_n437_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n351_), .A2(new_n348_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT31), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT90), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(KEYINPUT90), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n440_), .A2(new_n443_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n447_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT91), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n440_), .A2(new_n443_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n448_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT91), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n440_), .A2(new_n443_), .A3(new_n450_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n453_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT29), .B1(new_n369_), .B2(new_n379_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT95), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n387_), .A2(new_n391_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(KEYINPUT95), .A3(KEYINPUT29), .ZN(new_n464_));
  INV_X1    g263(.A(G228gat), .ZN(new_n465_));
  INV_X1    g264(.A(G233gat), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n462_), .A2(new_n235_), .A3(new_n464_), .A4(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT100), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n307_), .A2(new_n467_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT100), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n464_), .A4(new_n462_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n468_), .B1(new_n235_), .B2(new_n460_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G78gat), .B(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT101), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G22gat), .B(G50gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT28), .B1(new_n463_), .B2(KEYINPUT29), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n463_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n483_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n484_), .A3(new_n482_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n475_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n490_), .B1(new_n491_), .B2(new_n479_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n481_), .A2(new_n492_), .A3(KEYINPUT102), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT102), .ZN(new_n494_));
  INV_X1    g293(.A(new_n490_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n491_), .A2(new_n479_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n494_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n478_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n490_), .B1(new_n477_), .B2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n491_), .A2(new_n478_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n493_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n424_), .A2(new_n459_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT33), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n413_), .A2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n317_), .A2(new_n326_), .A3(new_n206_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(new_n327_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n411_), .A2(new_n412_), .A3(KEYINPUT33), .A4(new_n336_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n404_), .A2(KEYINPUT108), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n511_), .A2(new_n405_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n404_), .A2(KEYINPUT108), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n336_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n380_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n399_), .A2(new_n405_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT109), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT109), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n399_), .A2(new_n520_), .A3(new_n405_), .A4(new_n517_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n514_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .A4(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n317_), .A2(new_n326_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT32), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n524_), .B1(new_n525_), .B2(new_n206_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT20), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n429_), .B2(new_n235_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n316_), .B1(new_n528_), .B2(new_n417_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n420_), .ZN(new_n530_));
  OAI211_X1 g329(.A(KEYINPUT32), .B(new_n205_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n414_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n523_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n503_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n481_), .A2(new_n492_), .A3(KEYINPUT102), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n495_), .B1(new_n491_), .B2(new_n478_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(new_n491_), .B2(new_n478_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT102), .B1(new_n481_), .B2(new_n492_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n535_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT110), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n424_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n422_), .B1(new_n508_), .B2(new_n327_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n206_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n543_), .B(KEYINPUT27), .C1(new_n330_), .C2(new_n206_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n542_), .A2(new_n410_), .A3(new_n413_), .A4(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT110), .B1(new_n503_), .B2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n534_), .A2(new_n541_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT92), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n459_), .B(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n505_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G15gat), .B(G22gat), .ZN(new_n551_));
  INV_X1    g350(.A(G1gat), .ZN(new_n552_));
  INV_X1    g351(.A(G8gat), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT14), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G1gat), .B(G8gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G29gat), .B(G36gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G43gat), .B(G50gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(KEYINPUT15), .Z(new_n562_));
  OAI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(new_n557_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT78), .B1(new_n557_), .B2(new_n560_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n557_), .A2(new_n560_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n565_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G113gat), .B(G141gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G169gat), .B(G197gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT79), .B1(new_n571_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT79), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n566_), .A2(new_n577_), .A3(new_n570_), .A4(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n571_), .A2(new_n575_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  OR3_X1    g381(.A1(new_n550_), .A2(KEYINPUT111), .A3(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT111), .B1(new_n550_), .B2(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT34), .Z(new_n587_));
  INV_X1    g386(.A(KEYINPUT35), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n588_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT70), .Z(new_n592_));
  XOR2_X1   g391(.A(G85gat), .B(G92gat), .Z(new_n593_));
  NOR2_X1   g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT6), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n593_), .B1(new_n596_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT8), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT64), .B(G92gat), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT9), .B1(new_n603_), .B2(G85gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n605_));
  NOR2_X1   g404(.A1(G85gat), .A2(G92gat), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(new_n606_), .B2(KEYINPUT65), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(KEYINPUT65), .B2(new_n605_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n604_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT66), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(G106gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(KEYINPUT10), .B(G99gat), .Z(new_n613_));
  AOI21_X1  g412(.A(new_n599_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n602_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n592_), .B1(new_n615_), .B2(new_n560_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n590_), .B1(new_n616_), .B2(KEYINPUT69), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n616_), .B1(new_n562_), .B2(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI221_X1 g418(.A(new_n616_), .B1(KEYINPUT69), .B2(new_n590_), .C1(new_n562_), .C2(new_n615_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G190gat), .B(G218gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G134gat), .B(G162gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n621_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n626_), .B(KEYINPUT36), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT73), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n621_), .B2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n619_), .A2(KEYINPUT73), .A3(new_n620_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n629_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT74), .B(KEYINPUT37), .Z(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT75), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT75), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n635_), .A2(new_n639_), .A3(new_n636_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n629_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n621_), .A2(new_n630_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n638_), .A2(new_n640_), .B1(KEYINPUT37), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(G231gat), .A2(G233gat), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n557_), .B(new_n645_), .Z(new_n646_));
  XNOR2_X1  g445(.A(G57gat), .B(G64gat), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT11), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT11), .ZN(new_n649_));
  XOR2_X1   g448(.A(G71gat), .B(G78gat), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n646_), .B(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(G127gat), .B(G155gat), .Z(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT16), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G183gat), .B(G211gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT17), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n654_), .A2(new_n659_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(KEYINPUT76), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT17), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n654_), .A2(new_n662_), .A3(new_n658_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(KEYINPUT76), .ZN(new_n664_));
  INV_X1    g463(.A(new_n660_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT77), .B1(new_n644_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n653_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n611_), .A2(new_n614_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(new_n602_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n615_), .A2(new_n653_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT12), .A3(new_n671_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n615_), .A2(KEYINPUT12), .A3(new_n653_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(G230gat), .A2(G233gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT67), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n670_), .A2(new_n677_), .A3(new_n671_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n675_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n615_), .A2(KEYINPUT67), .A3(new_n653_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n676_), .A2(new_n681_), .ZN(new_n682_));
  XOR2_X1   g481(.A(G120gat), .B(G148gat), .Z(new_n683_));
  XNOR2_X1  g482(.A(G176gat), .B(G204gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n685_), .B(new_n686_), .Z(new_n687_));
  NAND2_X1  g486(.A1(new_n682_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n687_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n676_), .A2(new_n681_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT13), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n688_), .A2(KEYINPUT13), .A3(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n643_), .A2(KEYINPUT37), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n635_), .A2(new_n639_), .A3(new_n636_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n639_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT77), .ZN(new_n701_));
  INV_X1    g500(.A(new_n666_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n667_), .A2(new_n696_), .A3(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n585_), .A2(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n414_), .A2(KEYINPUT112), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n414_), .A2(KEYINPUT112), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n705_), .A2(new_n552_), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT38), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n550_), .A2(new_n635_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n695_), .A2(new_n582_), .A3(new_n666_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n414_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G1gat), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n710_), .A2(new_n711_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n712_), .A2(new_n717_), .A3(new_n718_), .ZN(G1324gat));
  NOR2_X1   g518(.A1(new_n332_), .A2(new_n423_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n585_), .A2(new_n704_), .A3(new_n553_), .A4(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G8gat), .B1(new_n715_), .B2(new_n720_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(KEYINPUT39), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(KEYINPUT39), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT40), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1325gat));
  OAI21_X1  g527(.A(G15gat), .B1(new_n715_), .B2(new_n549_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT41), .Z(new_n730_));
  INV_X1    g529(.A(G15gat), .ZN(new_n731_));
  INV_X1    g530(.A(new_n549_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n705_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1326gat));
  XNOR2_X1  g533(.A(new_n539_), .B(KEYINPUT113), .ZN(new_n735_));
  OAI21_X1  g534(.A(G22gat), .B1(new_n715_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT42), .ZN(new_n737_));
  INV_X1    g536(.A(G22gat), .ZN(new_n738_));
  INV_X1    g537(.A(new_n735_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n705_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(G1327gat));
  NAND2_X1  g540(.A1(new_n635_), .A2(new_n666_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n695_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G29gat), .B1(new_n745_), .B2(new_n414_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n695_), .A2(new_n582_), .A3(new_n702_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n547_), .A2(new_n549_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n504_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n750_), .B2(new_n644_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n550_), .A2(new_n700_), .A3(KEYINPUT43), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n747_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT114), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755_));
  INV_X1    g554(.A(new_n747_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n750_), .A2(new_n748_), .A3(new_n644_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n550_), .B2(new_n700_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n754_), .A2(new_n755_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(KEYINPUT44), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n709_), .A2(G29gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n746_), .B1(new_n764_), .B2(new_n765_), .ZN(G1328gat));
  XNOR2_X1  g565(.A(KEYINPUT115), .B(KEYINPUT46), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(G36gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n720_), .B1(new_n759_), .B2(KEYINPUT44), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n762_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n720_), .A2(G36gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n745_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n772_), .B1(new_n745_), .B2(new_n773_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n768_), .B1(new_n771_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n745_), .A2(new_n773_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT45), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n774_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n721_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT44), .B1(new_n753_), .B2(KEYINPUT114), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n761_), .B2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n781_), .B(new_n767_), .C1(new_n784_), .C2(new_n769_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n778_), .A2(new_n785_), .ZN(G1329gat));
  INV_X1    g585(.A(G43gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n755_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n753_), .A2(KEYINPUT114), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n763_), .B(new_n788_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n745_), .A2(new_n732_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n787_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT116), .B(KEYINPUT47), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n791_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1330gat));
  AOI21_X1  g598(.A(G50gat), .B1(new_n745_), .B2(new_n739_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n539_), .A2(G50gat), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n764_), .B2(new_n802_), .ZN(G1331gat));
  NOR2_X1   g602(.A1(new_n666_), .A2(new_n581_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NOR4_X1   g604(.A1(new_n550_), .A2(new_n696_), .A3(new_n635_), .A4(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(G57gat), .B1(new_n807_), .B2(new_n716_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n550_), .A2(new_n581_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n667_), .A2(new_n809_), .A3(new_n695_), .A4(new_n703_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n708_), .A2(G57gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n808_), .B1(new_n810_), .B2(new_n811_), .ZN(G1332gat));
  OR3_X1    g611(.A1(new_n810_), .A2(G64gat), .A3(new_n720_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n806_), .A2(new_n721_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT48), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n814_), .A2(new_n815_), .A3(G64gat), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n814_), .B2(G64gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT117), .ZN(G1333gat));
  OAI21_X1  g618(.A(G71gat), .B1(new_n807_), .B2(new_n549_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT49), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n549_), .A2(G71gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n810_), .B2(new_n822_), .ZN(G1334gat));
  OAI21_X1  g622(.A(G78gat), .B1(new_n807_), .B2(new_n735_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT50), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n735_), .A2(G78gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n810_), .B2(new_n826_), .ZN(G1335gat));
  INV_X1    g626(.A(G85gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n695_), .A2(new_n582_), .A3(new_n666_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n830_), .B2(new_n414_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n809_), .A2(new_n695_), .A3(new_n666_), .A4(new_n635_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n832_), .A2(G85gat), .A3(new_n708_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1336gat));
  INV_X1    g633(.A(new_n832_), .ZN(new_n835_));
  AOI21_X1  g634(.A(G92gat), .B1(new_n835_), .B2(new_n721_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n721_), .A2(new_n603_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(KEYINPUT118), .Z(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n830_), .B2(new_n838_), .ZN(G1337gat));
  NAND2_X1  g638(.A1(new_n830_), .A2(new_n732_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n459_), .A2(new_n613_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n840_), .A2(G99gat), .B1(new_n835_), .B2(new_n841_), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g642(.A1(new_n835_), .A2(new_n612_), .A3(new_n539_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n830_), .A2(new_n539_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(G106gat), .ZN(new_n847_));
  AOI211_X1 g646(.A(KEYINPUT52), .B(new_n612_), .C1(new_n830_), .C2(new_n539_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n844_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT53), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n851_), .B(new_n844_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1339gat));
  NOR2_X1   g652(.A1(new_n695_), .A2(new_n805_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n700_), .A2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT54), .ZN(new_n856_));
  INV_X1    g655(.A(new_n635_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n581_), .A2(new_n690_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n672_), .A2(new_n679_), .A3(new_n673_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n676_), .A2(KEYINPUT55), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n679_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n689_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n860_), .A2(KEYINPUT56), .A3(new_n863_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n858_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n564_), .B1(new_n563_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n869_), .B2(new_n563_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n574_), .B1(new_n569_), .B2(new_n564_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n579_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n857_), .B1(new_n868_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(KEYINPUT57), .B(new_n857_), .C1(new_n868_), .C2(new_n875_), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n690_), .A2(new_n579_), .A3(new_n873_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n867_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT56), .B1(new_n860_), .B2(new_n863_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n880_), .B(KEYINPUT58), .C1(new_n881_), .C2(new_n882_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n878_), .B(new_n879_), .C1(new_n700_), .C2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n666_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n539_), .B1(new_n856_), .B2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n708_), .A2(new_n721_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n459_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n890_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(G113gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n895_), .A2(new_n896_), .A3(new_n581_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n856_), .B2(new_n889_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(KEYINPUT59), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n894_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n890_), .B(new_n893_), .C1(new_n899_), .C2(KEYINPUT59), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n582_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n897_), .B1(new_n903_), .B2(new_n896_), .ZN(G1340gat));
  INV_X1    g703(.A(G120gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n696_), .B2(KEYINPUT60), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n895_), .B(new_n906_), .C1(KEYINPUT60), .C2(new_n905_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n696_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n905_), .ZN(G1341gat));
  NAND3_X1  g708(.A1(new_n895_), .A2(new_n339_), .A3(new_n702_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n666_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n339_), .ZN(G1342gat));
  AOI21_X1  g711(.A(G134gat), .B1(new_n895_), .B2(new_n635_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n901_), .A2(new_n902_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT121), .B(G134gat), .Z(new_n915_));
  NOR2_X1   g714(.A1(new_n700_), .A2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n913_), .B1(new_n914_), .B2(new_n916_), .ZN(G1343gat));
  NAND2_X1  g716(.A1(new_n549_), .A2(new_n539_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n856_), .B2(new_n889_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n919_), .A2(new_n581_), .A3(new_n891_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g720(.A1(new_n919_), .A2(new_n695_), .A3(new_n891_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g722(.A1(new_n856_), .A2(new_n889_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n918_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n924_), .A2(new_n702_), .A3(new_n891_), .A4(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n919_), .A2(KEYINPUT122), .A3(new_n702_), .A4(new_n891_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT61), .B(G155gat), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n928_), .A2(new_n929_), .A3(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1346gat));
  NAND2_X1  g732(.A1(new_n919_), .A2(new_n891_), .ZN(new_n934_));
  OAI21_X1  g733(.A(G162gat), .B1(new_n934_), .B2(new_n700_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n635_), .A2(new_n363_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n934_), .B2(new_n936_), .ZN(G1347gat));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n549_), .A2(new_n720_), .A3(new_n709_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT123), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n739_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n924_), .A2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n582_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n938_), .B1(new_n943_), .B2(new_n236_), .ZN(new_n944_));
  OAI211_X1 g743(.A(KEYINPUT62), .B(G169gat), .C1(new_n942_), .C2(new_n582_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n255_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n944_), .A2(new_n945_), .A3(new_n946_), .ZN(G1348gat));
  INV_X1    g746(.A(new_n942_), .ZN(new_n948_));
  AOI21_X1  g747(.A(G176gat), .B1(new_n948_), .B2(new_n695_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n950_));
  OR2_X1    g749(.A1(new_n890_), .A2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n890_), .A2(new_n950_), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n940_), .A2(new_n240_), .A3(new_n696_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n949_), .B1(new_n953_), .B2(new_n954_), .ZN(G1349gat));
  NOR3_X1   g754(.A1(new_n942_), .A2(new_n263_), .A3(new_n666_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n940_), .A2(new_n666_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n951_), .A2(new_n952_), .A3(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n956_), .B1(new_n958_), .B2(new_n248_), .ZN(G1350gat));
  OAI21_X1  g758(.A(G190gat), .B1(new_n942_), .B2(new_n700_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n635_), .A2(new_n264_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n942_), .B2(new_n961_), .ZN(G1351gat));
  NOR2_X1   g761(.A1(new_n720_), .A2(new_n414_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n919_), .A2(new_n581_), .A3(new_n963_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n964_), .B1(KEYINPUT125), .B2(new_n218_), .ZN(new_n965_));
  XOR2_X1   g764(.A(KEYINPUT125), .B(G197gat), .Z(new_n966_));
  AOI21_X1  g765(.A(new_n965_), .B1(new_n964_), .B2(new_n966_), .ZN(G1352gat));
  AND2_X1   g766(.A1(new_n919_), .A2(new_n963_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n695_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g769(.A(new_n666_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n971_));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n972_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n973_));
  OR3_X1    g772(.A1(new_n972_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974_));
  AOI22_X1  g773(.A1(new_n968_), .A2(new_n971_), .B1(new_n973_), .B2(new_n974_), .ZN(new_n975_));
  AND2_X1   g774(.A1(new_n968_), .A2(new_n971_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n975_), .B1(new_n976_), .B2(new_n974_), .ZN(G1354gat));
  AOI21_X1  g776(.A(G218gat), .B1(new_n968_), .B2(new_n635_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n644_), .A2(G218gat), .ZN(new_n979_));
  XNOR2_X1  g778(.A(new_n979_), .B(KEYINPUT127), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n978_), .B1(new_n968_), .B2(new_n980_), .ZN(G1355gat));
endmodule


