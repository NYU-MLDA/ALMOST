//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n966_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206_));
  INV_X1    g005(.A(G85gat), .ZN(new_n207_));
  INV_X1    g006(.A(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n206_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n206_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n205_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT10), .B(G99gat), .Z(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(KEYINPUT64), .B(new_n212_), .C1(new_n220_), .C2(new_n206_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n214_), .A2(new_n217_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT65), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT7), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n227_), .B2(new_n224_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT8), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n204_), .B1(new_n222_), .B2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n234_));
  INV_X1    g033(.A(new_n220_), .ZN(new_n235_));
  AOI211_X1 g034(.A(new_n235_), .B(new_n231_), .C1(new_n229_), .C2(new_n203_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n233_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G57gat), .B(G64gat), .Z(new_n238_));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G71gat), .B(G78gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n243_), .A3(KEYINPUT11), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n237_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(KEYINPUT12), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n237_), .A2(new_n249_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n245_), .A2(KEYINPUT12), .A3(new_n246_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n252_), .B1(new_n237_), .B2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G230gat), .ZN(new_n256_));
  INV_X1    g055(.A(G233gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n252_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n258_), .B1(new_n261_), .B2(new_n250_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G120gat), .B(G148gat), .ZN(new_n264_));
  INV_X1    g063(.A(G204gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT5), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT68), .B1(new_n263_), .B2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n271_), .A2(new_n272_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT13), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n271_), .A2(new_n272_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT13), .B1(new_n278_), .B2(new_n273_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G22gat), .B(G50gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT80), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT81), .B1(G141gat), .B2(G148gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT82), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n289_), .A2(KEYINPUT82), .A3(new_n290_), .A4(new_n291_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n287_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT3), .ZN(new_n298_));
  NAND3_X1  g097(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT79), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n298_), .B(new_n299_), .C1(new_n301_), .C2(KEYINPUT2), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n286_), .B1(new_n296_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n285_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n284_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT79), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n300_), .B(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n297_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n281_), .B1(new_n310_), .B2(KEYINPUT29), .ZN(new_n311_));
  AOI211_X1 g110(.A(new_n287_), .B(new_n301_), .C1(new_n284_), .C2(new_n305_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT2), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n308_), .A2(new_n313_), .B1(KEYINPUT3), .B2(new_n297_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n314_), .A2(new_n299_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n315_), .B2(new_n286_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317_));
  INV_X1    g116(.A(new_n281_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT83), .B(KEYINPUT28), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n311_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n311_), .B2(new_n319_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n321_), .A2(new_n322_), .A3(KEYINPUT87), .ZN(new_n323_));
  INV_X1    g122(.A(G228gat), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n324_), .A2(new_n257_), .A3(KEYINPUT86), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G211gat), .B(G218gat), .Z(new_n327_));
  INV_X1    g126(.A(G197gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n328_), .A2(G204gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(KEYINPUT84), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT84), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G197gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n329_), .B1(new_n333_), .B2(G204gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT21), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n327_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n330_), .A2(new_n332_), .A3(new_n265_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT85), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n265_), .B2(G197gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n328_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT21), .B1(new_n337_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n333_), .A2(G204gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n329_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n335_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n336_), .A2(new_n342_), .B1(new_n345_), .B2(new_n327_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n310_), .B2(KEYINPUT29), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT86), .B1(new_n324_), .B2(new_n257_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n326_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G78gat), .B(G106gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT84), .B(G197gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n344_), .B1(new_n352_), .B2(new_n265_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(KEYINPUT21), .A3(new_n327_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n335_), .B(new_n344_), .C1(new_n352_), .C2(new_n265_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n327_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n339_), .A2(new_n340_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n330_), .A2(new_n332_), .A3(new_n265_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n335_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n354_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n325_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n350_), .A2(new_n351_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n351_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n325_), .B1(new_n362_), .B2(new_n348_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n347_), .A2(new_n326_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n323_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n364_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n311_), .A2(new_n319_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n320_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n311_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT87), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n377_), .A3(new_n374_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n351_), .B1(new_n350_), .B2(new_n363_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n369_), .A2(new_n376_), .A3(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  XNOR2_X1  g183(.A(G15gat), .B(G43gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT31), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G127gat), .B(G134gat), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n388_), .A2(G113gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(G113gat), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n389_), .A2(G120gat), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(G120gat), .B1(new_n389_), .B2(new_n390_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT23), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n395_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT78), .B(G176gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n400_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT30), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT25), .B(G183gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT26), .B(G190gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(G169gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n268_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n413_), .A2(KEYINPUT24), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(KEYINPUT24), .A3(new_n394_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n411_), .A2(new_n397_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n407_), .A2(new_n408_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n408_), .B1(new_n407_), .B2(new_n416_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n393_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n407_), .A2(new_n416_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT30), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n391_), .A2(new_n392_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n417_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n387_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n420_), .A2(new_n424_), .A3(new_n387_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n384_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n427_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n384_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n429_), .A2(new_n425_), .A3(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n381_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n310_), .A2(new_n393_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n423_), .A2(new_n303_), .A3(new_n309_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(KEYINPUT4), .A3(new_n435_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n437_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n310_), .A2(new_n393_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G1gat), .B(G29gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G57gat), .B(G85gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n438_), .A2(new_n443_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT92), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT33), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n438_), .A2(new_n443_), .A3(new_n452_), .A4(new_n448_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT93), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n449_), .A2(new_n451_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n457_), .B(KEYINPUT88), .Z(new_n458_));
  XOR2_X1   g257(.A(new_n458_), .B(KEYINPUT19), .Z(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n405_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n403_), .A2(KEYINPUT89), .A3(new_n404_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n401_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n396_), .B(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n394_), .B1(new_n466_), .B2(new_n398_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n416_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT20), .B1(new_n361_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n342_), .A2(new_n356_), .A3(new_n355_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n470_), .A2(new_n354_), .B1(new_n407_), .B2(new_n416_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n460_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n361_), .A2(new_n468_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n470_), .A2(new_n407_), .A3(new_n416_), .A4(new_n354_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(KEYINPUT20), .A4(new_n459_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G8gat), .B(G36gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G64gat), .B(G92gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n472_), .A2(new_n475_), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n436_), .A2(new_n440_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n439_), .A2(new_n437_), .A3(new_n442_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n448_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n456_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n450_), .A2(new_n490_), .A3(new_n451_), .A4(new_n453_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n455_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  AND4_X1   g291(.A1(KEYINPUT20), .A2(new_n473_), .A3(new_n474_), .A4(new_n460_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n411_), .A2(new_n397_), .A3(new_n415_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n403_), .A2(KEYINPUT89), .A3(new_n404_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT89), .B1(new_n403_), .B2(new_n404_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n402_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n495_), .A2(new_n414_), .B1(new_n498_), .B2(new_n400_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n494_), .B1(new_n346_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n421_), .A2(new_n361_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n460_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(KEYINPUT32), .B(new_n480_), .C1(new_n493_), .C2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n503_), .B(KEYINPUT94), .Z(new_n504_));
  AOI21_X1  g303(.A(new_n448_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n449_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n472_), .A2(new_n475_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT32), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n508_), .B1(new_n509_), .B2(new_n481_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n504_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n433_), .B1(new_n492_), .B2(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n370_), .A2(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n432_), .B1(new_n513_), .B2(new_n369_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT98), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n459_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n516_));
  AND4_X1   g315(.A1(KEYINPUT20), .A2(new_n473_), .A3(new_n474_), .A4(new_n459_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n480_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT97), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n480_), .B(KEYINPUT96), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n520_), .B1(new_n493_), .B2(new_n502_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT97), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n483_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT27), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n482_), .A2(new_n483_), .A3(KEYINPUT27), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n515_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  AOI211_X1 g327(.A(KEYINPUT98), .B(new_n526_), .C1(new_n524_), .C2(KEYINPUT27), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n514_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n428_), .A2(new_n431_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n381_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n526_), .B1(new_n524_), .B2(KEYINPUT27), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n507_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n506_), .A2(KEYINPUT95), .A3(new_n449_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n512_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G1gat), .B(G8gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT74), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544_));
  INV_X1    g343(.A(G1gat), .ZN(new_n545_));
  INV_X1    g344(.A(G8gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n543_), .A2(new_n548_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(G43gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT69), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT69), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G43gat), .ZN(new_n555_));
  INV_X1    g354(.A(G50gat), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n553_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n556_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G29gat), .B(G36gat), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n553_), .A2(new_n555_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(G50gat), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n564_), .B2(new_n557_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n551_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n551_), .A2(new_n567_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT15), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n573_), .B1(new_n561_), .B2(new_n565_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n560_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n564_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(KEYINPUT15), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n572_), .B1(new_n551_), .B2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n571_), .B1(new_n570_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G113gat), .B(G141gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(new_n412_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n328_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n580_), .B(new_n583_), .Z(new_n584_));
  NOR2_X1   g383(.A1(new_n541_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT99), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n541_), .B2(new_n584_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n280_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT71), .B(G134gat), .ZN(new_n590_));
  INV_X1    g389(.A(G162gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n222_), .A2(new_n232_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n234_), .B1(new_n598_), .B2(new_n203_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n236_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n578_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT70), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT35), .B(new_n597_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n599_), .A2(new_n567_), .A3(new_n600_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n597_), .A2(KEYINPUT35), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n604_), .B(new_n606_), .C1(new_n578_), .C2(new_n237_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n578_), .B2(new_n237_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n603_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n595_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT72), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n603_), .A2(new_n607_), .ZN(new_n613_));
  NOR4_X1   g412(.A1(new_n233_), .A2(new_n236_), .A3(new_n566_), .A4(new_n234_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n601_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT70), .B1(new_n237_), .B2(new_n578_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n615_), .A2(KEYINPUT35), .A3(new_n597_), .A4(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n594_), .B(KEYINPUT36), .Z(new_n618_));
  NAND3_X1  g417(.A1(new_n613_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT72), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n620_), .B(new_n595_), .C1(new_n608_), .C2(new_n610_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n612_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(KEYINPUT73), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT37), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n624_), .A2(new_n619_), .A3(new_n612_), .A4(new_n621_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n551_), .B(new_n630_), .Z(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(new_n249_), .Z(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT16), .B(G183gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(G211gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT17), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n631_), .B(new_n247_), .ZN(new_n638_));
  XOR2_X1   g437(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT76), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n632_), .A2(new_n637_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT77), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n629_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n589_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n540_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n545_), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT38), .ZN(new_n649_));
  INV_X1    g448(.A(new_n622_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n644_), .A2(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n277_), .A2(new_n279_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n585_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n540_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n649_), .A2(new_n654_), .ZN(G1324gat));
  NOR2_X1   g454(.A1(new_n528_), .A2(new_n529_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G8gat), .B1(new_n653_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT39), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n646_), .A2(new_n546_), .A3(new_n656_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g463(.A(G15gat), .B1(new_n653_), .B2(new_n432_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT41), .Z(new_n666_));
  INV_X1    g465(.A(G15gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n646_), .A2(new_n667_), .A3(new_n531_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1326gat));
  XOR2_X1   g468(.A(new_n381_), .B(KEYINPUT101), .Z(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G22gat), .B1(new_n653_), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT42), .ZN(new_n673_));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n646_), .A2(new_n674_), .A3(new_n670_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT102), .Z(G1327gat));
  NOR2_X1   g476(.A1(new_n643_), .A2(new_n622_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n589_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n647_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n682_));
  INV_X1    g481(.A(new_n584_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n644_), .B(new_n683_), .C1(new_n277_), .C2(new_n279_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n622_), .A2(new_n625_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n685_), .A2(KEYINPUT103), .A3(new_n627_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT103), .B1(new_n685_), .B2(new_n627_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n688_), .B2(new_n541_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n685_), .A2(new_n690_), .A3(new_n627_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n370_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n321_), .A2(new_n322_), .ZN(new_n693_));
  OAI22_X1  g492(.A1(new_n323_), .A2(new_n368_), .B1(new_n693_), .B2(new_n364_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n531_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT27), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n522_), .B1(new_n508_), .B2(new_n480_), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT97), .B(new_n481_), .C1(new_n472_), .C2(new_n475_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n696_), .B1(new_n699_), .B2(new_n521_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT98), .B1(new_n700_), .B2(new_n526_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n533_), .A2(new_n515_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n695_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n381_), .A2(new_n533_), .A3(new_n531_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n540_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n492_), .A2(new_n511_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n433_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n691_), .B1(new_n705_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n684_), .B1(new_n689_), .B2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n682_), .B1(new_n711_), .B2(KEYINPUT44), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n647_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n713_));
  OAI22_X1  g512(.A1(new_n686_), .A2(new_n687_), .B1(new_n713_), .B2(new_n512_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n709_), .B1(new_n714_), .B2(KEYINPUT43), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716_));
  NOR4_X1   g515(.A1(new_n715_), .A2(KEYINPUT104), .A3(new_n716_), .A4(new_n684_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n712_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(new_n540_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n711_), .A2(KEYINPUT44), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n681_), .B1(new_n720_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(new_n684_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n726_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n685_), .A2(KEYINPUT103), .A3(new_n627_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n705_), .A2(new_n708_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n690_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n725_), .B1(new_n731_), .B2(new_n709_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n657_), .B1(new_n732_), .B2(new_n716_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n733_), .B1(new_n712_), .B2(new_n717_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT105), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(new_n733_), .C1(new_n712_), .C2(new_n717_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n735_), .A2(G36gat), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT106), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n735_), .A2(new_n740_), .A3(G36gat), .A4(new_n737_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n657_), .A2(G36gat), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT107), .B1(new_n679_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n589_), .A2(new_n745_), .A3(new_n678_), .A4(new_n742_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n744_), .A2(KEYINPUT45), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT45), .B1(new_n744_), .B2(new_n746_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n739_), .A2(new_n741_), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT46), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT46), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n750_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1329gat));
  NAND4_X1  g555(.A1(new_n718_), .A2(G43gat), .A3(new_n531_), .A4(new_n722_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT109), .B(G43gat), .Z(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n679_), .B2(new_n432_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g560(.A(G50gat), .B1(new_n680_), .B2(new_n670_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n719_), .A2(new_n381_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n721_), .A2(new_n556_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n763_), .B2(new_n764_), .ZN(G1331gat));
  NAND4_X1  g564(.A1(new_n280_), .A2(new_n730_), .A3(new_n651_), .A4(new_n584_), .ZN(new_n766_));
  INV_X1    g565(.A(G57gat), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n540_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n730_), .A2(new_n584_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT110), .Z(new_n770_));
  NOR2_X1   g569(.A1(new_n770_), .A2(new_n652_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n647_), .A3(new_n645_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n768_), .B1(new_n772_), .B2(new_n767_), .ZN(G1332gat));
  OAI21_X1  g572(.A(G64gat), .B1(new_n766_), .B2(new_n657_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT48), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n771_), .A2(new_n645_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n657_), .A2(G64gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(G1333gat));
  OAI21_X1  g577(.A(G71gat), .B1(new_n766_), .B2(new_n432_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT49), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n432_), .A2(G71gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n776_), .B2(new_n781_), .ZN(G1334gat));
  OAI21_X1  g581(.A(G78gat), .B1(new_n766_), .B2(new_n671_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT111), .Z(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT50), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n671_), .A2(G78gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n776_), .B2(new_n786_), .ZN(G1335gat));
  OR4_X1    g586(.A1(new_n643_), .A2(new_n715_), .A3(new_n652_), .A4(new_n683_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n788_), .A2(new_n207_), .A3(new_n540_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n771_), .A2(new_n678_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n647_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n791_), .B2(new_n207_), .ZN(G1336gat));
  AOI21_X1  g591(.A(G92gat), .B1(new_n790_), .B2(new_n656_), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT112), .Z(new_n794_));
  NAND2_X1  g593(.A1(new_n656_), .A2(G92gat), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT113), .Z(new_n796_));
  NOR2_X1   g595(.A1(new_n788_), .A2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n794_), .A2(new_n797_), .ZN(G1337gat));
  NAND3_X1  g597(.A1(new_n790_), .A2(new_n215_), .A3(new_n531_), .ZN(new_n799_));
  OAI21_X1  g598(.A(G99gat), .B1(new_n788_), .B2(new_n432_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g601(.A(new_n381_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n790_), .A2(new_n216_), .A3(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT114), .ZN(new_n805_));
  OAI21_X1  g604(.A(G106gat), .B1(new_n788_), .B2(new_n381_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT52), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT53), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n805_), .A2(new_n810_), .A3(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1339gat));
  NAND3_X1  g611(.A1(new_n652_), .A2(new_n645_), .A3(new_n584_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT54), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n258_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT55), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n260_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n255_), .A2(KEYINPUT55), .A3(new_n259_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n269_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n815_), .B1(new_n820_), .B2(KEYINPUT115), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n251_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(KEYINPUT55), .B2(new_n816_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n819_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n270_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(KEYINPUT56), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n263_), .A2(new_n270_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n584_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n821_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n580_), .A2(new_n583_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n568_), .A2(new_n569_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n583_), .C1(new_n569_), .C2(new_n579_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n278_), .A2(new_n273_), .A3(new_n833_), .A4(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n821_), .A2(new_n827_), .A3(KEYINPUT116), .A4(new_n829_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n832_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n622_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT57), .B1(new_n838_), .B2(new_n622_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n833_), .A2(new_n835_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n825_), .B2(KEYINPUT56), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n828_), .B1(new_n820_), .B2(new_n815_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n843_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n848_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n845_), .A2(new_n846_), .A3(KEYINPUT117), .A4(KEYINPUT58), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n629_), .A4(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n841_), .A2(new_n842_), .A3(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n814_), .B1(new_n854_), .B2(new_n643_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n703_), .A2(new_n647_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  XOR2_X1   g658(.A(new_n813_), .B(KEYINPUT54), .Z(new_n860_));
  NAND2_X1  g659(.A1(new_n839_), .A2(new_n840_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(KEYINPUT119), .A3(new_n852_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n842_), .B2(new_n853_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n841_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n862_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n860_), .B1(new_n866_), .B2(new_n644_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n857_), .B(KEYINPUT118), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n859_), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n858_), .A2(new_n859_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G113gat), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n584_), .ZN(new_n872_));
  AOI21_X1  g671(.A(G113gat), .B1(new_n858_), .B2(new_n683_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1340gat));
  OAI21_X1  g673(.A(G120gat), .B1(new_n870_), .B2(new_n652_), .ZN(new_n875_));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n652_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n858_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n876_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(G1341gat));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n870_), .A2(new_n880_), .A3(new_n644_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G127gat), .B1(new_n858_), .B2(new_n643_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1342gat));
  INV_X1    g682(.A(G134gat), .ZN(new_n884_));
  INV_X1    g683(.A(new_n629_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n870_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G134gat), .B1(new_n858_), .B2(new_n650_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1343gat));
  NOR2_X1   g687(.A1(new_n856_), .A2(new_n540_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n656_), .A2(new_n531_), .A3(new_n381_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n584_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT120), .B(G141gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1344gat));
  INV_X1    g693(.A(new_n891_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n280_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n643_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT61), .B(G155gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1346gat));
  NOR3_X1   g699(.A1(new_n891_), .A2(new_n591_), .A3(new_n688_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n895_), .A2(new_n650_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n591_), .B2(new_n902_), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n657_), .A2(new_n647_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n531_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n867_), .A2(new_n670_), .A3(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n905_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n842_), .A2(new_n853_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n841_), .B1(new_n910_), .B2(KEYINPUT119), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n643_), .B1(new_n911_), .B2(new_n864_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n671_), .B(new_n909_), .C1(new_n912_), .C2(new_n860_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT121), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n908_), .A2(new_n914_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n915_), .B(new_n683_), .C1(new_n497_), .C2(new_n496_), .ZN(new_n916_));
  AOI211_X1 g715(.A(KEYINPUT62), .B(new_n412_), .C1(new_n906_), .C2(new_n683_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n906_), .A2(new_n683_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(G169gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n916_), .B1(new_n917_), .B2(new_n920_), .ZN(G1348gat));
  NAND3_X1  g720(.A1(new_n855_), .A2(new_n381_), .A3(new_n909_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n922_), .A2(new_n268_), .A3(new_n652_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n915_), .A2(new_n280_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(new_n402_), .ZN(G1349gat));
  NOR2_X1   g724(.A1(new_n644_), .A2(new_n409_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n906_), .A2(new_n907_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n913_), .A2(KEYINPUT121), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n922_), .A2(new_n644_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(G183gat), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n929_), .A2(new_n930_), .A3(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n926_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n908_), .B2(new_n914_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT122), .B1(new_n936_), .B2(new_n932_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n937_), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n915_), .A2(new_n650_), .A3(new_n410_), .ZN(new_n939_));
  INV_X1    g738(.A(G190gat), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n885_), .B1(new_n908_), .B2(new_n914_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n939_), .B1(new_n940_), .B2(new_n941_), .ZN(G1351gat));
  AND2_X1   g741(.A1(new_n855_), .A2(new_n532_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n904_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n584_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(new_n328_), .ZN(G1352gat));
  NAND3_X1  g745(.A1(new_n943_), .A2(new_n280_), .A3(new_n904_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n947_), .B1(KEYINPUT123), .B2(G204gat), .ZN(new_n948_));
  NAND2_X1  g747(.A1(KEYINPUT123), .A2(G204gat), .ZN(new_n949_));
  MUX2_X1   g748(.A(new_n947_), .B(new_n948_), .S(new_n949_), .Z(G1353gat));
  NAND4_X1  g749(.A1(new_n855_), .A2(new_n643_), .A3(new_n532_), .A4(new_n904_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  AND2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  OR3_X1    g752(.A1(new_n951_), .A2(new_n952_), .A3(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n951_), .A2(new_n955_), .A3(new_n952_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(new_n951_), .B2(new_n952_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n954_), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(KEYINPUT125), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n960_));
  OAI211_X1 g759(.A(new_n954_), .B(new_n960_), .C1(new_n957_), .C2(new_n956_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n959_), .A2(new_n961_), .ZN(G1354gat));
  XOR2_X1   g761(.A(KEYINPUT127), .B(G218gat), .Z(new_n963_));
  NOR3_X1   g762(.A1(new_n944_), .A2(new_n885_), .A3(new_n963_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n943_), .A2(new_n650_), .A3(new_n904_), .ZN(new_n965_));
  XOR2_X1   g764(.A(new_n965_), .B(KEYINPUT126), .Z(new_n966_));
  AOI21_X1  g765(.A(new_n964_), .B1(new_n966_), .B2(new_n963_), .ZN(G1355gat));
endmodule


