//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT73), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n205_), .B(KEYINPUT15), .Z(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT10), .B(G99gat), .Z(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G106gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT9), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT6), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT9), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n211_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  OR3_X1    g025(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(new_n212_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT8), .B1(new_n212_), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n229_), .B(new_n231_), .Z(new_n232_));
  NAND4_X1  g031(.A1(new_n211_), .A2(new_n221_), .A3(KEYINPUT67), .A4(new_n222_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n225_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n206_), .A2(new_n234_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n225_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n205_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT34), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT35), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT74), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n235_), .A2(new_n238_), .A3(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n241_), .A2(new_n242_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n245_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n235_), .A2(new_n238_), .A3(new_n247_), .A4(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G190gat), .B(G218gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G134gat), .B(G162gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n249_), .A2(KEYINPUT36), .A3(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(KEYINPUT36), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n255_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT37), .ZN(new_n257_));
  NOR3_X1   g056(.A1(new_n253_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n249_), .A2(KEYINPUT75), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n255_), .B1(new_n249_), .B2(KEYINPUT75), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n253_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n258_), .B1(new_n263_), .B2(new_n257_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT76), .B(G15gat), .ZN(new_n265_));
  INV_X1    g064(.A(G22gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G1gat), .ZN(new_n268_));
  INV_X1    g067(.A(G8gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT14), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G1gat), .B(G8gat), .Z(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n271_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n271_), .B(new_n272_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n275_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(G231gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G57gat), .B(G64gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G71gat), .B(G78gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n286_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n282_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n282_), .A2(new_n292_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G127gat), .B(G155gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(G183gat), .B(G211gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT17), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n299_), .A2(KEYINPUT71), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n299_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(KEYINPUT17), .B2(new_n303_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n293_), .A2(new_n294_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n301_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n264_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT80), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT23), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(G183gat), .A3(G190gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G169gat), .ZN(new_n316_));
  INV_X1    g115(.A(G176gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT24), .A3(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n315_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n325_));
  INV_X1    g124(.A(G183gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(KEYINPUT83), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n325_), .B(KEYINPUT25), .C1(new_n326_), .C2(KEYINPUT83), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT84), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(KEYINPUT82), .A2(KEYINPUT25), .A3(G183gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n329_), .A2(new_n330_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT26), .ZN(new_n335_));
  INV_X1    g134(.A(G190gat), .ZN(new_n336_));
  OAI211_X1 g135(.A(KEYINPUT84), .B(new_n335_), .C1(new_n336_), .C2(KEYINPUT85), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT85), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G190gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n335_), .B1(new_n340_), .B2(KEYINPUT84), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n324_), .B1(new_n334_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n311_), .A2(new_n313_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n344_), .B(new_n345_), .C1(G183gat), .C2(G190gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT22), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n346_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n343_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(G71gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(G99gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n351_), .B(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G127gat), .B(G134gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT87), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G113gat), .B(G120gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G15gat), .B(G43gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT86), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT30), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n362_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n358_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n370_));
  INV_X1    g169(.A(G197gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n370_), .B1(new_n371_), .B2(G204gat), .ZN(new_n372_));
  INV_X1    g171(.A(G204gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(G204gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT21), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n371_), .B2(G204gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n373_), .A2(KEYINPUT92), .A3(G197gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT21), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .A4(new_n375_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n377_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n381_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n379_), .A2(new_n375_), .A3(new_n380_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(G141gat), .ZN(new_n394_));
  INV_X1    g193(.A(G148gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(KEYINPUT3), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(G141gat), .B2(G148gat), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G141gat), .A2(G148gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT2), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT89), .B1(new_n399_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n396_), .A2(new_n398_), .ZN(new_n406_));
  AND3_X1   g205(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT89), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n393_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n391_), .B1(KEYINPUT1), .B2(new_n389_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(KEYINPUT1), .B2(new_n389_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G141gat), .A2(G148gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n414_), .A2(new_n416_), .A3(new_n400_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT90), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n406_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n410_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n392_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n414_), .A2(new_n416_), .A3(new_n400_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n369_), .B(new_n388_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n412_), .A2(new_n417_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n388_), .B1(new_n428_), .B2(new_n426_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(G228gat), .A3(G233gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G78gat), .B(G106gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n427_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n425_), .A2(new_n426_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT28), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT28), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n425_), .A2(new_n438_), .A3(new_n426_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G22gat), .B(G50gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n437_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n438_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n443_));
  AOI211_X1 g242(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n418_), .C2(new_n424_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n442_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT93), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n441_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n441_), .B2(new_n445_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n434_), .B(new_n435_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n441_), .A2(new_n445_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n450_), .A2(KEYINPUT93), .B1(new_n434_), .B2(new_n435_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G1gat), .B(G29gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G57gat), .B(G85gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n361_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n360_), .B(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n418_), .A2(new_n424_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n428_), .A2(new_n362_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n458_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(KEYINPUT4), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n461_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n465_), .B1(new_n469_), .B2(new_n464_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G226gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT19), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT20), .B1(new_n351_), .B2(new_n388_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n382_), .A2(new_n383_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n474_), .A2(new_n377_), .B1(new_n386_), .B2(new_n385_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n319_), .B(KEYINPUT95), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n316_), .A2(KEYINPUT22), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n348_), .A2(G169gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n317_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n346_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT96), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n346_), .A2(new_n476_), .A3(KEYINPUT96), .A4(new_n479_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT25), .B(G183gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT26), .B(G190gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n485_), .A2(new_n486_), .B1(new_n487_), .B2(new_n321_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n318_), .A2(new_n319_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n489_), .A2(new_n487_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n490_), .A3(new_n315_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n475_), .B1(new_n484_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n472_), .B1(new_n473_), .B2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G8gat), .B(G36gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G64gat), .B(G92gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n351_), .A2(new_n388_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n484_), .A2(new_n475_), .A3(new_n491_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n472_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT20), .A4(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n493_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT98), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n493_), .A2(KEYINPUT98), .A3(new_n503_), .A4(new_n499_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n343_), .A2(new_n350_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n509_), .B2(new_n475_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n484_), .A2(new_n491_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n388_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n502_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  AND4_X1   g312(.A1(KEYINPUT20), .A2(new_n500_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n498_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n506_), .A2(new_n507_), .A3(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n470_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n464_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n468_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n467_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n458_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n461_), .A2(new_n464_), .A3(new_n462_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT100), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT100), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n461_), .A2(new_n462_), .A3(new_n525_), .A4(new_n464_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .A4(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT33), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(new_n526_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n531_), .A2(KEYINPUT33), .A3(new_n522_), .A4(new_n521_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n517_), .A2(new_n529_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT103), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n464_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n458_), .B1(new_n535_), .B2(new_n530_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n527_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n499_), .A2(KEYINPUT32), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n491_), .A2(new_n480_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n539_), .B1(new_n540_), .B2(new_n388_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n541_), .A2(KEYINPUT102), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n500_), .B1(new_n541_), .B2(KEYINPUT102), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n472_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n510_), .A2(new_n502_), .A3(new_n512_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n538_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n513_), .A2(new_n514_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n547_), .B2(new_n538_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n534_), .B1(new_n537_), .B2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n533_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n537_), .A2(new_n534_), .A3(new_n548_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n453_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n536_), .A2(new_n527_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT27), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n544_), .A2(new_n545_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n498_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n504_), .A2(KEYINPUT27), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n554_), .A2(new_n516_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n434_), .A2(new_n435_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n440_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n443_), .A2(new_n444_), .A3(new_n442_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT93), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n441_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n559_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n553_), .B(new_n558_), .C1(new_n564_), .C2(new_n451_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT104), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n453_), .A2(KEYINPUT104), .A3(new_n558_), .A4(new_n553_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n368_), .B1(new_n552_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n453_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n571_), .A2(new_n558_), .A3(new_n553_), .A4(new_n367_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G120gat), .B(G148gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT69), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n234_), .B2(new_n292_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n229_), .B(new_n231_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n224_), .B2(new_n223_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n583_), .A2(KEYINPUT69), .A3(new_n291_), .A4(new_n233_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n581_), .B(new_n584_), .C1(new_n291_), .C2(new_n236_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT70), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n292_), .B1(new_n234_), .B2(KEYINPUT12), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT71), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT12), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n583_), .B2(new_n233_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n234_), .A2(new_n591_), .A3(KEYINPUT12), .A4(new_n291_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n587_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n589_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n586_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n579_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n585_), .A2(new_n588_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT70), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n602_), .A2(new_n597_), .A3(new_n589_), .A4(new_n578_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT13), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G229gat), .A2(G233gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n280_), .A2(new_n237_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n280_), .A2(new_n237_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n608_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n276_), .A2(new_n279_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n206_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n609_), .A3(new_n607_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT81), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G169gat), .B(G197gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n620_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(new_n615_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n606_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n573_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n310_), .A2(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n628_), .A2(G1gat), .A3(new_n553_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT105), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT38), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT38), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n308_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n573_), .A2(new_n263_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT106), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n573_), .A2(new_n636_), .A3(new_n263_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n633_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n639_), .B2(new_n553_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n631_), .A2(new_n632_), .A3(new_n640_), .ZN(G1324gat));
  INV_X1    g440(.A(new_n628_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n558_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n269_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n269_), .B1(new_n638_), .B2(new_n643_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n644_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(G1325gat));
  INV_X1    g450(.A(G15gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n638_), .B2(new_n367_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT41), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n642_), .A2(new_n652_), .A3(new_n367_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1326gat));
  AOI21_X1  g455(.A(new_n266_), .B1(new_n638_), .B2(new_n453_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT42), .Z(new_n658_));
  NAND3_X1  g457(.A1(new_n642_), .A2(new_n266_), .A3(new_n453_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1327gat));
  NOR2_X1   g459(.A1(new_n263_), .A2(new_n308_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n573_), .A2(new_n626_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  OR3_X1    g462(.A1(new_n663_), .A2(G29gat), .A3(new_n553_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n626_), .A2(new_n307_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  INV_X1    g466(.A(new_n264_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n573_), .B2(new_n668_), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT43), .B(new_n264_), .C1(new_n570_), .C2(new_n572_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT44), .B(new_n666_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n537_), .A3(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n675_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT107), .B1(new_n675_), .B2(G29gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n664_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT108), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(new_n664_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1328gat));
  NOR2_X1   g481(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n558_), .A2(G36gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n662_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n684_), .B1(new_n662_), .B2(new_n685_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT45), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n688_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT45), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n686_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n683_), .B1(new_n689_), .B2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n673_), .A2(new_n643_), .A3(new_n674_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1329gat));
  AND2_X1   g497(.A1(new_n673_), .A2(new_n674_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(G43gat), .A3(new_n367_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G43gat), .B1(new_n662_), .B2(new_n367_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g503(.A(G50gat), .B1(new_n662_), .B2(new_n453_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n453_), .A2(G50gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n699_), .B2(new_n706_), .ZN(G1331gat));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n604_), .B(KEYINPUT13), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n624_), .B(new_n709_), .C1(new_n570_), .C2(new_n572_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n310_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n708_), .B1(new_n711_), .B2(new_n553_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT111), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n307_), .A2(new_n624_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n606_), .A2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n553_), .A2(new_n708_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(G1332gat));
  INV_X1    g517(.A(new_n711_), .ZN(new_n719_));
  INV_X1    g518(.A(G64gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n643_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n716_), .A2(new_n643_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(G64gat), .ZN(new_n724_));
  AOI211_X1 g523(.A(KEYINPUT48), .B(new_n720_), .C1(new_n716_), .C2(new_n643_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(G1333gat));
  NAND3_X1  g525(.A1(new_n719_), .A2(new_n353_), .A3(new_n367_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n716_), .A2(new_n367_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(G71gat), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G71gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1334gat));
  INV_X1    g531(.A(G78gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n719_), .A2(new_n733_), .A3(new_n453_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n716_), .A2(new_n453_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G78gat), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT50), .B(new_n733_), .C1(new_n716_), .C2(new_n453_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1335gat));
  AND2_X1   g538(.A1(new_n710_), .A2(new_n661_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n537_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n669_), .A2(new_n670_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n709_), .A2(new_n308_), .A3(new_n624_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n537_), .A2(G85gat), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT113), .Z(new_n746_));
  AOI21_X1  g545(.A(new_n741_), .B1(new_n744_), .B2(new_n746_), .ZN(G1336gat));
  NAND2_X1  g546(.A1(new_n742_), .A2(new_n743_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G92gat), .B1(new_n748_), .B2(new_n558_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n740_), .A2(new_n216_), .A3(new_n643_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1337gat));
  AND4_X1   g550(.A1(new_n207_), .A2(new_n710_), .A3(new_n367_), .A4(new_n661_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n752_), .A2(KEYINPUT114), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(KEYINPUT114), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n753_), .A2(new_n754_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n755_));
  OR2_X1    g554(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n756_));
  OAI21_X1  g555(.A(G99gat), .B1(new_n748_), .B2(new_n368_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1338gat));
  OAI21_X1  g559(.A(G106gat), .B1(new_n748_), .B2(new_n571_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(KEYINPUT116), .A3(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n764_));
  OAI211_X1 g563(.A(G106gat), .B(new_n764_), .C1(new_n748_), .C2(new_n571_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n740_), .A2(new_n208_), .A3(new_n453_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT53), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n763_), .A2(new_n769_), .A3(new_n765_), .A4(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1339gat));
  INV_X1    g570(.A(KEYINPUT57), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n607_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT119), .A3(new_n620_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT119), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n613_), .A2(new_n205_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n608_), .B1(new_n776_), .B2(new_n609_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n775_), .B1(new_n777_), .B2(new_n622_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n614_), .A2(new_n609_), .A3(new_n608_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n774_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n623_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n600_), .B2(new_n603_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n624_), .A2(new_n603_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n594_), .A2(new_n587_), .A3(new_n596_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n234_), .A2(new_n591_), .A3(KEYINPUT12), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT12), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n583_), .A2(new_n788_), .A3(new_n233_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(new_n292_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n588_), .B1(new_n790_), .B2(new_n595_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT55), .B(new_n588_), .C1(new_n790_), .C2(new_n595_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n786_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n784_), .B1(new_n795_), .B2(new_n579_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n783_), .B1(new_n796_), .B2(KEYINPUT118), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n597_), .A2(KEYINPUT55), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n791_), .A2(new_n792_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n785_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n578_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n784_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n782_), .B1(new_n797_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n253_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n772_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n796_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n795_), .A2(new_n784_), .A3(new_n579_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n603_), .A2(new_n623_), .A3(new_n780_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n807_), .A2(new_n809_), .A3(KEYINPUT58), .A4(new_n808_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n668_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n604_), .A2(new_n623_), .A3(new_n780_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n800_), .C2(new_n578_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n624_), .A2(new_n603_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n795_), .A2(new_n579_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n819_), .B2(KEYINPUT118), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n815_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(KEYINPUT57), .A4(new_n263_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n806_), .A2(new_n814_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n797_), .A2(new_n803_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n805_), .B1(new_n825_), .B2(new_n815_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n822_), .B1(new_n826_), .B2(KEYINPUT57), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n307_), .B1(new_n824_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n258_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n714_), .B(new_n829_), .C1(KEYINPUT37), .C2(new_n805_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT117), .B1(new_n830_), .B2(new_n606_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n709_), .A2(new_n832_), .A3(new_n264_), .A4(new_n714_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(KEYINPUT54), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT117), .B(new_n835_), .C1(new_n830_), .C2(new_n606_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n828_), .A2(new_n838_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n453_), .A2(new_n643_), .A3(new_n553_), .A4(new_n368_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n625_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843_));
  OR3_X1    g642(.A1(new_n842_), .A2(new_n843_), .A3(G113gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n842_), .B2(G113gat), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n841_), .B(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n624_), .A2(G113gat), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n844_), .A2(new_n845_), .B1(new_n847_), .B2(new_n848_), .ZN(G1340gat));
  XNOR2_X1  g648(.A(new_n841_), .B(KEYINPUT59), .ZN(new_n850_));
  OAI21_X1  g649(.A(G120gat), .B1(new_n850_), .B2(new_n709_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n841_), .ZN(new_n852_));
  INV_X1    g651(.A(G120gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n709_), .B2(KEYINPUT60), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n852_), .B(new_n854_), .C1(KEYINPUT60), .C2(new_n853_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n855_), .ZN(G1341gat));
  OAI21_X1  g655(.A(G127gat), .B1(new_n850_), .B2(new_n307_), .ZN(new_n857_));
  OR3_X1    g656(.A1(new_n841_), .A2(G127gat), .A3(new_n307_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1342gat));
  OAI21_X1  g658(.A(G134gat), .B1(new_n850_), .B2(new_n264_), .ZN(new_n860_));
  OR3_X1    g659(.A1(new_n841_), .A2(G134gat), .A3(new_n263_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1343gat));
  NOR2_X1   g661(.A1(new_n571_), .A2(new_n367_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n828_), .B2(new_n838_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n558_), .A3(new_n537_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n625_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT122), .B(G141gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n866_), .A2(new_n709_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n395_), .ZN(G1345gat));
  INV_X1    g670(.A(new_n866_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n308_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  OR3_X1    g674(.A1(new_n866_), .A2(G162gat), .A3(new_n263_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G162gat), .B1(new_n866_), .B2(new_n264_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1347gat));
  NAND2_X1  g677(.A1(new_n553_), .A2(new_n367_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n879_), .A2(new_n453_), .A3(new_n558_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n828_), .B2(new_n838_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n316_), .B1(new_n882_), .B2(new_n624_), .ZN(new_n883_));
  OR3_X1    g682(.A1(new_n883_), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n839_), .A2(new_n880_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n625_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n883_), .A2(KEYINPUT123), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT62), .B1(new_n883_), .B2(KEYINPUT123), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n884_), .B(new_n887_), .C1(new_n888_), .C2(new_n889_), .ZN(G1348gat));
  NOR2_X1   g689(.A1(new_n885_), .A2(new_n709_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n317_), .A2(KEYINPUT124), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n317_), .A2(KEYINPUT124), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n891_), .B2(new_n893_), .ZN(G1349gat));
  NOR2_X1   g694(.A1(new_n885_), .A2(new_n307_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n485_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n326_), .B2(new_n896_), .ZN(G1350gat));
  NOR2_X1   g697(.A1(new_n885_), .A2(new_n264_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n805_), .A2(new_n486_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT125), .ZN(new_n901_));
  OAI22_X1  g700(.A1(new_n899_), .A2(new_n336_), .B1(new_n885_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  OAI221_X1 g703(.A(KEYINPUT126), .B1(new_n885_), .B2(new_n901_), .C1(new_n899_), .C2(new_n336_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1351gat));
  NOR2_X1   g705(.A1(new_n558_), .A2(new_n537_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n839_), .A2(new_n863_), .A3(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT127), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n865_), .A2(KEYINPUT127), .A3(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G197gat), .B1(new_n912_), .B2(new_n624_), .ZN(new_n913_));
  AOI211_X1 g712(.A(new_n371_), .B(new_n625_), .C1(new_n910_), .C2(new_n911_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1352gat));
  INV_X1    g714(.A(new_n911_), .ZN(new_n916_));
  AOI21_X1  g715(.A(KEYINPUT127), .B1(new_n865_), .B2(new_n907_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n606_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(G204gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n912_), .A2(new_n373_), .A3(new_n606_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1353gat));
  OR2_X1    g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n912_), .B2(new_n308_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT63), .B(G211gat), .ZN(new_n924_));
  AOI211_X1 g723(.A(new_n307_), .B(new_n924_), .C1(new_n910_), .C2(new_n911_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1354gat));
  INV_X1    g725(.A(G218gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n912_), .A2(new_n927_), .A3(new_n805_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n264_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(G1355gat));
endmodule


