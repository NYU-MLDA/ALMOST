//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n981_, new_n982_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n991_,
    new_n992_, new_n994_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1004_, new_n1005_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  OR3_X1    g002(.A1(new_n203_), .A2(KEYINPUT77), .A3(KEYINPUT22), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT78), .B(G176gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT22), .B1(new_n203_), .B2(KEYINPUT77), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n208_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n209_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n202_), .B(new_n207_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT25), .B(G183gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(KEYINPUT24), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n202_), .ZN(new_n222_));
  INV_X1    g021(.A(G183gat), .ZN(new_n223_));
  INV_X1    g022(.A(G190gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT23), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n210_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .A4(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n216_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT80), .ZN(new_n229_));
  INV_X1    g028(.A(G204gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(G197gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT86), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(G197gat), .B2(new_n230_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n232_), .B1(new_n234_), .B2(new_n231_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT87), .ZN(new_n236_));
  AND2_X1   g035(.A1(G211gat), .A2(G218gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G211gat), .A2(G218gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G211gat), .ZN(new_n240_));
  INV_X1    g039(.A(G218gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G211gat), .A2(G218gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(KEYINPUT87), .A3(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n239_), .A2(new_n244_), .A3(KEYINPUT21), .ZN(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n230_), .A2(G197gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n239_), .A2(new_n244_), .B1(new_n249_), .B2(KEYINPUT21), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n232_), .B(new_n251_), .C1(new_n231_), .C2(new_n234_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n235_), .A2(new_n245_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n216_), .A2(new_n254_), .A3(new_n227_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n229_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT20), .ZN(new_n257_));
  INV_X1    g056(.A(new_n202_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT22), .B(G169gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n205_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT93), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n215_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n226_), .A2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(new_n260_), .B2(KEYINPUT93), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n219_), .A2(new_n222_), .A3(new_n221_), .ZN(new_n266_));
  OAI22_X1  g065(.A1(new_n262_), .A2(new_n265_), .B1(new_n214_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n245_), .A2(new_n235_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n250_), .A2(new_n252_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n257_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n256_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G226gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G8gat), .B(G36gat), .ZN(new_n278_));
  INV_X1    g077(.A(G92gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT18), .B(G64gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n255_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n254_), .B1(new_n216_), .B2(new_n227_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n270_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n266_), .A2(new_n214_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n205_), .A2(new_n259_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n202_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT93), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n289_), .A2(new_n290_), .B1(new_n263_), .B2(new_n226_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n287_), .B1(new_n291_), .B2(new_n261_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n257_), .B1(new_n292_), .B2(new_n253_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n286_), .A2(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n277_), .B(new_n283_), .C1(new_n276_), .C2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n253_), .B1(new_n229_), .B2(new_n255_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT20), .B1(new_n267_), .B2(new_n270_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n276_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n275_), .B1(new_n256_), .B2(new_n271_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n282_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT27), .B1(new_n295_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT96), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n302_), .B(new_n276_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n256_), .A2(new_n271_), .A3(new_n275_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n294_), .A2(new_n276_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT96), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n283_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n295_), .A2(KEYINPUT27), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT97), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT27), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n298_), .A2(new_n299_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n283_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n303_), .A2(new_n304_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n302_), .B1(new_n294_), .B2(new_n276_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n282_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT97), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n301_), .B1(new_n310_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n229_), .A2(new_n255_), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT30), .B(G15gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT31), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n320_), .B(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G227gat), .A2(G233gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n323_), .A2(new_n324_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G127gat), .B(G134gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(KEYINPUT81), .B(G43gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G71gat), .B(G99gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OR3_X1    g134(.A1(new_n326_), .A2(new_n327_), .A3(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n335_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n319_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(KEYINPUT95), .B(KEYINPUT0), .Z(new_n340_));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G57gat), .B(G85gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  INV_X1    g145(.A(G141gat), .ZN(new_n347_));
  INV_X1    g146(.A(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G155gat), .ZN(new_n350_));
  INV_X1    g149(.A(G162gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT1), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(G155gat), .B2(G162gat), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n350_), .A2(new_n351_), .A3(KEYINPUT1), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n346_), .B(new_n349_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(G141gat), .A3(G148gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n346_), .A2(KEYINPUT82), .A3(KEYINPUT2), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT3), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(G141gat), .B2(G148gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n359_), .A2(new_n363_), .A3(new_n364_), .A4(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G155gat), .B(G162gat), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n360_), .A2(new_n362_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n364_), .B1(new_n371_), .B2(new_n359_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n355_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n330_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n330_), .B(new_n355_), .C1(new_n370_), .C2(new_n372_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(KEYINPUT4), .A3(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n377_), .B(KEYINPUT94), .C1(KEYINPUT4), .C2(new_n375_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT94), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n375_), .A2(new_n379_), .A3(KEYINPUT4), .A4(new_n376_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n345_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n376_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n345_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n344_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n377_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT94), .B1(new_n375_), .B2(KEYINPUT4), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n380_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n383_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n384_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n344_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n385_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n396_));
  AOI211_X1 g195(.A(new_n396_), .B(new_n253_), .C1(new_n373_), .C2(KEYINPUT29), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n397_), .B2(KEYINPUT88), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n253_), .B1(new_n373_), .B2(KEYINPUT29), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT88), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n373_), .A2(KEYINPUT29), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(KEYINPUT85), .A3(new_n270_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT88), .ZN(new_n403_));
  INV_X1    g202(.A(new_n395_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n406_), .B(KEYINPUT89), .Z(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n398_), .A2(new_n400_), .A3(new_n405_), .A4(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT88), .B1(new_n399_), .B2(KEYINPUT85), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n411_), .A2(new_n404_), .B1(KEYINPUT88), .B2(new_n399_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n412_), .B2(new_n398_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n414_));
  OR3_X1    g213(.A1(new_n373_), .A2(KEYINPUT29), .A3(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G22gat), .B(G50gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n414_), .B1(new_n373_), .B2(KEYINPUT29), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n416_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n419_));
  OAI22_X1  g218(.A1(new_n410_), .A2(new_n413_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT90), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n418_), .A2(new_n419_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n405_), .A2(new_n400_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n411_), .A2(new_n404_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n407_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n423_), .B1(new_n426_), .B2(new_n409_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT90), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n409_), .A2(KEYINPUT91), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT91), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n412_), .A2(new_n430_), .A3(new_n398_), .A4(new_n408_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n406_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n429_), .A2(new_n423_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n422_), .A2(new_n428_), .A3(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n339_), .A2(new_n394_), .A3(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n427_), .B2(KEYINPUT90), .ZN(new_n436_));
  AOI211_X1 g235(.A(new_n421_), .B(new_n423_), .C1(new_n426_), .C2(new_n409_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n301_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n313_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n317_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n393_), .B(new_n439_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT98), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT98), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n434_), .A2(new_n319_), .A3(new_n444_), .A4(new_n393_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n295_), .A2(new_n300_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n344_), .B1(new_n382_), .B2(new_n345_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n388_), .B2(new_n345_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n392_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n392_), .A2(new_n450_), .ZN(new_n453_));
  OAI211_X1 g252(.A(KEYINPUT32), .B(new_n283_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT32), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n312_), .B1(new_n455_), .B2(new_n282_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  OAI22_X1  g256(.A1(new_n452_), .A2(new_n453_), .B1(new_n393_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n438_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n443_), .A2(new_n445_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n338_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n435_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G169gat), .B(G197gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT76), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G113gat), .B(G141gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT75), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT74), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT69), .B(G43gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G29gat), .ZN(new_n472_));
  INV_X1    g271(.A(G36gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G29gat), .A2(G36gat), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n474_), .A2(G50gat), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(G50gat), .B1(new_n474_), .B2(new_n475_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n471_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n475_), .ZN(new_n479_));
  INV_X1    g278(.A(G50gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n474_), .A2(G50gat), .A3(new_n475_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n470_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G1gat), .ZN(new_n485_));
  AND2_X1   g284(.A1(KEYINPUT72), .A2(G8gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(KEYINPUT72), .A2(G8gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n485_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(KEYINPUT14), .A2(G1gat), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(G8gat), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(new_n489_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G1gat), .ZN(new_n495_));
  INV_X1    g294(.A(G8gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n491_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  AOI211_X1 g297(.A(new_n469_), .B(new_n484_), .C1(new_n493_), .C2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n493_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n484_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT74), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n498_), .A2(new_n484_), .A3(new_n493_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT73), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n468_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n500_), .A2(new_n501_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n469_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n500_), .A2(KEYINPUT74), .A3(new_n501_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT73), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n504_), .B(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n512_), .A3(KEYINPUT75), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n467_), .B1(new_n506_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT15), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n484_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n478_), .A2(new_n483_), .A3(KEYINPUT15), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n500_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n512_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n521_), .A2(new_n467_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n466_), .B1(new_n514_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n467_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n510_), .A2(new_n512_), .A3(KEYINPUT75), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT75), .B1(new_n510_), .B2(new_n512_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n521_), .A2(new_n467_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n466_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n523_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G230gat), .A2(G233gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(G71gat), .B(G78gat), .Z(new_n533_));
  INV_X1    g332(.A(G57gat), .ZN(new_n534_));
  INV_X1    g333(.A(G64gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT11), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G57gat), .A2(G64gat), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT65), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n538_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(KEYINPUT11), .ZN(new_n543_));
  AND2_X1   g342(.A1(G57gat), .A2(G64gat), .ZN(new_n544_));
  NOR2_X1   g343(.A1(G57gat), .A2(G64gat), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n541_), .B(KEYINPUT11), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n540_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT11), .B1(new_n544_), .B2(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT65), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n550_), .A2(new_n539_), .A3(new_n533_), .A4(new_n546_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n548_), .A2(KEYINPUT66), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT66), .B1(new_n548_), .B2(new_n551_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G85gat), .B(G92gat), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT9), .ZN(new_n557_));
  INV_X1    g356(.A(G85gat), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n558_), .A2(new_n279_), .A3(KEYINPUT9), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G99gat), .A2(G106gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT6), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT6), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(G99gat), .A3(G106gat), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n559_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT10), .B(G99gat), .Z(new_n565_));
  INV_X1    g364(.A(G106gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n557_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT8), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n561_), .A2(new_n563_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT64), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT7), .ZN(new_n573_));
  INV_X1    g372(.A(G99gat), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n566_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n561_), .A2(new_n563_), .A3(KEYINPUT64), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n572_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n569_), .B1(new_n580_), .B2(new_n556_), .ZN(new_n581_));
  AOI211_X1 g380(.A(KEYINPUT8), .B(new_n555_), .C1(new_n578_), .C2(new_n570_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n568_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n554_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n578_), .A2(new_n570_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n569_), .A3(new_n556_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT64), .B1(new_n561_), .B2(new_n563_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(new_n577_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n555_), .B1(new_n588_), .B2(new_n579_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n586_), .B1(new_n589_), .B2(new_n569_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n590_), .B(new_n568_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n532_), .B1(new_n584_), .B2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT67), .B(KEYINPUT12), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT66), .ZN(new_n595_));
  INV_X1    g394(.A(new_n551_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n550_), .A2(new_n546_), .B1(new_n539_), .B2(new_n533_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n548_), .A2(KEYINPUT66), .A3(new_n551_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n568_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n561_), .A2(new_n563_), .A3(KEYINPUT64), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n602_), .A2(new_n587_), .A3(new_n577_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT8), .B1(new_n603_), .B2(new_n555_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n601_), .B1(new_n604_), .B2(new_n586_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n594_), .B1(new_n600_), .B2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n596_), .A2(new_n597_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n583_), .A2(KEYINPUT12), .A3(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n606_), .A2(new_n532_), .A3(new_n591_), .A4(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT68), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n608_), .A2(new_n591_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n612_), .A2(KEYINPUT68), .A3(new_n532_), .A4(new_n606_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n592_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(new_n230_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT5), .B(G176gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  NOR2_X1   g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  AOI211_X1 g419(.A(new_n592_), .B(new_n620_), .C1(new_n611_), .C2(new_n613_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n622_), .A2(KEYINPUT13), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(KEYINPUT13), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n462_), .A2(new_n531_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n500_), .B(new_n627_), .Z(new_n628_));
  OR2_X1    g427(.A1(new_n628_), .A2(new_n607_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(new_n240_), .ZN(new_n631_));
  XOR2_X1   g430(.A(KEYINPUT16), .B(G183gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(KEYINPUT17), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n607_), .B2(new_n628_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n628_), .B(new_n600_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n633_), .B(KEYINPUT17), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT35), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n519_), .A2(new_n583_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n484_), .B(new_n568_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT34), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n641_), .A2(KEYINPUT70), .A3(new_n644_), .A4(new_n642_), .ZN(new_n645_));
  OAI211_X1 g444(.A(KEYINPUT70), .B(new_n642_), .C1(new_n605_), .C2(new_n518_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT34), .ZN(new_n647_));
  INV_X1    g446(.A(G232gat), .ZN(new_n648_));
  INV_X1    g447(.A(G233gat), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n645_), .A2(new_n647_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n640_), .B(new_n643_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n645_), .A2(new_n647_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n650_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(KEYINPUT35), .A3(new_n652_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(G190gat), .B(G218gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(G134gat), .B(G162gat), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n660_), .B(new_n661_), .Z(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT36), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT36), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n655_), .A2(new_n665_), .A3(new_n658_), .A4(new_n662_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n664_), .A2(KEYINPUT37), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n666_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n663_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n659_), .B2(KEYINPUT71), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT71), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n655_), .A2(new_n671_), .A3(new_n658_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n668_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n639_), .B(new_n667_), .C1(new_n673_), .C2(KEYINPUT37), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n626_), .A2(new_n675_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n676_), .A2(G1gat), .A3(new_n393_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT38), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT38), .ZN(new_n679_));
  INV_X1    g478(.A(new_n639_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n673_), .A2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n626_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n485_), .B1(new_n682_), .B2(new_n394_), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n678_), .A2(new_n679_), .A3(new_n683_), .ZN(G1324gat));
  INV_X1    g483(.A(new_n676_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n319_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n685_), .B(new_n686_), .C1(new_n487_), .C2(new_n486_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n682_), .A2(new_n686_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G8gat), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(KEYINPUT39), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(KEYINPUT39), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n692_), .B(new_n694_), .ZN(G1325gat));
  INV_X1    g494(.A(G15gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n682_), .B2(new_n338_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(KEYINPUT41), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(KEYINPUT41), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n685_), .A2(new_n696_), .A3(new_n338_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n699_), .A2(new_n700_), .A3(new_n701_), .ZN(G1326gat));
  INV_X1    g501(.A(G22gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n682_), .B2(new_n434_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT42), .Z(new_n705_));
  NAND3_X1  g504(.A1(new_n685_), .A2(new_n703_), .A3(new_n434_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1327gat));
  NOR3_X1   g506(.A1(new_n653_), .A2(new_n654_), .A3(new_n640_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n643_), .A2(new_n640_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n657_), .B2(new_n652_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT71), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n672_), .A3(new_n663_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n666_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(new_n639_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n626_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT103), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n626_), .A2(new_n717_), .A3(new_n714_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n472_), .A3(new_n394_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT37), .B1(new_n712_), .B2(new_n666_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n667_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n434_), .A2(new_n319_), .A3(new_n393_), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n726_), .A2(KEYINPUT98), .B1(new_n438_), .B2(new_n458_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n338_), .B1(new_n727_), .B2(new_n445_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n721_), .B(new_n725_), .C1(new_n728_), .C2(new_n435_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n462_), .B2(new_n724_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n625_), .A2(new_n531_), .A3(new_n639_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(KEYINPUT100), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT100), .ZN(new_n736_));
  INV_X1    g535(.A(new_n732_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n738_), .B2(KEYINPUT44), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n735_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n460_), .A2(new_n461_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n435_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n721_), .B1(new_n743_), .B2(new_n725_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n462_), .A2(KEYINPUT43), .A3(new_n724_), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT44), .B(new_n732_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT101), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT101), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n738_), .A2(new_n748_), .A3(KEYINPUT44), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n740_), .A2(new_n750_), .A3(new_n394_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT102), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G29gat), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n751_), .A2(new_n752_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n720_), .B1(new_n754_), .B2(new_n755_), .ZN(G1328gat));
  INV_X1    g555(.A(KEYINPUT46), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n739_), .A2(new_n735_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n473_), .B1(new_n758_), .B2(new_n686_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n716_), .A2(new_n473_), .A3(new_n686_), .A4(new_n718_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n757_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n740_), .A2(new_n750_), .A3(new_n686_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G36gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n760_), .B(KEYINPUT45), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(KEYINPUT46), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n763_), .A2(new_n767_), .ZN(G1329gat));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n740_), .A2(new_n750_), .A3(new_n338_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(G43gat), .ZN(new_n771_));
  INV_X1    g570(.A(G43gat), .ZN(new_n772_));
  AND4_X1   g571(.A1(new_n772_), .A2(new_n716_), .A3(new_n338_), .A4(new_n718_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n769_), .B1(new_n771_), .B2(new_n774_), .ZN(new_n775_));
  AOI211_X1 g574(.A(KEYINPUT47), .B(new_n773_), .C1(new_n770_), .C2(G43gat), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1330gat));
  NAND3_X1  g576(.A1(new_n719_), .A2(new_n480_), .A3(new_n434_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n758_), .A2(new_n434_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n480_), .ZN(G1331gat));
  INV_X1    g579(.A(new_n625_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n531_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n743_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n681_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(G57gat), .A3(new_n394_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n784_), .A2(new_n674_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n534_), .B1(new_n790_), .B2(new_n393_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT104), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n792_), .B2(new_n791_), .ZN(G1332gat));
  AOI21_X1  g593(.A(new_n535_), .B1(new_n787_), .B2(new_n686_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT105), .B(KEYINPUT48), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n796_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n789_), .A2(new_n535_), .A3(new_n686_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n797_), .A2(new_n798_), .A3(new_n799_), .ZN(G1333gat));
  INV_X1    g599(.A(G71gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n787_), .B2(new_n338_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT106), .B(KEYINPUT49), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n803_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n789_), .A2(new_n801_), .A3(new_n338_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(G1334gat));
  INV_X1    g606(.A(G78gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n787_), .B2(new_n434_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n810_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n789_), .A2(new_n808_), .A3(new_n434_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(G1335gat));
  NAND3_X1  g613(.A1(new_n731_), .A2(new_n680_), .A3(new_n783_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n815_), .A2(new_n558_), .A3(new_n393_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n785_), .A2(new_n714_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G85gat), .B1(new_n818_), .B2(new_n394_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n816_), .A2(new_n819_), .ZN(G1336gat));
  NOR3_X1   g619(.A1(new_n815_), .A2(new_n279_), .A3(new_n319_), .ZN(new_n821_));
  AOI21_X1  g620(.A(G92gat), .B1(new_n818_), .B2(new_n686_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n815_), .B2(new_n461_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n338_), .A2(new_n565_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n817_), .B2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g626(.A1(new_n818_), .A2(new_n566_), .A3(new_n434_), .ZN(new_n828_));
  OAI21_X1  g627(.A(G106gat), .B1(new_n815_), .B2(new_n438_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n829_), .A2(KEYINPUT52), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(KEYINPUT52), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n828_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT53), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n828_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1339gat));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n467_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n529_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n530_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n837_), .B1(new_n622_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT55), .B1(new_n611_), .B2(new_n613_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n608_), .A2(new_n591_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n593_), .B1(new_n554_), .B2(new_n583_), .ZN(new_n845_));
  OAI211_X1 g644(.A(G230gat), .B(G233gat), .C1(new_n844_), .C2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n609_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n620_), .B1(new_n843_), .B2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(KEYINPUT108), .A2(KEYINPUT56), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n523_), .A2(new_n530_), .B1(new_n614_), .B2(new_n618_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n620_), .B(new_n850_), .C1(new_n843_), .C2(new_n848_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n514_), .A2(new_n522_), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n856_), .A2(new_n529_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(KEYINPUT109), .C1(new_n619_), .C2(new_n621_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n842_), .A2(new_n855_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n713_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT110), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(KEYINPUT57), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864_));
  INV_X1    g663(.A(new_n621_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n857_), .B(new_n865_), .C1(KEYINPUT56), .C2(new_n849_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n849_), .A2(KEYINPUT56), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n849_), .A2(KEYINPUT56), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n841_), .A2(new_n621_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n870_), .A2(KEYINPUT58), .A3(new_n867_), .A4(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n869_), .B(new_n872_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n859_), .B(new_n713_), .C1(new_n861_), .C2(KEYINPUT57), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n863_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n680_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT112), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n623_), .A2(new_n531_), .A3(new_n624_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT54), .B1(new_n674_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n878_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n724_), .A2(new_n880_), .A3(new_n881_), .A4(new_n639_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n875_), .A2(new_n884_), .A3(new_n680_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n877_), .A2(new_n883_), .A3(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n339_), .A2(new_n434_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n394_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(KEYINPUT59), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(G113gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n531_), .A2(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT113), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n888_), .B1(new_n876_), .B2(new_n883_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT111), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n895_), .A2(new_n896_), .A3(KEYINPUT59), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n895_), .B2(KEYINPUT59), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n890_), .B(new_n893_), .C1(new_n898_), .C2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n891_), .B1(new_n895_), .B2(new_n531_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT114), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n900_), .A2(KEYINPUT114), .A3(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1340gat));
  OAI21_X1  g705(.A(new_n890_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G120gat), .B1(new_n907_), .B2(new_n781_), .ZN(new_n908_));
  INV_X1    g707(.A(G120gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n781_), .B2(KEYINPUT60), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n910_), .B1(KEYINPUT60), .B2(new_n909_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n908_), .B1(new_n895_), .B2(new_n911_), .ZN(G1341gat));
  AOI21_X1  g711(.A(G127gat), .B1(new_n894_), .B2(new_n639_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT115), .ZN(new_n914_));
  INV_X1    g713(.A(new_n907_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n639_), .A2(G127gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(G1342gat));
  AOI21_X1  g716(.A(G134gat), .B1(new_n894_), .B2(new_n673_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT116), .Z(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT117), .B(G134gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n725_), .A2(new_n920_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT118), .Z(new_n922_));
  AOI21_X1  g721(.A(new_n919_), .B1(new_n915_), .B2(new_n922_), .ZN(G1343gat));
  NAND2_X1  g722(.A1(new_n876_), .A2(new_n883_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n438_), .A2(new_n338_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n319_), .A2(new_n394_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n924_), .A2(new_n925_), .A3(new_n927_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(KEYINPUT119), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n782_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n625_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g732(.A1(new_n929_), .A2(new_n639_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(KEYINPUT120), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n929_), .A2(new_n936_), .A3(new_n639_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT61), .B(G155gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n935_), .A2(new_n937_), .A3(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n938_), .ZN(new_n940_));
  OR2_X1    g739(.A1(new_n928_), .A2(KEYINPUT119), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n928_), .A2(KEYINPUT119), .ZN(new_n942_));
  AOI211_X1 g741(.A(KEYINPUT120), .B(new_n680_), .C1(new_n941_), .C2(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n936_), .B1(new_n929_), .B2(new_n639_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n940_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n939_), .A2(new_n945_), .ZN(G1346gat));
  NOR2_X1   g745(.A1(new_n713_), .A2(G162gat), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n929_), .A2(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n724_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(new_n351_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(KEYINPUT121), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n948_), .B(new_n952_), .C1(new_n351_), .C2(new_n949_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1347gat));
  NOR2_X1   g753(.A1(new_n319_), .A2(new_n394_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n338_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n956_), .A2(new_n531_), .ZN(new_n957_));
  XOR2_X1   g756(.A(new_n957_), .B(KEYINPUT122), .Z(new_n958_));
  NOR2_X1   g757(.A1(new_n958_), .A2(new_n434_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n203_), .B1(new_n886_), .B2(new_n959_), .ZN(new_n960_));
  XOR2_X1   g759(.A(new_n960_), .B(KEYINPUT62), .Z(new_n961_));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n956_), .A2(new_n434_), .ZN(new_n963_));
  AND3_X1   g762(.A1(new_n886_), .A2(new_n962_), .A3(new_n963_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n962_), .B1(new_n886_), .B2(new_n963_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n966_), .A2(new_n782_), .A3(new_n259_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n961_), .A2(new_n967_), .ZN(G1348gat));
  AND2_X1   g767(.A1(new_n924_), .A2(new_n963_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n969_), .A2(G176gat), .A3(new_n625_), .ZN(new_n970_));
  XOR2_X1   g769(.A(new_n970_), .B(KEYINPUT125), .Z(new_n971_));
  NAND2_X1  g770(.A1(new_n886_), .A2(new_n963_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(KEYINPUT123), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n886_), .A2(new_n962_), .A3(new_n963_), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n973_), .A2(new_n625_), .A3(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(new_n205_), .ZN(new_n976_));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n975_), .A2(KEYINPUT124), .A3(new_n205_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n971_), .B1(new_n978_), .B2(new_n979_), .ZN(G1349gat));
  AOI21_X1  g779(.A(G183gat), .B1(new_n969_), .B2(new_n639_), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n680_), .A2(new_n217_), .ZN(new_n982_));
  AOI21_X1  g781(.A(new_n981_), .B1(new_n966_), .B2(new_n982_), .ZN(G1350gat));
  NAND4_X1  g782(.A1(new_n973_), .A2(new_n218_), .A3(new_n673_), .A4(new_n974_), .ZN(new_n984_));
  NOR3_X1   g783(.A1(new_n964_), .A2(new_n965_), .A3(new_n724_), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n984_), .B1(new_n985_), .B2(new_n224_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n986_), .A2(KEYINPUT126), .ZN(new_n987_));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n988_));
  OAI211_X1 g787(.A(new_n984_), .B(new_n988_), .C1(new_n985_), .C2(new_n224_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n987_), .A2(new_n989_), .ZN(G1351gat));
  AND3_X1   g789(.A1(new_n924_), .A2(new_n925_), .A3(new_n955_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n991_), .A2(new_n782_), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n992_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g792(.A1(new_n991_), .A2(new_n625_), .ZN(new_n994_));
  XNOR2_X1  g793(.A(new_n994_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g794(.A1(new_n991_), .A2(new_n639_), .ZN(new_n996_));
  XNOR2_X1  g795(.A(KEYINPUT63), .B(G211gat), .ZN(new_n997_));
  NOR2_X1   g796(.A1(new_n996_), .A2(new_n997_), .ZN(new_n998_));
  INV_X1    g797(.A(KEYINPUT63), .ZN(new_n999_));
  NAND3_X1  g798(.A1(new_n996_), .A2(new_n999_), .A3(new_n240_), .ZN(new_n1000_));
  OR2_X1    g799(.A1(new_n1000_), .A2(KEYINPUT127), .ZN(new_n1001_));
  NAND2_X1  g800(.A1(new_n1000_), .A2(KEYINPUT127), .ZN(new_n1002_));
  AOI21_X1  g801(.A(new_n998_), .B1(new_n1001_), .B2(new_n1002_), .ZN(G1354gat));
  AOI21_X1  g802(.A(G218gat), .B1(new_n991_), .B2(new_n673_), .ZN(new_n1004_));
  NOR2_X1   g803(.A1(new_n724_), .A2(new_n241_), .ZN(new_n1005_));
  AOI21_X1  g804(.A(new_n1004_), .B1(new_n991_), .B2(new_n1005_), .ZN(G1355gat));
endmodule


