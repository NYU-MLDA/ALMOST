//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n874_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT69), .ZN(new_n203_));
  XOR2_X1   g002(.A(G134gat), .B(G162gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT36), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G232gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT34), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT7), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G85gat), .B(G92gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n210_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n212_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n211_), .B(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n215_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n218_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(KEYINPUT65), .A3(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n219_), .A2(KEYINPUT8), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT9), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G85gat), .A3(G92gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT10), .B(G99gat), .ZN(new_n228_));
  OAI221_X1 g027(.A(new_n227_), .B1(new_n218_), .B2(new_n226_), .C1(G106gat), .C2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(new_n213_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT65), .B1(new_n222_), .B2(new_n223_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G29gat), .B(G36gat), .Z(new_n234_));
  XOR2_X1   g033(.A(G43gat), .B(G50gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n225_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(KEYINPUT15), .Z(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(new_n225_), .B2(new_n233_), .ZN(new_n239_));
  OAI211_X1 g038(.A(KEYINPUT35), .B(new_n209_), .C1(new_n237_), .C2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n225_), .A2(new_n233_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n238_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n209_), .A2(KEYINPUT35), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n209_), .A2(KEYINPUT35), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n225_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .A4(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n240_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n207_), .B1(new_n248_), .B2(KEYINPUT70), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n250_));
  INV_X1    g049(.A(new_n207_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n240_), .A2(new_n247_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n205_), .A2(new_n206_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT37), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n249_), .A2(new_n252_), .B1(new_n248_), .B2(new_n254_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n257_), .A2(KEYINPUT37), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(KEYINPUT37), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G57gat), .B(G64gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT66), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n266_), .A2(KEYINPUT11), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(KEYINPUT11), .ZN(new_n268_));
  XOR2_X1   g067(.A(G71gat), .B(G78gat), .Z(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n268_), .A2(new_n269_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G15gat), .B(G22gat), .ZN(new_n273_));
  INV_X1    g072(.A(G1gat), .ZN(new_n274_));
  INV_X1    g073(.A(G8gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT14), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G1gat), .B(G8gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n272_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G231gat), .A2(G233gat), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G127gat), .B(G155gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G183gat), .B(G211gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT17), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT17), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n283_), .A2(new_n294_), .A3(new_n284_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n264_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT73), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(G127gat), .B(G134gat), .Z(new_n301_));
  XOR2_X1   g100(.A(G113gat), .B(G120gat), .Z(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  INV_X1    g102(.A(G155gat), .ZN(new_n304_));
  INV_X1    g103(.A(G162gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(KEYINPUT79), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT79), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(G155gat), .B2(G162gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT81), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n311_), .B1(new_n313_), .B2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n310_), .A2(KEYINPUT1), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n306_), .A2(new_n308_), .B1(KEYINPUT1), .B2(new_n310_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(KEYINPUT80), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n310_), .A2(KEYINPUT1), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n309_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT80), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G141gat), .B(G148gat), .Z(new_n328_));
  AOI21_X1  g127(.A(new_n319_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n303_), .B1(new_n329_), .B2(KEYINPUT90), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n307_), .A2(G155gat), .A3(G162gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT79), .B1(new_n304_), .B2(new_n305_), .ZN(new_n332_));
  OAI211_X1 g131(.A(KEYINPUT80), .B(new_n323_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n320_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n321_), .A2(KEYINPUT80), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n328_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n318_), .A2(new_n313_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n337_), .A2(new_n339_), .A3(new_n303_), .A4(KEYINPUT90), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n300_), .B1(new_n330_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G85gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT0), .B(G57gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n337_), .A2(KEYINPUT90), .A3(new_n339_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n303_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n347_), .B1(new_n350_), .B2(new_n340_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n300_), .B(KEYINPUT91), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n303_), .A2(new_n347_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n352_), .B1(new_n329_), .B2(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n342_), .B(new_n346_), .C1(new_n351_), .C2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT95), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n342_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n346_), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n355_), .A2(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n357_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G78gat), .B(G106gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(KEYINPUT21), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT21), .ZN(new_n368_));
  INV_X1    g167(.A(new_n366_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n364_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G211gat), .B(G218gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n369_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n371_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT83), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n367_), .A2(new_n371_), .A3(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n372_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n329_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G228gat), .ZN(new_n381_));
  INV_X1    g180(.A(G233gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n337_), .A2(new_n339_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT29), .ZN(new_n386_));
  INV_X1    g185(.A(new_n383_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n378_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n363_), .B1(new_n384_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI211_X1 g190(.A(KEYINPUT85), .B(new_n363_), .C1(new_n384_), .C2(new_n388_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n384_), .A2(new_n388_), .A3(new_n363_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT86), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n384_), .A2(new_n388_), .A3(KEYINPUT86), .A4(new_n363_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT28), .B1(new_n385_), .B2(KEYINPUT29), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT28), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n329_), .A2(new_n401_), .A3(new_n379_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n399_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(G22gat), .B(G50gat), .Z(new_n405_));
  NAND3_X1  g204(.A1(new_n400_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n405_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n406_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n403_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n393_), .A2(new_n398_), .A3(new_n407_), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n394_), .A2(KEYINPUT84), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n380_), .A2(new_n383_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n387_), .B1(new_n386_), .B2(new_n378_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n362_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n389_), .A2(KEYINPUT84), .A3(new_n394_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n410_), .A2(new_n407_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n411_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT24), .ZN(new_n422_));
  INV_X1    g221(.A(G169gat), .ZN(new_n423_));
  INV_X1    g222(.A(G176gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G183gat), .A2(G190gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT23), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(G190gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT26), .B1(new_n431_), .B2(KEYINPUT75), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT75), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT26), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(G190gat), .ZN(new_n435_));
  INV_X1    g234(.A(G183gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT25), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT25), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G183gat), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n432_), .A2(new_n435_), .A3(new_n437_), .A4(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n423_), .A2(new_n424_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G169gat), .A2(G176gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(KEYINPUT24), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n430_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(G169gat), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n428_), .B(new_n429_), .C1(G183gat), .C2(G190gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT76), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n444_), .A2(KEYINPUT76), .A3(new_n448_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G15gat), .B(G43gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G71gat), .B(G99gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n456_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT78), .B(KEYINPUT31), .Z(new_n460_));
  OR2_X1    g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n460_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464_));
  XOR2_X1   g263(.A(new_n464_), .B(KEYINPUT77), .Z(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT30), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(new_n303_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n461_), .A2(new_n467_), .A3(new_n462_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n359_), .A2(new_n360_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n376_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT83), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n373_), .A2(new_n374_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n474_), .A2(new_n475_), .B1(new_n476_), .B2(new_n370_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n451_), .A2(new_n477_), .A3(new_n452_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n425_), .A2(new_n428_), .A3(KEYINPUT88), .A4(new_n429_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT25), .B(G183gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT26), .B(G190gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n482_), .A2(new_n443_), .A3(new_n483_), .A4(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n448_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n479_), .B1(new_n488_), .B2(new_n378_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n478_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G226gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G8gat), .B(G36gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G64gat), .B(G92gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n487_), .A2(new_n448_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n479_), .B1(new_n500_), .B2(new_n477_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n493_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n452_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT76), .B1(new_n444_), .B2(new_n448_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n378_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n494_), .A2(new_n499_), .A3(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n507_), .A2(KEYINPUT27), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n477_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT20), .B1(new_n488_), .B2(new_n378_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n493_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n478_), .A2(new_n489_), .A3(new_n502_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n499_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n508_), .A2(new_n515_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n509_), .A2(new_n510_), .A3(new_n493_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n502_), .B1(new_n478_), .B2(new_n489_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n514_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n499_), .B1(new_n494_), .B2(new_n506_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n516_), .B1(KEYINPUT27), .B2(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n421_), .A2(new_n473_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n361_), .B1(new_n411_), .B2(new_n420_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n522_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT92), .B(KEYINPUT33), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n342_), .A2(new_n346_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n350_), .A2(new_n340_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n354_), .B1(new_n529_), .B2(KEYINPUT4), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n527_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT4), .B1(new_n330_), .B2(new_n341_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n354_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n358_), .B1(new_n529_), .B2(new_n300_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT33), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n352_), .B1(new_n330_), .B2(new_n341_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n300_), .B1(new_n329_), .B2(new_n353_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n537_), .B(new_n358_), .C1(new_n351_), .C2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n521_), .A2(new_n531_), .A3(new_n536_), .A4(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT93), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n514_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n539_), .A2(new_n507_), .A3(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n544_), .A2(KEYINPUT93), .A3(new_n531_), .A4(new_n536_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n494_), .A2(KEYINPUT94), .A3(new_n506_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n499_), .A2(KEYINPUT32), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT94), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n511_), .A2(new_n512_), .A3(new_n547_), .ZN(new_n549_));
  OAI22_X1  g348(.A1(new_n546_), .A2(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(new_n545_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n415_), .A2(KEYINPUT85), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n389_), .A2(new_n390_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(new_n419_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n416_), .A2(new_n417_), .B1(new_n410_), .B2(new_n407_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n525_), .A2(new_n526_), .B1(new_n552_), .B2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n524_), .B1(new_n559_), .B2(new_n471_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n279_), .A2(new_n236_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT74), .ZN(new_n566_));
  INV_X1    g365(.A(new_n236_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(new_n280_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n566_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n242_), .A2(new_n280_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n569_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n564_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n571_), .A2(new_n575_), .A3(new_n564_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G120gat), .B(G148gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n272_), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n241_), .A2(KEYINPUT67), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n241_), .A2(new_n587_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n225_), .A2(new_n272_), .A3(new_n233_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(KEYINPUT67), .A3(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n588_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(KEYINPUT12), .A3(new_n590_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT12), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n241_), .A2(new_n595_), .A3(new_n587_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n592_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n586_), .B1(new_n593_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n593_), .A2(new_n597_), .A3(new_n586_), .ZN(new_n600_));
  OR3_X1    g399(.A1(new_n599_), .A2(KEYINPUT13), .A3(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT13), .B1(new_n599_), .B2(new_n600_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n580_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n560_), .A2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n299_), .A2(new_n274_), .A3(new_n361_), .A4(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT38), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT97), .Z(new_n608_));
  NAND2_X1  g407(.A1(new_n552_), .A2(new_n558_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n421_), .A2(new_n472_), .A3(new_n526_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n471_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n523_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n256_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n614_), .A2(new_n297_), .A3(new_n603_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n274_), .B1(new_n615_), .B2(new_n361_), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n605_), .A2(KEYINPUT96), .A3(new_n606_), .ZN(new_n617_));
  OAI21_X1  g416(.A(KEYINPUT96), .B1(new_n605_), .B2(new_n606_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n616_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n608_), .A2(new_n619_), .ZN(G1324gat));
  NAND2_X1  g419(.A1(new_n299_), .A2(new_n604_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n621_), .A2(G8gat), .A3(new_n526_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT98), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n275_), .B1(new_n615_), .B2(new_n522_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT39), .Z(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n623_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  NAND2_X1  g428(.A1(new_n615_), .A2(new_n471_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G15gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT100), .Z(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(KEYINPUT41), .ZN(new_n633_));
  OR3_X1    g432(.A1(new_n621_), .A2(G15gat), .A3(new_n612_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(KEYINPUT41), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(G1326gat));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n615_), .B2(new_n421_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT42), .Z(new_n639_));
  NOR2_X1   g438(.A1(new_n558_), .A2(G22gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT101), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n639_), .B1(new_n621_), .B2(new_n641_), .ZN(G1327gat));
  NOR2_X1   g441(.A1(new_n297_), .A2(new_n259_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n604_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(G29gat), .B1(new_n644_), .B2(new_n361_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n471_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n646_), .B(new_n263_), .C1(new_n647_), .C2(new_n523_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT102), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n560_), .A2(new_n650_), .A3(new_n646_), .A4(new_n263_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT43), .B1(new_n613_), .B2(new_n264_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n649_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n603_), .A2(new_n296_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT44), .B1(new_n653_), .B2(new_n654_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n361_), .A2(G29gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n645_), .B1(new_n657_), .B2(new_n658_), .ZN(G1328gat));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n655_), .A2(new_n656_), .A3(new_n526_), .ZN(new_n665_));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n656_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n654_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n522_), .A3(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(KEYINPUT103), .A3(G36gat), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n667_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n526_), .A2(G36gat), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n560_), .A2(new_n603_), .A3(new_n643_), .A4(new_n673_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT104), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT104), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT45), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n679_), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n660_), .A2(new_n661_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n663_), .B1(new_n672_), .B2(new_n684_), .ZN(new_n685_));
  AOI211_X1 g484(.A(new_n662_), .B(new_n683_), .C1(new_n667_), .C2(new_n671_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1329gat));
  AOI21_X1  g486(.A(G43gat), .B1(new_n644_), .B2(new_n471_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n471_), .A2(G43gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n657_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g490(.A(G50gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n644_), .A2(new_n692_), .A3(new_n421_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n657_), .A2(new_n421_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(KEYINPUT106), .ZN(new_n695_));
  OAI21_X1  g494(.A(G50gat), .B1(new_n694_), .B2(KEYINPUT106), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n695_), .B2(new_n696_), .ZN(G1331gat));
  NAND2_X1  g496(.A1(new_n601_), .A2(new_n602_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n299_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n613_), .A2(new_n579_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT107), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n472_), .B1(new_n703_), .B2(KEYINPUT108), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(KEYINPUT108), .B2(new_n703_), .ZN(new_n705_));
  INV_X1    g504(.A(G57gat), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n577_), .A2(new_n292_), .A3(new_n295_), .A4(new_n578_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n698_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n614_), .A2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n472_), .A2(KEYINPUT109), .ZN(new_n710_));
  MUX2_X1   g509(.A(KEYINPUT109), .B(new_n710_), .S(G57gat), .Z(new_n711_));
  AOI22_X1  g510(.A1(new_n705_), .A2(new_n706_), .B1(new_n709_), .B2(new_n711_), .ZN(G1332gat));
  INV_X1    g511(.A(G64gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n709_), .B2(new_n522_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT48), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n522_), .A2(new_n713_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n703_), .B2(new_n716_), .ZN(G1333gat));
  INV_X1    g516(.A(G71gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n709_), .B2(new_n471_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT110), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n720_), .A2(KEYINPUT49), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(KEYINPUT49), .ZN(new_n722_));
  INV_X1    g521(.A(new_n703_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n718_), .A3(new_n471_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n721_), .A2(new_n722_), .A3(new_n724_), .ZN(G1334gat));
  NAND2_X1  g524(.A1(new_n709_), .A2(new_n421_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G78gat), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT50), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n558_), .A2(G78gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT111), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n728_), .B1(new_n703_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT112), .ZN(G1335gat));
  AND4_X1   g531(.A1(new_n256_), .A2(new_n702_), .A3(new_n296_), .A4(new_n699_), .ZN(new_n733_));
  INV_X1    g532(.A(G85gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n361_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n698_), .A2(new_n297_), .A3(new_n579_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n653_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737_), .B2(new_n472_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1336gat));
  INV_X1    g538(.A(G92gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n733_), .A2(new_n740_), .A3(new_n522_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G92gat), .B1(new_n737_), .B2(new_n526_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  INV_X1    g542(.A(new_n228_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n733_), .A2(new_n744_), .A3(new_n471_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n653_), .A2(new_n471_), .A3(new_n736_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(G99gat), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n746_), .A3(G99gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g550(.A(G106gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n733_), .A2(new_n752_), .A3(new_n421_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n653_), .A2(new_n421_), .A3(new_n736_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(G106gat), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n754_), .A3(G106gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XOR2_X1   g557(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(G1339gat));
  XNOR2_X1  g559(.A(new_n707_), .B(KEYINPUT115), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n698_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT54), .B1(new_n762_), .B2(new_n263_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n264_), .A2(new_n698_), .A3(new_n764_), .A4(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n564_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n574_), .A2(new_n569_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OR3_X1    g570(.A1(new_n771_), .A2(new_n576_), .A3(KEYINPUT118), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT118), .B1(new_n771_), .B2(new_n576_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n600_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n772_), .A2(new_n773_), .B1(new_n774_), .B2(new_n598_), .ZN(new_n775_));
  OR3_X1    g574(.A1(new_n597_), .A2(KEYINPUT116), .A3(KEYINPUT55), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n594_), .A2(new_n592_), .A3(new_n596_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT55), .B1(new_n597_), .B2(KEYINPUT116), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n586_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT56), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n774_), .A2(new_n579_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n779_), .B2(new_n586_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n786_), .B2(new_n781_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n775_), .B1(new_n783_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n768_), .B1(new_n788_), .B2(new_n256_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n775_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n780_), .A2(new_n781_), .A3(KEYINPUT56), .ZN(new_n791_));
  INV_X1    g590(.A(new_n784_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n790_), .B1(new_n793_), .B2(new_n782_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT57), .A3(new_n259_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n600_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n779_), .A2(new_n785_), .A3(new_n586_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n796_), .B1(new_n799_), .B2(new_n786_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n786_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n801_), .A2(KEYINPUT58), .A3(new_n798_), .A4(new_n797_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n802_), .A3(new_n263_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n789_), .A2(new_n795_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n767_), .B1(new_n804_), .B2(new_n296_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n558_), .A2(new_n526_), .A3(new_n471_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n472_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G113gat), .B1(new_n807_), .B2(new_n579_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n804_), .A2(new_n296_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n766_), .ZN(new_n810_));
  OR3_X1    g609(.A1(new_n806_), .A2(KEYINPUT119), .A3(new_n472_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT119), .B1(new_n806_), .B2(new_n472_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n810_), .A2(KEYINPUT120), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n805_), .B2(new_n814_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n816_), .B(new_n818_), .C1(new_n807_), .C2(new_n812_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n579_), .A2(G113gat), .ZN(new_n821_));
  XOR2_X1   g620(.A(new_n821_), .B(KEYINPUT121), .Z(new_n822_));
  AOI21_X1  g621(.A(new_n808_), .B1(new_n820_), .B2(new_n822_), .ZN(G1340gat));
  OAI21_X1  g622(.A(G120gat), .B1(new_n819_), .B2(new_n698_), .ZN(new_n824_));
  INV_X1    g623(.A(G120gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n698_), .B2(KEYINPUT60), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n807_), .B(new_n826_), .C1(KEYINPUT60), .C2(new_n825_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n827_), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n807_), .B2(new_n297_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n297_), .A2(G127gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT122), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n820_), .B2(new_n831_), .ZN(G1342gat));
  OAI21_X1  g631(.A(G134gat), .B1(new_n819_), .B2(new_n264_), .ZN(new_n833_));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n807_), .A2(new_n834_), .A3(new_n256_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1343gat));
  NOR2_X1   g635(.A1(new_n805_), .A2(new_n472_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n558_), .A2(new_n522_), .A3(new_n471_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n579_), .A3(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT123), .B(G141gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n838_), .ZN(new_n842_));
  OR3_X1    g641(.A1(new_n842_), .A2(G148gat), .A3(new_n698_), .ZN(new_n843_));
  OAI21_X1  g642(.A(G148gat), .B1(new_n842_), .B2(new_n698_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1345gat));
  XNOR2_X1  g644(.A(KEYINPUT61), .B(G155gat), .ZN(new_n846_));
  OR3_X1    g645(.A1(new_n842_), .A2(new_n296_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n842_), .B2(new_n296_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1346gat));
  OAI21_X1  g648(.A(G162gat), .B1(new_n842_), .B2(new_n264_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n256_), .A2(new_n305_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n842_), .B2(new_n851_), .ZN(G1347gat));
  NOR3_X1   g651(.A1(new_n421_), .A2(new_n473_), .A3(new_n526_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR4_X1   g653(.A1(new_n805_), .A2(KEYINPUT22), .A3(new_n580_), .A4(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n856_));
  OR3_X1    g655(.A1(new_n855_), .A2(new_n856_), .A3(G169gat), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n805_), .A2(new_n854_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n856_), .A3(new_n579_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n859_), .B(G169gat), .C1(new_n856_), .C2(new_n855_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n857_), .A2(new_n860_), .ZN(G1348gat));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n699_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n424_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT124), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n862_), .A2(new_n865_), .A3(new_n424_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT125), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n862_), .B2(new_n424_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n858_), .A2(KEYINPUT125), .A3(G176gat), .A4(new_n699_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n864_), .A2(new_n866_), .B1(new_n868_), .B2(new_n869_), .ZN(G1349gat));
  NAND2_X1  g669(.A1(new_n858_), .A2(new_n297_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n484_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n436_), .B2(new_n871_), .ZN(G1350gat));
  INV_X1    g672(.A(new_n858_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G190gat), .B1(new_n874_), .B2(new_n264_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n858_), .A2(new_n256_), .A3(new_n485_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1351gat));
  NAND3_X1  g676(.A1(new_n525_), .A2(new_n522_), .A3(new_n612_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n805_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n579_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n699_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n297_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  AND2_X1   g684(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n884_), .B2(new_n885_), .ZN(G1354gat));
  OR2_X1    g687(.A1(new_n805_), .A2(new_n878_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT127), .B(G218gat), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n889_), .A2(new_n264_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT126), .B1(new_n889_), .B2(new_n259_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n879_), .A2(new_n893_), .A3(new_n256_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n891_), .B1(new_n895_), .B2(new_n890_), .ZN(G1355gat));
endmodule


