//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(G99gat), .ZN(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT64), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n217_), .A2(new_n206_), .A3(new_n207_), .A4(new_n208_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n210_), .A2(new_n215_), .A3(new_n216_), .A4(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G85gat), .ZN(new_n220_));
  INV_X1    g019(.A(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(G71gat), .A2(G78gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G71gat), .A2(G78gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G57gat), .B(G64gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(KEYINPUT11), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n231_), .B2(KEYINPUT11), .ZN(new_n234_));
  INV_X1    g033(.A(G64gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G57gat), .ZN(new_n236_));
  INV_X1    g035(.A(G57gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G64gat), .ZN(new_n238_));
  AND4_X1   g037(.A1(new_n233_), .A2(new_n236_), .A3(new_n238_), .A4(KEYINPUT11), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n232_), .B1(new_n234_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(new_n238_), .A3(KEYINPUT11), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT65), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n238_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n236_), .A2(new_n238_), .A3(new_n233_), .A4(KEYINPUT11), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n242_), .A2(new_n245_), .A3(new_n230_), .A4(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n240_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n219_), .A2(KEYINPUT8), .A3(new_n224_), .ZN(new_n249_));
  OR2_X1    g048(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n208_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n222_), .A2(KEYINPUT9), .A3(new_n223_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n223_), .A2(KEYINPUT9), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n215_), .A2(new_n252_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n227_), .A2(new_n248_), .A3(new_n249_), .A4(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G230gat), .A2(G233gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT67), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(new_n260_), .A3(new_n257_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n227_), .A2(new_n255_), .A3(new_n249_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n248_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n263_), .A2(KEYINPUT12), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT12), .B1(new_n263_), .B2(new_n264_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n249_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT8), .B1(new_n219_), .B2(new_n224_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n255_), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(new_n248_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n257_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n263_), .A2(new_n264_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(KEYINPUT66), .A3(new_n256_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n262_), .A2(new_n267_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n205_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n276_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n271_), .B2(new_n248_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n263_), .A2(KEYINPUT12), .A3(new_n264_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n256_), .A2(new_n260_), .A3(new_n257_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n260_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n282_), .B(new_n283_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(KEYINPUT68), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n279_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n205_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT69), .B1(new_n277_), .B2(new_n290_), .ZN(new_n291_));
  AND4_X1   g090(.A1(KEYINPUT69), .A2(new_n280_), .A3(new_n286_), .A4(new_n290_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT13), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(KEYINPUT13), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G232gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT34), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT35), .ZN(new_n300_));
  XOR2_X1   g099(.A(G29gat), .B(G36gat), .Z(new_n301_));
  XOR2_X1   g100(.A(G43gat), .B(G50gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT15), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n300_), .B1(new_n304_), .B2(new_n263_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n303_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n305_), .B1(new_n306_), .B2(new_n263_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n299_), .A2(KEYINPUT35), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G190gat), .B(G218gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G134gat), .B(G162gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n312_), .A2(KEYINPUT36), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n312_), .B(KEYINPUT36), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n309_), .A2(new_n317_), .ZN(new_n318_));
  OR3_X1    g117(.A1(new_n315_), .A2(new_n318_), .A3(KEYINPUT37), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT37), .B1(new_n315_), .B2(new_n318_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G15gat), .B(G22gat), .ZN(new_n323_));
  INV_X1    g122(.A(G1gat), .ZN(new_n324_));
  INV_X1    g123(.A(G8gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT14), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G1gat), .B(G8gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G231gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(new_n248_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G127gat), .B(G155gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT70), .B(KEYINPUT16), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G183gat), .B(G211gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT17), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n337_), .A2(KEYINPUT17), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n332_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n332_), .A2(new_n338_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT71), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n297_), .A2(new_n322_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n344_), .A2(new_n345_), .ZN(new_n347_));
  XOR2_X1   g146(.A(KEYINPUT84), .B(G204gat), .Z(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(G197gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G197gat), .ZN(new_n353_));
  OAI22_X1  g152(.A1(new_n349_), .A2(new_n350_), .B1(new_n353_), .B2(G204gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT21), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G197gat), .A2(G204gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT84), .B(G204gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(G197gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(KEYINPUT21), .ZN(new_n359_));
  XOR2_X1   g158(.A(G211gat), .B(G218gat), .Z(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(KEYINPUT21), .A3(new_n360_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n370_));
  INV_X1    g169(.A(G141gat), .ZN(new_n371_));
  INV_X1    g170(.A(G148gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G141gat), .A2(G148gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT80), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n373_), .B(new_n374_), .C1(new_n376_), .C2(KEYINPUT2), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n376_), .A2(KEYINPUT2), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n369_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT81), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n366_), .A2(KEYINPUT1), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n366_), .B1(new_n368_), .B2(KEYINPUT1), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n384_), .B2(new_n383_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n371_), .A2(new_n372_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n375_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT29), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n365_), .B1(KEYINPUT86), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(KEYINPUT86), .B2(new_n390_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(G228gat), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n392_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n389_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT29), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n396_), .B(new_n364_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G22gat), .B(G50gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n398_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n400_), .A2(new_n401_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n407_), .A2(KEYINPUT28), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n409_), .B(KEYINPUT87), .Z(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(KEYINPUT28), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n408_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n411_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n415_));
  OAI22_X1  g214(.A1(new_n405_), .A2(new_n406_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n398_), .A2(new_n402_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n403_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n415_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n398_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n413_), .A4(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT90), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G169gat), .A2(G176gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT24), .ZN(new_n431_));
  OR3_X1    g230(.A1(KEYINPUT75), .A2(G169gat), .A3(G176gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  MUX2_X1   g233(.A(KEYINPUT24), .B(new_n431_), .S(new_n434_), .Z(new_n435_));
  INV_X1    g234(.A(G183gat), .ZN(new_n436_));
  INV_X1    g235(.A(G190gat), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n436_), .A2(new_n437_), .A3(KEYINPUT23), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT23), .B1(new_n436_), .B2(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT25), .B(G183gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT26), .B(G190gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n435_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT22), .B(G169gat), .ZN(new_n446_));
  INV_X1    g245(.A(G176gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT76), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n440_), .B(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(new_n438_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G183gat), .A2(G190gat), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n448_), .B(new_n430_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n445_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n429_), .B1(new_n364_), .B2(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n450_), .A2(new_n438_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT74), .B1(new_n436_), .B2(KEYINPUT25), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n443_), .B(new_n457_), .C1(new_n442_), .C2(KEYINPUT74), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n435_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n448_), .B(KEYINPUT77), .Z(new_n460_));
  OAI21_X1  g259(.A(new_n441_), .B1(G183gat), .B2(G190gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n430_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n455_), .B1(new_n364_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G226gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT19), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n445_), .A2(new_n453_), .A3(KEYINPUT92), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n454_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n365_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n429_), .B1(new_n364_), .B2(new_n463_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n468_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(KEYINPUT32), .B(new_n428_), .C1(new_n467_), .C2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n364_), .A2(new_n454_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n476_), .A2(KEYINPUT88), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(KEYINPUT88), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n468_), .B(new_n473_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n464_), .A2(new_n466_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n428_), .A2(KEYINPUT32), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n475_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G225gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n389_), .B(KEYINPUT82), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G127gat), .B(G134gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G113gat), .B(G120gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(new_n490_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n389_), .A2(new_n490_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n485_), .B(new_n491_), .C1(new_n494_), .C2(new_n487_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n492_), .A2(new_n493_), .A3(new_n484_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G1gat), .B(G29gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G85gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT0), .B(G57gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  AND3_X1   g299(.A1(new_n495_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n483_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT93), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n479_), .A2(new_n428_), .A3(new_n480_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n428_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n495_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT33), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT33), .A4(new_n500_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n500_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(new_n494_), .B2(new_n484_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT91), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n491_), .B(new_n484_), .C1(new_n494_), .C2(new_n487_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n517_), .B(new_n513_), .C1(new_n494_), .C2(new_n484_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n508_), .A2(new_n511_), .A3(new_n512_), .A4(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n483_), .B(new_n521_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n422_), .A2(new_n504_), .A3(new_n520_), .A4(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G71gat), .B(G99gat), .ZN(new_n524_));
  INV_X1    g323(.A(G43gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G227gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(G15gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n526_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n463_), .B(KEYINPUT30), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT78), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n530_), .A2(new_n531_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n529_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n532_), .B2(new_n529_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n490_), .B(KEYINPUT31), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n535_), .B(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n501_), .A2(new_n502_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT27), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n540_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n467_), .A2(new_n474_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n505_), .B(KEYINPUT27), .C1(new_n428_), .C2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n539_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n416_), .A2(new_n421_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n538_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n543_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n539_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n535_), .B(new_n536_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n523_), .A2(new_n546_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n304_), .A2(new_n329_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n327_), .B(new_n328_), .Z(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n303_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n553_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n306_), .A2(new_n329_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT73), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(new_n558_), .A3(KEYINPUT73), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n556_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n557_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G169gat), .B(G197gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n567_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n557_), .B2(new_n563_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR4_X1   g371(.A1(new_n346_), .A2(new_n347_), .A3(new_n552_), .A4(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n324_), .A3(new_n549_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT38), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT95), .B1(new_n315_), .B2(new_n318_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n314_), .B(new_n578_), .C1(new_n309_), .C2(new_n317_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n552_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n297_), .A2(new_n572_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT94), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n581_), .A2(new_n584_), .A3(new_n342_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n324_), .B1(new_n585_), .B2(new_n549_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n576_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n575_), .B2(new_n574_), .ZN(G1324gat));
  NAND3_X1  g387(.A1(new_n573_), .A2(new_n325_), .A3(new_n547_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n547_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(G8gat), .ZN(new_n592_));
  AOI211_X1 g391(.A(KEYINPUT39), .B(new_n325_), .C1(new_n585_), .C2(new_n547_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n589_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT40), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(G1325gat));
  INV_X1    g395(.A(G15gat), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n585_), .B2(new_n538_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT41), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n573_), .A2(new_n597_), .A3(new_n538_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(G1326gat));
  INV_X1    g400(.A(G22gat), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n585_), .B2(new_n545_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT42), .Z(new_n604_));
  NAND3_X1  g403(.A1(new_n573_), .A2(new_n602_), .A3(new_n545_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(G1327gat));
  OAI21_X1  g405(.A(KEYINPUT43), .B1(new_n321_), .B2(KEYINPUT96), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n523_), .A2(new_n546_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n548_), .A2(new_n551_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n322_), .B(new_n608_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n552_), .B2(new_n321_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n343_), .A4(new_n584_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT44), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT97), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n613_), .A2(new_n617_), .A3(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n613_), .A2(new_n614_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n549_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G29gat), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n552_), .A2(new_n572_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n297_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n580_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n343_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n624_), .A2(new_n625_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT98), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n624_), .A2(new_n631_), .A3(new_n625_), .A4(new_n628_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n539_), .A2(G29gat), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT99), .Z(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n623_), .A2(new_n636_), .ZN(G1328gat));
  INV_X1    g436(.A(new_n547_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(G36gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n630_), .A2(new_n632_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT45), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT45), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n630_), .A2(new_n642_), .A3(new_n632_), .A4(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n547_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n646_));
  INV_X1    g445(.A(G36gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n644_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT46), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n644_), .B(KEYINPUT46), .C1(new_n646_), .C2(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1329gat));
  NAND2_X1  g451(.A1(new_n633_), .A2(new_n538_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n525_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n550_), .A2(new_n525_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n618_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n617_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n621_), .B(new_n655_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n654_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT47), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT47), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n654_), .A2(new_n658_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1330gat));
  INV_X1    g462(.A(G50gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n633_), .A2(new_n664_), .A3(new_n545_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n620_), .A2(new_n422_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n619_), .A2(KEYINPUT100), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G50gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT100), .B1(new_n619_), .B2(new_n666_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1331gat));
  NAND2_X1  g469(.A1(new_n297_), .A2(new_n572_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n552_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n343_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT101), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n237_), .A3(new_n549_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n671_), .A2(new_n343_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n581_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G57gat), .B1(new_n679_), .B2(new_n539_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(G1332gat));
  AOI21_X1  g480(.A(new_n235_), .B1(new_n678_), .B2(new_n547_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT48), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n675_), .A2(new_n235_), .A3(new_n547_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1333gat));
  INV_X1    g484(.A(G71gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n678_), .B2(new_n538_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT49), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n675_), .A2(new_n686_), .A3(new_n538_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1334gat));
  INV_X1    g489(.A(G78gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n675_), .A2(new_n691_), .A3(new_n545_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT50), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n678_), .A2(new_n545_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G78gat), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT50), .B(new_n691_), .C1(new_n678_), .C2(new_n545_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT102), .ZN(G1335gat));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n672_), .B2(new_n628_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n628_), .ZN(new_n701_));
  NOR4_X1   g500(.A1(new_n552_), .A2(KEYINPUT103), .A3(new_n701_), .A4(new_n671_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G85gat), .B1(new_n703_), .B2(new_n549_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n612_), .A2(new_n343_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n671_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n611_), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n539_), .A2(new_n220_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT104), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n704_), .B1(new_n708_), .B2(new_n710_), .ZN(G1336gat));
  OAI21_X1  g510(.A(G92gat), .B1(new_n707_), .B2(new_n638_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n703_), .A2(new_n221_), .A3(new_n547_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT105), .Z(G1337gat));
  AND3_X1   g514(.A1(new_n538_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717_));
  AOI22_X1  g516(.A1(new_n703_), .A2(new_n716_), .B1(new_n717_), .B2(KEYINPUT51), .ZN(new_n718_));
  OAI21_X1  g517(.A(G99gat), .B1(new_n707_), .B2(new_n550_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n717_), .A2(KEYINPUT51), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1338gat));
  OAI21_X1  g521(.A(G106gat), .B1(new_n707_), .B2(new_n422_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n422_), .A2(G106gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n726_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT52), .B(G106gat), .C1(new_n707_), .C2(new_n422_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n725_), .A2(new_n729_), .A3(new_n730_), .A4(new_n732_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1339gat));
  INV_X1    g535(.A(KEYINPUT58), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n291_), .A2(new_n292_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT114), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n561_), .A2(new_n562_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n556_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n556_), .B1(new_n554_), .B2(new_n303_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n567_), .B1(new_n553_), .B2(new_n742_), .ZN(new_n743_));
  AOI22_X1  g542(.A1(new_n564_), .A2(new_n567_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n738_), .A2(new_n739_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT56), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n257_), .B1(new_n267_), .B2(new_n256_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n284_), .A2(new_n285_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n282_), .A2(new_n283_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT55), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n262_), .A2(new_n751_), .A3(new_n267_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n747_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n746_), .B1(new_n753_), .B2(new_n290_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n290_), .A2(new_n746_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n753_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n745_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n739_), .B1(new_n738_), .B2(new_n744_), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT115), .B(new_n737_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n759_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n737_), .A2(KEYINPUT115), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n757_), .A4(new_n745_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(new_n322_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n753_), .B2(new_n756_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n256_), .ZN(new_n768_));
  OAI211_X1 g567(.A(G230gat), .B(G233gat), .C1(new_n749_), .C2(new_n768_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n748_), .A2(KEYINPUT55), .A3(new_n749_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n751_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(KEYINPUT112), .A3(new_n755_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n754_), .A2(new_n767_), .A3(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n571_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n571_), .B(KEYINPUT111), .C1(new_n291_), .C2(new_n292_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n774_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n744_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n580_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n765_), .B1(new_n781_), .B2(KEYINPUT113), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n783_), .B(new_n580_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n764_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n781_), .A2(KEYINPUT57), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n342_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n673_), .A2(new_n295_), .A3(new_n572_), .A4(new_n296_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT54), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n791_), .A2(KEYINPUT110), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(KEYINPUT110), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n795_));
  OR3_X1    g594(.A1(new_n790_), .A2(new_n795_), .A3(KEYINPUT54), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n790_), .B2(KEYINPUT54), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n794_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n789_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n548_), .A2(new_n549_), .A3(new_n538_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT59), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n786_), .B1(new_n785_), .B2(KEYINPUT116), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n764_), .B(new_n806_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n627_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n792_), .A2(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n801_), .A2(KEYINPUT59), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n804_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n572_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n572_), .A2(G113gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n803_), .B2(new_n814_), .ZN(G1340gat));
  OAI21_X1  g614(.A(G120gat), .B1(new_n812_), .B2(new_n625_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT60), .ZN(new_n817_));
  AOI21_X1  g616(.A(G120gat), .B1(new_n297_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n817_), .B2(G120gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n800_), .A2(new_n802_), .A3(new_n819_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT117), .Z(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(new_n821_), .ZN(G1341gat));
  INV_X1    g621(.A(G127gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n803_), .B2(new_n343_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT118), .B(new_n823_), .C1(new_n803_), .C2(new_n343_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n810_), .A2(new_n811_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n803_), .B2(KEYINPUT59), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n788_), .A2(new_n823_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n830_), .B2(new_n831_), .ZN(G1342gat));
  INV_X1    g631(.A(G134gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n321_), .A2(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT119), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n800_), .A2(new_n580_), .A3(new_n802_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n830_), .A2(new_n835_), .B1(new_n833_), .B2(new_n836_), .ZN(G1343gat));
  AOI21_X1  g636(.A(new_n809_), .B1(new_n788_), .B2(new_n787_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n422_), .A2(new_n538_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n638_), .A3(new_n549_), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(KEYINPUT120), .Z(new_n841_));
  NOR2_X1   g640(.A1(new_n838_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n571_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n297_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n842_), .A2(new_n849_), .A3(new_n627_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n842_), .B2(new_n627_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n848_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n852_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n850_), .A3(new_n847_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1346gat));
  AOI21_X1  g655(.A(G162gat), .B1(new_n842_), .B2(new_n580_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n322_), .A2(G162gat), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(KEYINPUT122), .Z(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n842_), .B2(new_n859_), .ZN(G1347gat));
  NOR2_X1   g659(.A1(new_n638_), .A2(new_n549_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n422_), .A3(new_n538_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n571_), .B(new_n863_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n446_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(G169gat), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT123), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n866_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n867_), .A2(KEYINPUT123), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(KEYINPUT62), .A3(new_n868_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1348gat));
  NAND4_X1  g673(.A1(new_n800_), .A2(G176gat), .A3(new_n297_), .A4(new_n863_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n810_), .A2(new_n625_), .A3(new_n862_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(G176gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT124), .ZN(G1349gat));
  NOR2_X1   g677(.A1(new_n838_), .A2(new_n862_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G183gat), .B1(new_n879_), .B2(new_n627_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n810_), .A2(new_n862_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n788_), .A2(new_n442_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(G1350gat));
  NAND3_X1  g682(.A1(new_n881_), .A2(new_n443_), .A3(new_n580_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n322_), .B(new_n863_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n885_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT125), .B1(new_n885_), .B2(G190gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT126), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n884_), .B(new_n890_), .C1(new_n886_), .C2(new_n887_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1351gat));
  NAND2_X1  g691(.A1(new_n839_), .A2(new_n861_), .ZN(new_n893_));
  OR3_X1    g692(.A1(new_n838_), .A2(KEYINPUT127), .A3(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT127), .B1(new_n838_), .B2(new_n893_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G197gat), .B1(new_n896_), .B2(new_n571_), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n353_), .B(new_n572_), .C1(new_n894_), .C2(new_n895_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1352gat));
  AOI21_X1  g698(.A(G204gat), .B1(new_n896_), .B2(new_n297_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n348_), .B(new_n625_), .C1(new_n894_), .C2(new_n895_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1353gat));
  OR2_X1    g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n896_), .B2(new_n342_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT63), .B(G211gat), .ZN(new_n905_));
  AOI211_X1 g704(.A(new_n788_), .B(new_n905_), .C1(new_n894_), .C2(new_n895_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1354gat));
  INV_X1    g706(.A(G218gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n896_), .A2(new_n908_), .A3(new_n580_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n321_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n908_), .B2(new_n910_), .ZN(G1355gat));
endmodule


