//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT72), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G190gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(G218gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(G218gat), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n207_), .A2(KEYINPUT36), .A3(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT36), .B1(new_n207_), .B2(new_n208_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G232gat), .A2(G233gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT34), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT35), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AND3_X1   g016(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G85gat), .ZN(new_n225_));
  INV_X1    g024(.A(G92gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT9), .A3(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(KEYINPUT9), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n220_), .A2(new_n224_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  AND4_X1   g032(.A1(new_n220_), .A2(new_n224_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT67), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n227_), .A2(new_n228_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G99gat), .A2(G106gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT6), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n241_));
  NOR3_X1   g040(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT7), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n240_), .B(new_n241_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n245_));
  INV_X1    g044(.A(G99gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n222_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(KEYINPUT7), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n236_), .B(new_n237_), .C1(new_n244_), .C2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(KEYINPUT7), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n242_), .A2(new_n243_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(new_n220_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n236_), .B1(new_n253_), .B2(new_n237_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n233_), .B(new_n235_), .C1(new_n250_), .C2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G29gat), .B(G36gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G43gat), .B(G50gat), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n257_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT15), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT15), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n256_), .A2(new_n257_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n256_), .A2(new_n257_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n255_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT71), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n255_), .A2(new_n268_), .A3(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n258_), .A2(new_n259_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n271_), .B(new_n231_), .C1(new_n250_), .C2(new_n254_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(KEYINPUT35), .B2(new_n213_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n217_), .B1(new_n270_), .B2(new_n274_), .ZN(new_n275_));
  AOI211_X1 g074(.A(new_n216_), .B(new_n273_), .C1(new_n267_), .C2(new_n269_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n203_), .B(new_n211_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n269_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n268_), .B1(new_n255_), .B2(new_n265_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n274_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n216_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n270_), .A2(new_n217_), .A3(new_n274_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(new_n210_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n282_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n203_), .B1(new_n285_), .B2(new_n211_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n202_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n211_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n285_), .A2(KEYINPUT73), .A3(new_n211_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT37), .A4(new_n283_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G127gat), .B(G155gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT16), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G183gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(G211gat), .Z(new_n297_));
  INV_X1    g096(.A(KEYINPUT17), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT14), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT75), .B(G8gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(G1gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(G15gat), .B(G22gat), .Z(new_n305_));
  NOR3_X1   g104(.A1(new_n304_), .A2(KEYINPUT76), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307_));
  AND2_X1   g106(.A1(KEYINPUT75), .A2(G8gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(KEYINPUT75), .A2(G8gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(G1gat), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT14), .ZN(new_n311_));
  INV_X1    g110(.A(new_n305_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n307_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n301_), .B1(new_n306_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT76), .B1(new_n304_), .B2(new_n305_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n312_), .A3(new_n307_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n300_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G231gat), .A3(G233gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G231gat), .A2(G233gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n314_), .A2(new_n320_), .A3(new_n317_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G71gat), .B(G78gat), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G64gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G57gat), .ZN(new_n326_));
  INV_X1    g125(.A(G57gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G64gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT66), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT66), .B1(new_n326_), .B2(new_n328_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n324_), .B(KEYINPUT11), .C1(new_n329_), .C2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT11), .B1(new_n329_), .B2(new_n330_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT66), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n327_), .A2(G64gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n325_), .A2(G57gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT11), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT66), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n332_), .A2(new_n339_), .A3(new_n323_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n322_), .A2(new_n331_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n331_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n319_), .A2(new_n342_), .A3(new_n321_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n299_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n343_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n345_), .A2(new_n298_), .A3(new_n297_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n293_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT77), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G230gat), .A2(G233gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n351_), .B(KEYINPUT64), .Z(new_n352_));
  OAI21_X1  g151(.A(new_n237_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT8), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n234_), .B1(new_n354_), .B2(new_n249_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n342_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(new_n342_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n352_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n355_), .B2(new_n342_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n352_), .B1(new_n355_), .B2(new_n342_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n340_), .A2(KEYINPUT12), .A3(new_n331_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n255_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n366_));
  XNOR2_X1  g165(.A(G120gat), .B(G148gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G176gat), .B(G204gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n359_), .A2(new_n365_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n359_), .B2(new_n365_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT13), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT13), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT70), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G113gat), .B(G141gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(G169gat), .ZN(new_n381_));
  INV_X1    g180(.A(G197gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n314_), .A2(new_n271_), .A3(new_n317_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G229gat), .A2(G233gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n315_), .A2(new_n300_), .A3(new_n316_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n300_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n265_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT78), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n318_), .A2(new_n392_), .A3(new_n265_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n387_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n386_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n271_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n388_), .A2(new_n389_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n271_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n395_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n384_), .B1(new_n394_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n260_), .A2(new_n264_), .ZN(new_n402_));
  AOI211_X1 g201(.A(KEYINPUT78), .B(new_n402_), .C1(new_n314_), .C2(new_n317_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n392_), .B1(new_n318_), .B2(new_n265_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n399_), .B(new_n383_), .C1(new_n405_), .C2(new_n387_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n401_), .A2(new_n406_), .A3(KEYINPUT79), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n408_), .B(new_n384_), .C1(new_n394_), .C2(new_n400_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n350_), .A2(new_n379_), .A3(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT3), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT2), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G155gat), .B(G162gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n417_), .A2(KEYINPUT1), .ZN(new_n420_));
  INV_X1    g219(.A(new_n412_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n414_), .A3(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n419_), .A2(KEYINPUT88), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n417_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n420_), .A2(new_n423_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT28), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n431_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT89), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n432_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT28), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n433_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G22gat), .B(G50gat), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n436_), .A2(new_n442_), .A3(new_n440_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(KEYINPUT92), .A3(new_n445_), .ZN(new_n446_));
  OR3_X1    g245(.A1(new_n382_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n447_));
  INV_X1    g246(.A(G204gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G197gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT91), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n382_), .A2(G204gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n447_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G211gat), .B(G218gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT21), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n451_), .B2(new_n449_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT90), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n453_), .B1(new_n452_), .B2(KEYINPUT21), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n456_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G228gat), .A2(G233gat), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n460_), .B(new_n461_), .C1(new_n430_), .C2(new_n432_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n460_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n427_), .A2(new_n428_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(new_n432_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n462_), .B1(new_n466_), .B2(new_n461_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G78gat), .B(G106gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n446_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n471_));
  INV_X1    g270(.A(new_n445_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n442_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(new_n446_), .A3(new_n469_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G15gat), .B(G43gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G227gat), .A2(G233gat), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G71gat), .B(G99gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n481_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n483_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n477_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n480_), .B(new_n481_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n483_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(KEYINPUT86), .A3(new_n485_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G169gat), .A2(G176gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(KEYINPUT22), .B(G169gat), .Z(new_n494_));
  OAI21_X1  g293(.A(new_n493_), .B1(new_n494_), .B2(G176gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT80), .B(G183gat), .Z(new_n496_));
  XOR2_X1   g295(.A(KEYINPUT81), .B(G190gat), .Z(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G183gat), .A2(G190gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT23), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT23), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(G183gat), .A3(G190gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n503_), .A2(KEYINPUT83), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT83), .B1(new_n499_), .B2(KEYINPUT23), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n498_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT84), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n495_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OAI211_X1 g307(.A(KEYINPUT84), .B(new_n498_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(G169gat), .A2(G176gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT82), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(KEYINPUT24), .A3(new_n493_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n511_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT24), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n513_), .A2(new_n503_), .A3(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n496_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT26), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n497_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n524_));
  OAI22_X1  g323(.A1(new_n519_), .A2(new_n521_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n518_), .A2(new_n525_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n510_), .A2(KEYINPUT30), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT30), .B1(new_n510_), .B2(new_n526_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n488_), .B(new_n492_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT87), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n510_), .A2(new_n526_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n508_), .A2(new_n509_), .B1(new_n525_), .B2(new_n518_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT30), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT86), .B1(new_n491_), .B2(new_n485_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n529_), .A2(new_n530_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT31), .ZN(new_n539_));
  XOR2_X1   g338(.A(G127gat), .B(G134gat), .Z(new_n540_));
  XOR2_X1   g339(.A(G113gat), .B(G120gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT31), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n529_), .A2(new_n530_), .A3(new_n537_), .A4(new_n544_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n539_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n476_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n470_), .B(new_n475_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT27), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G8gat), .B(G36gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT18), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G64gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(new_n226_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n510_), .A2(new_n463_), .A3(new_n526_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT25), .B(G183gat), .Z(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT26), .B(G190gat), .Z(new_n559_));
  OAI21_X1  g358(.A(new_n513_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n505_), .B1(new_n503_), .B2(KEYINPUT83), .ZN(new_n561_));
  NOR3_X1   g360(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n561_), .A2(KEYINPUT94), .A3(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT94), .B1(new_n561_), .B2(new_n562_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n560_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n503_), .B1(G183gat), .B2(G190gat), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(new_n567_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n495_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n460_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n557_), .A2(new_n571_), .A3(KEYINPUT20), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G226gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT19), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT93), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n534_), .A2(new_n463_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n565_), .A2(new_n570_), .A3(new_n460_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT20), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n574_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(KEYINPUT96), .A2(new_n576_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n575_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n579_), .B1(new_n534_), .B2(new_n463_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n584_), .B2(new_n571_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n556_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n576_), .A2(KEYINPUT96), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n578_), .A2(new_n579_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n531_), .A2(new_n460_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n581_), .A3(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n587_), .A2(new_n589_), .A3(new_n556_), .A4(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n552_), .B1(new_n588_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n582_), .A2(KEYINPUT99), .A3(new_n556_), .A4(new_n587_), .ZN(new_n598_));
  OAI22_X1  g397(.A1(new_n580_), .A2(new_n581_), .B1(new_n575_), .B2(new_n572_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n556_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n552_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n598_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n595_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G1gat), .B(G29gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT0), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(new_n327_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(new_n225_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G225gat), .A2(G233gat), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n425_), .A2(new_n429_), .A3(new_n543_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(KEYINPUT4), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n464_), .A2(new_n542_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n613_), .A2(KEYINPUT97), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(KEYINPUT97), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(KEYINPUT4), .A3(new_n611_), .A4(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n612_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n613_), .B(KEYINPUT97), .Z(new_n619_));
  NAND4_X1  g418(.A1(new_n619_), .A2(KEYINPUT98), .A3(KEYINPUT4), .A4(new_n611_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n610_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n610_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n619_), .B2(new_n611_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n609_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n621_), .A2(new_n609_), .A3(new_n623_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n551_), .A2(new_n604_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n556_), .A2(KEYINPUT32), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n582_), .A2(new_n587_), .A3(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n599_), .A2(KEYINPUT32), .A3(new_n556_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n630_), .B(new_n631_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n624_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT33), .B(new_n609_), .C1(new_n621_), .C2(new_n623_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n618_), .A2(new_n620_), .A3(new_n610_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n619_), .A2(new_n622_), .A3(new_n611_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n608_), .A3(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n634_), .A2(new_n635_), .A3(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n588_), .A2(new_n594_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n632_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n548_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n628_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n411_), .A2(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n645_), .A2(G1gat), .A3(new_n627_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n625_), .A2(new_n626_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n648_));
  AOI22_X1  g447(.A1(new_n648_), .A2(new_n604_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n284_), .A2(new_n286_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n378_), .A2(new_n410_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n348_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n647_), .A3(new_n654_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n646_), .A2(KEYINPUT38), .B1(new_n655_), .B2(G1gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n646_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n657_), .A2(KEYINPUT100), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT100), .B1(new_n657_), .B2(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(G1324gat));
  NAND3_X1  g460(.A1(new_n651_), .A2(new_n603_), .A3(new_n654_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n662_), .A2(new_n663_), .A3(G8gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n662_), .B2(G8gat), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n604_), .A2(new_n303_), .ZN(new_n666_));
  OAI22_X1  g465(.A1(new_n664_), .A2(new_n665_), .B1(new_n645_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1325gat));
  NAND3_X1  g468(.A1(new_n651_), .A2(new_n548_), .A3(new_n654_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n670_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT41), .B1(new_n670_), .B2(G15gat), .ZN(new_n672_));
  INV_X1    g471(.A(new_n547_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n539_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(G15gat), .ZN(new_n676_));
  OAI22_X1  g475(.A1(new_n671_), .A2(new_n672_), .B1(new_n645_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT101), .ZN(G1326gat));
  OR3_X1    g477(.A1(new_n645_), .A2(G22gat), .A3(new_n476_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n651_), .A2(new_n654_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G22gat), .B1(new_n680_), .B2(new_n476_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT102), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n683_), .B(G22gat), .C1(new_n680_), .C2(new_n476_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n682_), .A2(KEYINPUT42), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT42), .B1(new_n682_), .B2(new_n684_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n679_), .B1(new_n685_), .B2(new_n686_), .ZN(G1327gat));
  NOR2_X1   g486(.A1(new_n653_), .A2(new_n347_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n644_), .B2(new_n293_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n293_), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT43), .B(new_n691_), .C1(new_n628_), .C2(new_n643_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n688_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n649_), .B2(new_n691_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n644_), .A2(new_n689_), .A3(new_n293_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT44), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n695_), .A2(new_n700_), .A3(new_n647_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G29gat), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n647_), .B(new_n603_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n641_), .A2(new_n642_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n650_), .B(new_n688_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT103), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n644_), .A2(new_n707_), .A3(new_n650_), .A4(new_n688_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n627_), .A2(G29gat), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT104), .Z(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n702_), .A2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  INV_X1    g513(.A(G36gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n604_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(new_n700_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n604_), .A2(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n706_), .A2(new_n708_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n714_), .B1(new_n717_), .B2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n603_), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n693_), .A2(new_n694_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G36gat), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n719_), .B(KEYINPUT45), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(KEYINPUT46), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n722_), .A2(new_n727_), .ZN(G1329gat));
  NAND3_X1  g527(.A1(new_n706_), .A2(new_n548_), .A3(new_n708_), .ZN(new_n729_));
  INV_X1    g528(.A(G43gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(G43gat), .B(new_n548_), .C1(new_n699_), .C2(KEYINPUT44), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(new_n724_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g533(.A(new_n476_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G50gat), .B1(new_n709_), .B2(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n695_), .A2(G50gat), .A3(new_n735_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n700_), .ZN(G1331gat));
  INV_X1    g537(.A(new_n379_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n410_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n739_), .A2(new_n348_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n651_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n627_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n378_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n350_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT105), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n649_), .A2(new_n740_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n647_), .A2(new_n327_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n743_), .B1(new_n748_), .B2(new_n749_), .ZN(G1332gat));
  NAND2_X1  g549(.A1(new_n603_), .A2(new_n325_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n651_), .A2(new_n603_), .A3(new_n741_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G64gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G64gat), .ZN(new_n755_));
  OAI22_X1  g554(.A1(new_n748_), .A2(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT106), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n758_));
  OAI221_X1 g557(.A(new_n758_), .B1(new_n754_), .B2(new_n755_), .C1(new_n748_), .C2(new_n751_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1333gat));
  OAI21_X1  g559(.A(G71gat), .B1(new_n742_), .B2(new_n675_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(KEYINPUT49), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(KEYINPUT49), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n675_), .A2(G71gat), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n762_), .A2(new_n763_), .B1(new_n748_), .B2(new_n764_), .ZN(G1334gat));
  NAND3_X1  g564(.A1(new_n651_), .A2(new_n735_), .A3(new_n741_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(G78gat), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n767_), .A2(new_n769_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n476_), .A2(G78gat), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n770_), .A2(new_n771_), .B1(new_n748_), .B2(new_n772_), .ZN(G1335gat));
  INV_X1    g572(.A(new_n650_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n649_), .A2(new_n774_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n739_), .A2(new_n347_), .A3(new_n740_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n647_), .A3(new_n776_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n777_), .A2(KEYINPUT108), .A3(new_n225_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT108), .B1(new_n777_), .B2(new_n225_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n744_), .A2(new_n347_), .A3(new_n740_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n647_), .A2(G85gat), .ZN(new_n782_));
  OAI22_X1  g581(.A1(new_n778_), .A2(new_n779_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT109), .ZN(G1336gat));
  AND2_X1   g583(.A1(new_n775_), .A2(new_n776_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G92gat), .B1(new_n785_), .B2(new_n603_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n781_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n603_), .A2(G92gat), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT110), .Z(new_n789_));
  AOI21_X1  g588(.A(new_n786_), .B1(new_n787_), .B2(new_n789_), .ZN(G1337gat));
  NAND4_X1  g589(.A1(new_n785_), .A2(new_n548_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n781_), .A2(new_n675_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n246_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g593(.A1(new_n785_), .A2(new_n222_), .A3(new_n735_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n735_), .B(new_n780_), .C1(new_n690_), .C2(new_n692_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(G106gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n796_), .B2(G106gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n795_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1339gat));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n365_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n361_), .A2(new_n364_), .A3(new_n356_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n352_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .A4(KEYINPUT55), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n370_), .A2(new_n812_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n811_), .A2(KEYINPUT113), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n370_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT113), .B1(new_n811_), .B2(new_n813_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n814_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n385_), .B(new_n395_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n386_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n819_), .A2(KEYINPUT112), .A3(new_n384_), .A4(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n384_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n385_), .A2(new_n395_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n822_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n821_), .A2(new_n826_), .A3(new_n406_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n827_), .A2(new_n372_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n805_), .B1(new_n818_), .B2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n827_), .A2(new_n372_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n811_), .A2(new_n815_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n812_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n811_), .A2(new_n813_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT58), .B(new_n830_), .C1(new_n836_), .C2(new_n814_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n829_), .A2(new_n293_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n827_), .A2(new_n374_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n407_), .A2(new_n371_), .A3(new_n409_), .ZN(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT111), .B(KEYINPUT56), .Z(new_n842_));
  NAND2_X1  g641(.A1(new_n831_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n833_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n840_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n839_), .B1(new_n845_), .B2(new_n650_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n407_), .A2(new_n371_), .A3(new_n409_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n833_), .B2(new_n843_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n774_), .B(KEYINPUT57), .C1(new_n848_), .C2(new_n840_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n838_), .A2(new_n846_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n378_), .A2(new_n740_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n691_), .A2(new_n851_), .A3(new_n347_), .A4(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n852_), .A2(new_n287_), .A3(new_n347_), .A4(new_n292_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT54), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n850_), .A2(new_n348_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n603_), .A2(new_n627_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n549_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n647_), .A2(new_n595_), .A3(new_n602_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT114), .B1(new_n861_), .B2(new_n549_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n856_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G113gat), .B1(new_n864_), .B2(new_n740_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT115), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n850_), .A2(new_n348_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n853_), .A2(new_n855_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n863_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(new_n870_), .A3(new_n873_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(KEYINPUT116), .A2(new_n872_), .B1(new_n874_), .B2(KEYINPUT59), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n872_), .A2(KEYINPUT116), .A3(KEYINPUT59), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT118), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n872_), .A2(KEYINPUT116), .A3(KEYINPUT59), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n874_), .A2(KEYINPUT59), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n873_), .B1(new_n864_), .B2(new_n871_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n878_), .B(new_n879_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n877_), .A2(new_n882_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n740_), .A2(G113gat), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n866_), .B1(new_n883_), .B2(new_n884_), .ZN(G1340gat));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n744_), .B2(G120gat), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n864_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n886_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n875_), .A2(new_n876_), .A3(new_n739_), .A4(new_n888_), .ZN(new_n890_));
  INV_X1    g689(.A(G120gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(G1341gat));
  AOI21_X1  g691(.A(G127gat), .B1(new_n864_), .B2(new_n347_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n347_), .A2(G127gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT119), .Z(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n883_), .B2(new_n895_), .ZN(G1342gat));
  INV_X1    g695(.A(G134gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n864_), .A2(new_n897_), .A3(new_n650_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n691_), .B1(new_n877_), .B2(new_n882_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1343gat));
  NOR2_X1   g699(.A1(new_n856_), .A2(new_n550_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n857_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n410_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT120), .B(G141gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1344gat));
  NOR2_X1   g704(.A1(new_n902_), .A2(new_n739_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT121), .B(G148gat), .Z(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1345gat));
  NOR2_X1   g707(.A1(new_n902_), .A2(new_n348_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT61), .B(G155gat), .Z(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  OAI21_X1  g710(.A(G162gat), .B1(new_n902_), .B2(new_n691_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n774_), .A2(G162gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n902_), .B2(new_n913_), .ZN(G1347gat));
  INV_X1    g713(.A(G169gat), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n604_), .A2(new_n647_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n858_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n915_), .B1(new_n918_), .B2(new_n740_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT123), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n856_), .A2(new_n410_), .A3(new_n917_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n922_), .B(KEYINPUT62), .C1(new_n923_), .C2(new_n915_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n920_), .A2(G169gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n923_), .B2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n918_), .A2(new_n740_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n928_), .A2(KEYINPUT122), .A3(new_n920_), .A4(G169gat), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n921_), .A2(new_n924_), .A3(new_n927_), .A4(new_n929_), .ZN(new_n930_));
  OR2_X1    g729(.A1(new_n928_), .A2(new_n494_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT124), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(new_n934_), .A3(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1348gat));
  AOI21_X1  g735(.A(G176gat), .B1(new_n918_), .B2(new_n378_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n379_), .A2(G176gat), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n918_), .B2(new_n938_), .ZN(G1349gat));
  AOI21_X1  g738(.A(new_n558_), .B1(KEYINPUT125), .B2(new_n496_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n496_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n918_), .A2(new_n347_), .ZN(new_n943_));
  MUX2_X1   g742(.A(new_n940_), .B(new_n942_), .S(new_n943_), .Z(G1350gat));
  INV_X1    g743(.A(new_n918_), .ZN(new_n945_));
  OAI21_X1  g744(.A(G190gat), .B1(new_n945_), .B2(new_n691_), .ZN(new_n946_));
  OR2_X1    g745(.A1(new_n774_), .A2(new_n559_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n945_), .B2(new_n947_), .ZN(G1351gat));
  NAND2_X1  g747(.A1(new_n901_), .A2(new_n916_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(new_n410_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(KEYINPUT126), .B(G197gat), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1352gat));
  NOR2_X1   g751(.A1(new_n949_), .A2(new_n739_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n954_), .B2(new_n448_), .ZN(new_n955_));
  XOR2_X1   g754(.A(KEYINPUT127), .B(G204gat), .Z(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n953_), .B2(new_n956_), .ZN(G1353gat));
  NOR2_X1   g756(.A1(new_n949_), .A2(new_n348_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  AND2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n958_), .B1(new_n959_), .B2(new_n960_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n961_), .B1(new_n958_), .B2(new_n959_), .ZN(G1354gat));
  OAI21_X1  g761(.A(G218gat), .B1(new_n949_), .B2(new_n691_), .ZN(new_n963_));
  OR2_X1    g762(.A1(new_n774_), .A2(G218gat), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n963_), .B1(new_n949_), .B2(new_n964_), .ZN(G1355gat));
endmodule


