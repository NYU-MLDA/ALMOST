//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT85), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT3), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(G141gat), .B2(G148gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n203_), .B1(new_n209_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n206_), .A2(new_n208_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n216_), .A2(KEYINPUT85), .A3(new_n212_), .A4(new_n213_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT86), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT86), .ZN(new_n222_));
  OR2_X1    g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n222_), .B1(new_n223_), .B2(new_n218_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n215_), .A2(new_n217_), .A3(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G141gat), .A2(G148gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT84), .B1(new_n218_), .B2(KEYINPUT1), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(KEYINPUT1), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n223_), .A3(new_n230_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n218_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n228_), .B(new_n210_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n202_), .B1(new_n226_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G197gat), .B(G204gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT21), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n235_), .A2(KEYINPUT89), .A3(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n236_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n238_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(G228gat), .B(G233gat), .C1(new_n234_), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n225_), .A2(new_n217_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n214_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT85), .B1(new_n245_), .B2(new_n216_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n233_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT87), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n226_), .A2(KEYINPUT87), .A3(new_n233_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(new_n202_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n253_));
  INV_X1    g052(.A(G228gat), .ZN(new_n254_));
  INV_X1    g053(.A(G233gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n243_), .B1(new_n252_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n243_), .B(new_n260_), .C1(new_n252_), .C2(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G22gat), .B(G50gat), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n265_), .B1(new_n251_), .B2(new_n202_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n265_), .ZN(new_n267_));
  AOI211_X1 g066(.A(KEYINPUT29), .B(new_n267_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n264_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n250_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT87), .B1(new_n226_), .B2(new_n233_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n202_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n267_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n251_), .A2(new_n202_), .A3(new_n265_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n263_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n261_), .A2(KEYINPUT90), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT91), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n262_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n277_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT91), .ZN(new_n283_));
  INV_X1    g082(.A(new_n262_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G225gat), .A2(G233gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G113gat), .B(G120gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n249_), .A2(new_n294_), .A3(new_n250_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n226_), .A2(new_n233_), .A3(new_n292_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n289_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(KEYINPUT4), .A3(new_n296_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT97), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n295_), .A2(KEYINPUT97), .A3(KEYINPUT4), .A4(new_n296_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n302_));
  AND4_X1   g101(.A1(new_n302_), .A2(new_n249_), .A3(new_n250_), .A4(new_n294_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n297_), .B1(new_n305_), .B2(new_n289_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G1gat), .B(G29gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G85gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT0), .B(G57gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n308_), .B(new_n309_), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n303_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n288_), .B1(new_n313_), .B2(new_n301_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n310_), .B1(new_n314_), .B2(new_n297_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G8gat), .B(G36gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G64gat), .B(G92gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT19), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G169gat), .ZN(new_n326_));
  INV_X1    g125(.A(G176gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n328_), .A2(KEYINPUT24), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT23), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G183gat), .A3(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n328_), .A2(KEYINPUT24), .A3(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n329_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(G190gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT25), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT79), .B1(new_n340_), .B2(G183gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT25), .B(G183gat), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n339_), .B(new_n341_), .C1(new_n342_), .C2(KEYINPUT79), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n343_), .A2(KEYINPUT80), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(KEYINPUT80), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n338_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n331_), .A2(new_n333_), .A3(KEYINPUT81), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n330_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n348_));
  INV_X1    g147(.A(G183gat), .ZN(new_n349_));
  INV_X1    g148(.A(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n348_), .A3(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G169gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n346_), .A2(new_n242_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT20), .ZN(new_n357_));
  NOR2_X1   g156(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n359_), .A2(new_n326_), .A3(new_n327_), .A4(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n360_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n328_), .B(new_n335_), .C1(new_n362_), .C2(new_n358_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n347_), .A2(new_n348_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT93), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n342_), .A2(new_n339_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n363_), .A3(new_n361_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT93), .B1(new_n370_), .B2(new_n365_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n353_), .B(new_n326_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n331_), .A2(new_n333_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT94), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n334_), .A2(new_n351_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT94), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n354_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n369_), .A2(new_n371_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT95), .B1(new_n379_), .B2(new_n253_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n357_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n253_), .A3(KEYINPUT95), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n325_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n379_), .A2(new_n253_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n242_), .B1(new_n346_), .B2(new_n355_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n325_), .A2(KEYINPUT20), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n322_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n389_));
  INV_X1    g188(.A(new_n355_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n343_), .A2(KEYINPUT80), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n343_), .A2(KEYINPUT80), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n393_), .B2(new_n338_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n389_), .B1(new_n394_), .B2(new_n242_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n379_), .A2(new_n253_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT95), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n395_), .A2(new_n398_), .A3(new_n382_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n387_), .B1(new_n399_), .B2(new_n324_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n322_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n388_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT27), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n375_), .A2(new_n354_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n370_), .B2(new_n365_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT99), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(KEYINPUT99), .B(new_n405_), .C1(new_n370_), .C2(new_n365_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n242_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT20), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT100), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n385_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(KEYINPUT100), .A3(KEYINPUT20), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n325_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  AND4_X1   g214(.A1(new_n325_), .A2(new_n395_), .A3(new_n398_), .A4(new_n382_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n322_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n404_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n403_), .A2(new_n404_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n287_), .A2(new_n317_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n401_), .A2(KEYINPUT32), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n400_), .A2(new_n421_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n300_), .A2(new_n288_), .A3(new_n301_), .A4(new_n304_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n295_), .A2(new_n289_), .A3(new_n296_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n428_), .A2(new_n311_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n402_), .A3(new_n388_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n306_), .A2(new_n311_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n431_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n315_), .A2(new_n433_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n426_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n420_), .B1(new_n437_), .B2(new_n287_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n394_), .A2(KEYINPUT30), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n346_), .A2(new_n355_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT30), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n439_), .A2(new_n442_), .A3(KEYINPUT82), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447_));
  INV_X1    g246(.A(G43gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(G15gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n449_), .B(new_n452_), .Z(new_n453_));
  NAND3_X1  g252(.A1(new_n445_), .A2(new_n446_), .A3(new_n453_), .ZN(new_n454_));
  OR3_X1    g253(.A1(new_n443_), .A2(new_n444_), .A3(new_n453_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n294_), .B(KEYINPUT31), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n454_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n317_), .A2(new_n461_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n419_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT101), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n281_), .A2(new_n286_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT101), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n461_), .A2(new_n312_), .A3(new_n315_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n419_), .A4(new_n468_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n438_), .A2(new_n462_), .B1(new_n465_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G15gat), .B(G22gat), .ZN(new_n471_));
  INV_X1    g270(.A(G1gat), .ZN(new_n472_));
  INV_X1    g271(.A(G8gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT14), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G1gat), .B(G8gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G29gat), .B(G36gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G43gat), .B(G50gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n477_), .B(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G229gat), .A2(G233gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n480_), .B(KEYINPUT15), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n477_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT77), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT77), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n487_), .A3(new_n477_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n477_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n480_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n482_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n483_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G113gat), .B(G141gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G169gat), .B(G197gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT78), .ZN(new_n499_));
  INV_X1    g298(.A(new_n497_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n492_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(new_n483_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT78), .B(new_n500_), .C1(new_n501_), .C2(new_n483_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n470_), .A2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(G85gat), .ZN(new_n510_));
  INV_X1    g309(.A(G92gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(KEYINPUT9), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT10), .B(G99gat), .ZN(new_n515_));
  OAI221_X1 g314(.A(new_n514_), .B1(KEYINPUT9), .B2(new_n513_), .C1(new_n515_), .C2(G106gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT6), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(G99gat), .A3(G106gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n520_), .A3(KEYINPUT64), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT64), .B1(new_n518_), .B2(new_n520_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n516_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n525_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n518_), .A2(new_n520_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n531_));
  INV_X1    g330(.A(G99gat), .ZN(new_n532_));
  INV_X1    g331(.A(G106gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(KEYINPUT66), .A3(new_n526_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n529_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n512_), .A2(new_n513_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT8), .ZN(new_n540_));
  INV_X1    g339(.A(new_n523_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n526_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n543_), .A3(new_n521_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT8), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n545_), .A2(KEYINPUT65), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(KEYINPUT65), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n537_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n524_), .B1(new_n540_), .B2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G57gat), .B(G64gat), .Z(new_n551_));
  INV_X1    g350(.A(KEYINPUT11), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT67), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n552_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G71gat), .B(G78gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(G57gat), .B(G64gat), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(KEYINPUT11), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .A4(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n555_), .B1(KEYINPUT11), .B2(new_n556_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n556_), .A2(new_n557_), .A3(KEYINPUT11), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n557_), .B1(new_n556_), .B2(KEYINPUT11), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n509_), .B1(new_n550_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n542_), .A2(new_n525_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n537_), .B1(new_n567_), .B2(new_n535_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n549_), .B1(new_n568_), .B2(new_n545_), .ZN(new_n569_));
  OR3_X1    g368(.A1(new_n516_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n564_), .A3(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n559_), .A2(new_n563_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n539_), .A2(KEYINPUT8), .B1(new_n544_), .B2(new_n548_), .ZN(new_n573_));
  OAI211_X1 g372(.A(KEYINPUT12), .B(new_n572_), .C1(new_n573_), .C2(new_n524_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n565_), .A2(new_n566_), .A3(new_n571_), .A4(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n566_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n571_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n564_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G120gat), .B(G148gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n575_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT71), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT71), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n575_), .A2(new_n579_), .A3(new_n587_), .A4(new_n584_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT70), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n575_), .A2(new_n579_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n584_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  AOI211_X1 g392(.A(KEYINPUT70), .B(new_n584_), .C1(new_n575_), .C2(new_n579_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n589_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n589_), .B(KEYINPUT13), .C1(new_n593_), .C2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n599_), .A2(new_n600_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n550_), .A2(new_n480_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n484_), .B1(new_n573_), .B2(new_n524_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT34), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT35), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(KEYINPUT35), .A3(new_n608_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(KEYINPUT35), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n605_), .A2(new_n606_), .A3(new_n612_), .A4(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT75), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT73), .B(KEYINPUT74), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n614_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n622_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n616_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n614_), .B(new_n615_), .C1(new_n627_), .C2(new_n623_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT37), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n626_), .A2(KEYINPUT37), .A3(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n477_), .B(KEYINPUT76), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(new_n572_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n572_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G127gat), .B(G155gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT16), .ZN(new_n641_));
  XOR2_X1   g440(.A(G183gat), .B(G211gat), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT17), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n643_), .A2(new_n644_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n639_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  OAI22_X1  g446(.A1(new_n637_), .A2(new_n638_), .B1(new_n644_), .B2(new_n643_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n633_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n604_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n507_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n472_), .A3(new_n316_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT38), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n470_), .A2(new_n629_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n649_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n599_), .A2(new_n506_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n317_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n653_), .A2(new_n654_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n655_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n655_), .A2(KEYINPUT102), .A3(new_n660_), .A4(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1324gat));
  XNOR2_X1  g465(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n667_));
  INV_X1    g466(.A(new_n419_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n656_), .A2(new_n668_), .A3(new_n658_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n473_), .B1(KEYINPUT104), .B2(KEYINPUT39), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n669_), .B(new_n670_), .C1(KEYINPUT104), .C2(KEYINPUT39), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n507_), .A2(new_n651_), .A3(new_n473_), .A4(new_n668_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT103), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n667_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  AND4_X1   g477(.A1(new_n677_), .A2(new_n674_), .A3(new_n673_), .A4(new_n667_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1325gat));
  OAI21_X1  g479(.A(G15gat), .B1(new_n659_), .B2(new_n462_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT41), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n652_), .A2(new_n451_), .A3(new_n461_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1326gat));
  XNOR2_X1  g483(.A(new_n287_), .B(KEYINPUT106), .ZN(new_n685_));
  OAI21_X1  g484(.A(G22gat), .B1(new_n659_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT42), .ZN(new_n687_));
  INV_X1    g486(.A(G22gat), .ZN(new_n688_));
  INV_X1    g487(.A(new_n685_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n652_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(G1327gat));
  INV_X1    g490(.A(new_n629_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n599_), .A2(new_n649_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n507_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n316_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n633_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT107), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT43), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n700_), .B1(new_n470_), .B2(new_n633_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n465_), .A2(new_n469_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n310_), .B(new_n434_), .C1(new_n314_), .C2(new_n297_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n403_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n436_), .A2(new_n703_), .A3(new_n704_), .A4(new_n430_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n425_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n316_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n466_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n461_), .B1(new_n709_), .B2(new_n420_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n697_), .B(new_n699_), .C1(new_n702_), .C2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n701_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n599_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n505_), .A3(new_n657_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT44), .B1(new_n712_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717_));
  AOI211_X1 g516(.A(new_n717_), .B(new_n714_), .C1(new_n701_), .C2(new_n711_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n316_), .A2(G29gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n696_), .B1(new_n719_), .B2(new_n720_), .ZN(G1328gat));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  INV_X1    g521(.A(G36gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n719_), .B2(new_n668_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n507_), .A2(new_n723_), .A3(new_n668_), .A4(new_n693_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT45), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n722_), .B1(new_n724_), .B2(new_n727_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n716_), .A2(new_n718_), .A3(new_n419_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT46), .B(new_n726_), .C1(new_n729_), .C2(new_n723_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1329gat));
  NOR4_X1   g530(.A1(new_n716_), .A2(new_n718_), .A3(new_n448_), .A4(new_n462_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G43gat), .B1(new_n695_), .B2(new_n461_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT47), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n462_), .A2(new_n448_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n719_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n734_), .A2(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n695_), .B2(new_n689_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n287_), .A2(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n719_), .B2(new_n741_), .ZN(G1331gat));
  NOR2_X1   g541(.A1(new_n470_), .A2(new_n505_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n650_), .A2(new_n713_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G57gat), .B1(new_n746_), .B2(new_n316_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n647_), .A2(new_n648_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n604_), .A2(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n656_), .A2(G57gat), .A3(new_n316_), .A4(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n750_), .A2(new_n751_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n747_), .A2(new_n752_), .A3(new_n753_), .ZN(G1332gat));
  NAND2_X1  g553(.A1(new_n656_), .A2(new_n749_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G64gat), .B1(new_n755_), .B2(new_n419_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT48), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n419_), .A2(G64gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n745_), .B2(new_n758_), .ZN(G1333gat));
  OR3_X1    g558(.A1(new_n745_), .A2(G71gat), .A3(new_n462_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G71gat), .B1(new_n755_), .B2(new_n462_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(KEYINPUT49), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(KEYINPUT49), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n760_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT109), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n766_), .B(new_n760_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1334gat));
  OAI21_X1  g567(.A(G78gat), .B1(new_n755_), .B2(new_n685_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT50), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n685_), .A2(G78gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n745_), .B2(new_n771_), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n692_), .A2(new_n649_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n743_), .A2(new_n604_), .A3(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n510_), .A3(new_n316_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n599_), .A2(new_n506_), .A3(new_n657_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n712_), .A2(KEYINPUT110), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n701_), .A2(new_n778_), .A3(new_n711_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n776_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(new_n316_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n775_), .B1(new_n781_), .B2(new_n510_), .ZN(G1336gat));
  NAND3_X1  g581(.A1(new_n774_), .A2(new_n511_), .A3(new_n668_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n780_), .A2(new_n668_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n511_), .ZN(G1337gat));
  AOI21_X1  g584(.A(new_n532_), .B1(new_n780_), .B2(new_n461_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n462_), .A2(new_n515_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n743_), .A2(new_n604_), .A3(new_n773_), .A4(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT111), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT112), .B(KEYINPUT51), .C1(new_n786_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n462_), .B(new_n776_), .C1(new_n777_), .C2(new_n779_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n792_), .B(new_n789_), .C1(new_n793_), .C2(new_n532_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n774_), .A2(new_n533_), .A3(new_n287_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n776_), .A2(new_n466_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n712_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n799_), .B2(G106gat), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT52), .B(new_n533_), .C1(new_n712_), .C2(new_n798_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n796_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g602(.A(new_n464_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n317_), .A2(new_n462_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n574_), .B(new_n571_), .C1(new_n578_), .C2(new_n508_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n576_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT55), .A3(new_n575_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n565_), .A2(new_n571_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n566_), .A4(new_n574_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n812_), .A2(KEYINPUT114), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT114), .B1(new_n812_), .B2(new_n815_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n584_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n809_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n812_), .A2(new_n815_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n584_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n812_), .A2(new_n815_), .A3(KEYINPUT114), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n819_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT56), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n589_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n820_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n482_), .B1(new_n490_), .B2(new_n480_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n482_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n500_), .B1(new_n481_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n489_), .A2(new_n829_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n832_), .B2(new_n831_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n595_), .A2(new_n498_), .A3(new_n834_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n808_), .B(new_n629_), .C1(new_n828_), .C2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n827_), .B1(new_n825_), .B2(KEYINPUT56), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n818_), .A2(new_n819_), .A3(new_n809_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n835_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT57), .B1(new_n839_), .B2(new_n692_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n836_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n834_), .A2(new_n498_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n809_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n809_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n818_), .B2(new_n847_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n823_), .A2(new_n824_), .A3(new_n847_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n843_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  OAI221_X1 g652(.A(new_n843_), .B1(new_n851_), .B2(KEYINPUT58), .C1(new_n848_), .C2(new_n849_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n697_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n649_), .B1(new_n841_), .B2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n597_), .A2(new_n748_), .A3(new_n598_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n597_), .A2(new_n748_), .A3(KEYINPUT113), .A4(new_n598_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n633_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT54), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n858_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n633_), .A4(new_n860_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n862_), .A2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT59), .B(new_n807_), .C1(new_n856_), .C2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  INV_X1    g667(.A(new_n835_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n505_), .A2(new_n589_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n821_), .A2(new_n822_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n592_), .A3(new_n824_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT115), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n870_), .B1(new_n873_), .B2(new_n809_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n869_), .B1(new_n874_), .B2(new_n826_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n808_), .B1(new_n875_), .B2(new_n629_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n839_), .A2(KEYINPUT57), .A3(new_n692_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n855_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n866_), .B1(new_n878_), .B2(new_n657_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n868_), .B1(new_n879_), .B2(new_n806_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n506_), .B1(new_n867_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(G113gat), .ZN(new_n882_));
  INV_X1    g681(.A(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n807_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n505_), .A2(new_n882_), .ZN(new_n885_));
  OAI22_X1  g684(.A1(new_n881_), .A2(new_n882_), .B1(new_n884_), .B2(new_n885_), .ZN(G1340gat));
  NOR2_X1   g685(.A1(new_n879_), .A2(new_n806_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n888_));
  AOI21_X1  g687(.A(G120gat), .B1(new_n599_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT119), .B1(new_n888_), .B2(G120gat), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n887_), .B(new_n891_), .C1(new_n889_), .C2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n604_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n867_), .B2(new_n880_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896_));
  OAI21_X1  g695(.A(G120gat), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  AOI211_X1 g696(.A(KEYINPUT120), .B(new_n894_), .C1(new_n867_), .C2(new_n880_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n893_), .B1(new_n897_), .B2(new_n898_), .ZN(G1341gat));
  INV_X1    g698(.A(G127gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n887_), .A2(new_n900_), .A3(new_n649_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n657_), .B1(new_n867_), .B2(new_n880_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n900_), .ZN(G1342gat));
  AOI21_X1  g702(.A(G134gat), .B1(new_n887_), .B2(new_n629_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n867_), .A2(new_n880_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT121), .B(G134gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n633_), .A2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n904_), .B1(new_n905_), .B2(new_n907_), .ZN(G1343gat));
  NAND4_X1  g707(.A1(new_n287_), .A2(new_n316_), .A3(new_n419_), .A4(new_n462_), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n909_), .B(KEYINPUT122), .Z(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n879_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n505_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n604_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g715(.A(KEYINPUT61), .B(G155gat), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n912_), .A2(new_n919_), .A3(new_n649_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n912_), .B2(new_n649_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n918_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n922_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n924_), .A2(new_n920_), .A3(new_n917_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1346gat));
  INV_X1    g725(.A(new_n912_), .ZN(new_n927_));
  OR3_X1    g726(.A1(new_n927_), .A2(G162gat), .A3(new_n692_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G162gat), .B1(new_n927_), .B2(new_n633_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n463_), .A2(new_n419_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n685_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n879_), .A2(new_n932_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT22), .B(G169gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(new_n505_), .A3(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n931_), .A2(new_n505_), .ZN(new_n936_));
  XOR2_X1   g735(.A(new_n936_), .B(KEYINPUT124), .Z(new_n937_));
  NAND3_X1  g736(.A1(new_n883_), .A2(new_n685_), .A3(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(KEYINPUT62), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n326_), .B1(new_n939_), .B2(KEYINPUT62), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n938_), .A2(new_n940_), .A3(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n940_), .B1(new_n938_), .B2(new_n941_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n935_), .B1(new_n943_), .B2(new_n944_), .ZN(G1348gat));
  NOR2_X1   g744(.A1(new_n879_), .A2(new_n287_), .ZN(new_n946_));
  AND4_X1   g745(.A1(G176gat), .A2(new_n946_), .A3(new_n604_), .A4(new_n931_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n879_), .A2(new_n713_), .A3(new_n932_), .ZN(new_n948_));
  OR3_X1    g747(.A1(new_n948_), .A2(KEYINPUT126), .A3(G176gat), .ZN(new_n949_));
  OAI21_X1  g748(.A(KEYINPUT126), .B1(new_n948_), .B2(G176gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n947_), .B1(new_n949_), .B2(new_n950_), .ZN(G1349gat));
  NAND3_X1  g750(.A1(new_n946_), .A2(new_n649_), .A3(new_n931_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n657_), .A2(new_n342_), .ZN(new_n953_));
  AOI22_X1  g752(.A1(new_n952_), .A2(new_n349_), .B1(new_n933_), .B2(new_n953_), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n933_), .A2(new_n339_), .A3(new_n629_), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n879_), .A2(new_n633_), .A3(new_n932_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n350_), .B2(new_n956_), .ZN(G1351gat));
  NOR4_X1   g756(.A1(new_n466_), .A2(new_n316_), .A3(new_n419_), .A4(new_n461_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n879_), .A2(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n505_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g761(.A1(new_n960_), .A2(new_n604_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g763(.A1(new_n879_), .A2(new_n657_), .A3(new_n959_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  OR3_X1    g766(.A1(new_n965_), .A2(KEYINPUT127), .A3(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(KEYINPUT127), .B1(new_n965_), .B2(new_n967_), .ZN(new_n969_));
  XOR2_X1   g768(.A(KEYINPUT63), .B(G211gat), .Z(new_n970_));
  AOI22_X1  g769(.A1(new_n968_), .A2(new_n969_), .B1(new_n965_), .B2(new_n970_), .ZN(G1354gat));
  INV_X1    g770(.A(G218gat), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n960_), .A2(new_n972_), .A3(new_n629_), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n879_), .A2(new_n633_), .A3(new_n959_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n973_), .B1(new_n972_), .B2(new_n974_), .ZN(G1355gat));
endmodule


