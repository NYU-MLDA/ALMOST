//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G231gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G57gat), .B(G64gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n213_));
  XOR2_X1   g012(.A(G71gat), .B(G78gat), .Z(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n214_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n211_), .B(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G127gat), .B(G155gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G183gat), .B(G211gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n226_));
  INV_X1    g025(.A(new_n224_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n220_), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n226_), .B1(new_n225_), .B2(new_n228_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n202_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n219_), .A2(new_n202_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n229_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G99gat), .A2(G106gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT6), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(G99gat), .A3(G106gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT65), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(new_n245_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT7), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n247_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G85gat), .B(G92gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n254_), .A2(KEYINPUT8), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n248_), .A2(KEYINPUT66), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n257_), .A2(new_n252_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n246_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n254_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT8), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n256_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT9), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(G85gat), .A3(G92gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(new_n254_), .B2(new_n265_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT64), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT10), .B(G99gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G106gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n247_), .A2(new_n272_), .A3(new_n250_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n264_), .B1(new_n268_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n267_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n273_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(KEYINPUT67), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n263_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G29gat), .B(G36gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G43gat), .B(G50gat), .Z(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT15), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n260_), .A2(new_n252_), .A3(new_n257_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT8), .B1(new_n286_), .B2(new_n254_), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n287_), .A2(new_n256_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n283_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n241_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT35), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n285_), .A2(KEYINPUT72), .A3(new_n289_), .A4(new_n240_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n292_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G190gat), .B(G218gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G134gat), .B(G162gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT36), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n299_), .B(KEYINPUT36), .Z(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  OAI22_X1  g103(.A1(new_n301_), .A2(new_n302_), .B1(new_n296_), .B2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT73), .B1(new_n296_), .B2(new_n300_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT37), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n304_), .B1(new_n296_), .B2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(new_n308_), .B2(new_n296_), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT75), .B(KEYINPUT37), .Z(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n301_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n237_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT78), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT12), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(new_n288_), .B2(new_n218_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n218_), .A2(new_n316_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n279_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G230gat), .A2(G233gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n276_), .A2(new_n277_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n263_), .A2(new_n322_), .A3(new_n218_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n317_), .A2(new_n320_), .A3(new_n321_), .A4(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n321_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n288_), .A2(new_n218_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n323_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G120gat), .B(G148gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT5), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G176gat), .B(G204gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n324_), .A2(new_n328_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT69), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n324_), .A2(new_n328_), .A3(KEYINPUT69), .A4(new_n333_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n324_), .A2(new_n328_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT68), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n324_), .A2(new_n328_), .A3(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n332_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT70), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n338_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n344_), .B1(new_n338_), .B2(new_n343_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT13), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n338_), .A2(new_n343_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT70), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT13), .B1(new_n351_), .B2(new_n345_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n315_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n348_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(KEYINPUT13), .A3(new_n345_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(KEYINPUT71), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n314_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT79), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n314_), .A2(new_n358_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G183gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT25), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G183gat), .ZN(new_n366_));
  INV_X1    g165(.A(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT26), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT26), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G190gat), .ZN(new_n370_));
  AND4_X1   g169(.A1(new_n364_), .A2(new_n366_), .A3(new_n368_), .A4(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT82), .ZN(new_n372_));
  INV_X1    g171(.A(G169gat), .ZN(new_n373_));
  INV_X1    g172(.A(G176gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT24), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT23), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n375_), .A2(KEYINPUT24), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n379_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n372_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G169gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n363_), .A2(new_n367_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n382_), .A2(new_n383_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G71gat), .B(G99gat), .ZN(new_n394_));
  INV_X1    g193(.A(G43gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n372_), .A2(new_n386_), .B1(new_n391_), .B2(new_n389_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n396_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G127gat), .B(G134gat), .Z(new_n402_));
  XOR2_X1   g201(.A(G113gat), .B(G120gat), .Z(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n401_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  INV_X1    g205(.A(G15gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT30), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT31), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n405_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n405_), .A2(new_n410_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G85gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT0), .B(G57gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT86), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G155gat), .ZN(new_n421_));
  INV_X1    g220(.A(G162gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n420_), .A2(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G141gat), .A2(G148gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT2), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT85), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n429_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n427_), .B1(new_n430_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n436_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n431_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT1), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(G155gat), .A3(G162gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n423_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT84), .B1(new_n425_), .B2(KEYINPUT1), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n425_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n442_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT87), .B1(new_n440_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n430_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n433_), .B(new_n434_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n420_), .B(new_n426_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n418_), .B2(new_n443_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n455_), .A2(new_n448_), .A3(new_n423_), .A4(new_n444_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(new_n431_), .A3(new_n441_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT87), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n450_), .A2(new_n459_), .A3(new_n404_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n404_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n440_), .A2(new_n449_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(KEYINPUT4), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT100), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G225gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n450_), .A2(new_n459_), .A3(new_n468_), .A4(new_n404_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .A4(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n460_), .A2(new_n463_), .A3(new_n466_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n467_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n465_), .B1(new_n474_), .B2(new_n464_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n417_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n464_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT100), .B1(new_n477_), .B2(new_n473_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n417_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n471_), .A4(new_n470_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n413_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n483_));
  INV_X1    g282(.A(G197gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT89), .B1(new_n484_), .B2(G204gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT89), .ZN(new_n486_));
  INV_X1    g285(.A(G204gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(G197gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(G204gat), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT21), .ZN(new_n495_));
  INV_X1    g294(.A(G218gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G211gat), .ZN(new_n497_));
  INV_X1    g296(.A(G211gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G218gat), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n494_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n493_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n483_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n489_), .A2(new_n492_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT91), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n505_), .A2(KEYINPUT92), .A3(new_n494_), .A4(new_n500_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n497_), .A2(new_n499_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n490_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n495_), .B1(G197gat), .B2(G204gat), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n489_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT90), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n511_), .A2(new_n512_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n507_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n377_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT96), .B1(new_n520_), .B2(new_n371_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT25), .B(G183gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT26), .B(G190gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT96), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n524_), .B(new_n525_), .C1(new_n377_), .C2(new_n519_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n521_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n375_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n384_), .B1(new_n528_), .B2(new_n519_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT97), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n391_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n391_), .A2(new_n531_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n389_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT98), .B1(new_n518_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT20), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n518_), .B2(new_n393_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G226gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT19), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n503_), .A2(new_n506_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT98), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n530_), .A4(new_n534_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n536_), .A2(new_n538_), .A3(new_n541_), .A4(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT99), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n537_), .B1(new_n542_), .B2(new_n398_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n518_), .A2(new_n535_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n540_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT20), .B1(new_n542_), .B2(new_n398_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(new_n540_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT99), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n536_), .A4(new_n544_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n546_), .A2(new_n550_), .A3(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G8gat), .B(G36gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT18), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G64gat), .B(G92gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n546_), .A2(new_n554_), .A3(new_n559_), .A4(new_n550_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT27), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n547_), .A2(new_n548_), .A3(new_n541_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT102), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT101), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n530_), .A2(new_n566_), .A3(new_n534_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n529_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n521_), .B2(new_n526_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n534_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT101), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n567_), .A2(new_n571_), .A3(new_n542_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n540_), .B1(new_n572_), .B2(new_n551_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT102), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n547_), .A2(new_n548_), .A3(new_n574_), .A4(new_n541_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n565_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n560_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n577_), .A2(new_n562_), .A3(KEYINPUT27), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n563_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G78gat), .B(G106gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(KEYINPUT93), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G22gat), .B(G50gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n450_), .A2(new_n459_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT28), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT29), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n586_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n584_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n590_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n584_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n588_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n583_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G228gat), .A2(G233gat), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n518_), .B(new_n597_), .C1(new_n585_), .C2(new_n587_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n462_), .A2(new_n587_), .ZN(new_n599_));
  OAI211_X1 g398(.A(G228gat), .B(G233gat), .C1(new_n542_), .C2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT94), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n598_), .A2(new_n603_), .A3(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n591_), .A2(new_n594_), .A3(new_n581_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n596_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n602_), .A2(new_n604_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n606_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n595_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n482_), .A2(new_n579_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n559_), .A2(KEYINPUT32), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n576_), .A2(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n546_), .A2(new_n554_), .A3(new_n550_), .A4(new_n613_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n481_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT103), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n481_), .A2(new_n615_), .A3(new_n616_), .A4(new_n619_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n460_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n469_), .A2(new_n466_), .ZN(new_n622_));
  AOI211_X1 g421(.A(new_n479_), .B(new_n621_), .C1(new_n464_), .C2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n480_), .B2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n472_), .A2(new_n475_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(KEYINPUT33), .A3(new_n479_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n561_), .A2(new_n625_), .A3(new_n562_), .A4(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n618_), .A2(new_n620_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n611_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n611_), .A2(new_n481_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n579_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n411_), .A2(new_n412_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT83), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n612_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n283_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(new_n209_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G229gat), .A2(G233gat), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n284_), .A2(new_n209_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n637_), .B(new_n209_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n639_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n640_), .A2(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G113gat), .B(G141gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G169gat), .B(G197gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n644_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n636_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n481_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(G1gat), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n360_), .A2(new_n362_), .A3(new_n652_), .A4(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT38), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n655_), .A2(KEYINPUT104), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT104), .B1(new_n655_), .B2(new_n656_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n310_), .A2(new_n301_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n636_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n662_), .A2(new_n358_), .A3(new_n650_), .A4(new_n236_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n663_), .A2(new_n653_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G1gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n665_), .B1(new_n656_), .B2(new_n655_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT105), .B1(new_n659_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n655_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n668_), .A2(KEYINPUT38), .B1(new_n664_), .B2(G1gat), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n669_), .B(new_n670_), .C1(new_n658_), .C2(new_n657_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n667_), .A2(new_n671_), .ZN(G1324gat));
  NOR2_X1   g471(.A1(new_n663_), .A2(new_n579_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT106), .B1(new_n673_), .B2(new_n205_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n360_), .A2(new_n652_), .A3(new_n362_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n579_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n205_), .ZN(new_n677_));
  OAI22_X1  g476(.A1(new_n674_), .A2(KEYINPUT39), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n663_), .A2(new_n579_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(new_n681_), .A3(G8gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(KEYINPUT39), .A3(new_n674_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n679_), .A2(KEYINPUT40), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n682_), .A2(KEYINPUT39), .A3(new_n674_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(new_n678_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(G1325gat));
  OAI21_X1  g487(.A(G15gat), .B1(new_n663_), .B2(new_n635_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT41), .Z(new_n690_));
  INV_X1    g489(.A(new_n635_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n407_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n675_), .B2(new_n692_), .ZN(G1326gat));
  OAI21_X1  g492(.A(G22gat), .B1(new_n663_), .B2(new_n611_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT42), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n611_), .A2(G22gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n675_), .B2(new_n696_), .ZN(G1327gat));
  NAND2_X1  g496(.A1(new_n661_), .A2(new_n237_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n357_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n652_), .ZN(new_n700_));
  OR3_X1    g499(.A1(new_n700_), .A2(G29gat), .A3(new_n653_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n307_), .A2(new_n312_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n636_), .B2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n482_), .A2(new_n579_), .A3(new_n611_), .ZN(new_n704_));
  AOI22_X1  g503(.A1(new_n629_), .A2(new_n611_), .B1(new_n579_), .B2(new_n631_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n691_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  INV_X1    g506(.A(new_n702_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n703_), .A2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n353_), .A2(new_n650_), .A3(new_n237_), .A4(new_n356_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT44), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  AOI211_X1 g513(.A(new_n714_), .B(new_n711_), .C1(new_n703_), .C2(new_n709_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n481_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G29gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n716_), .B2(new_n481_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n701_), .B1(new_n719_), .B2(new_n720_), .ZN(G1328gat));
  NOR3_X1   g520(.A1(new_n700_), .A2(G36gat), .A3(new_n579_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n716_), .B2(new_n676_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n707_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n712_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n714_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n712_), .B(KEYINPUT44), .C1(new_n727_), .C2(new_n728_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n730_), .A2(new_n725_), .A3(new_n676_), .A4(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G36gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n724_), .B1(new_n726_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n724_), .B(KEYINPUT46), .C1(new_n726_), .C2(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1329gat));
  NAND3_X1  g537(.A1(new_n716_), .A2(G43gat), .A3(new_n634_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT109), .B(G43gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(new_n700_), .B2(new_n635_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g542(.A(G50gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n611_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n611_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n699_), .A2(new_n652_), .A3(new_n746_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n716_), .A2(new_n745_), .B1(new_n744_), .B2(new_n747_), .ZN(G1331gat));
  AND4_X1   g547(.A1(new_n651_), .A2(new_n314_), .A3(new_n706_), .A4(new_n357_), .ZN(new_n749_));
  INV_X1    g548(.A(G57gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n481_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n357_), .A2(new_n651_), .A3(new_n236_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n706_), .A2(new_n660_), .ZN(new_n754_));
  OR3_X1    g553(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n481_), .A3(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n751_), .B1(new_n757_), .B2(new_n750_), .ZN(G1332gat));
  INV_X1    g557(.A(G64gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n749_), .A2(new_n759_), .A3(new_n676_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n755_), .A2(new_n676_), .A3(new_n756_), .ZN(new_n761_));
  XOR2_X1   g560(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(G64gat), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(G64gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(G1333gat));
  NOR2_X1   g564(.A1(new_n635_), .A2(G71gat), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT112), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n749_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n755_), .A2(new_n691_), .A3(new_n756_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G71gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G71gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(G1334gat));
  INV_X1    g572(.A(G78gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n749_), .A2(new_n774_), .A3(new_n746_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n755_), .A2(new_n746_), .A3(new_n756_), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(G78gat), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G78gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n775_), .B(KEYINPUT114), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1335gat));
  OR2_X1    g583(.A1(new_n710_), .A2(KEYINPUT115), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n710_), .A2(KEYINPUT115), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n357_), .A2(new_n651_), .A3(new_n237_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n357_), .A2(KEYINPUT116), .A3(new_n651_), .A4(new_n237_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n786_), .A3(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792_), .B2(new_n653_), .ZN(new_n793_));
  NOR4_X1   g592(.A1(new_n358_), .A2(new_n650_), .A3(new_n636_), .A4(new_n698_), .ZN(new_n794_));
  INV_X1    g593(.A(G85gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n481_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n793_), .A2(new_n796_), .A3(KEYINPUT117), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1336gat));
  OAI21_X1  g600(.A(G92gat), .B1(new_n792_), .B2(new_n579_), .ZN(new_n802_));
  INV_X1    g601(.A(G92gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n794_), .A2(new_n803_), .A3(new_n676_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1337gat));
  OAI21_X1  g604(.A(G99gat), .B1(new_n792_), .B2(new_n635_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n794_), .A2(new_n634_), .A3(new_n270_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT51), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n810_), .A3(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1338gat));
  NAND3_X1  g611(.A1(new_n794_), .A2(new_n271_), .A3(new_n746_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n611_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n710_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n814_), .B1(new_n816_), .B2(G106gat), .ZN(new_n817_));
  AOI211_X1 g616(.A(KEYINPUT52), .B(new_n271_), .C1(new_n815_), .C2(new_n710_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n813_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT53), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n813_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1339gat));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT119), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n327_), .B1(new_n279_), .B2(new_n319_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n321_), .B1(new_n827_), .B2(new_n317_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n324_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n827_), .A2(KEYINPUT55), .A3(new_n321_), .A4(new_n317_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n332_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n834_), .B(new_n333_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n644_), .A2(new_n649_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n641_), .A2(new_n638_), .A3(new_n643_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n649_), .B1(new_n642_), .B2(new_n639_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n338_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n826_), .B1(new_n836_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n843_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n825_), .B(new_n845_), .C1(new_n833_), .C2(new_n835_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n708_), .A3(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n650_), .B(new_n338_), .C1(new_n833_), .C2(new_n835_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n842_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n661_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n847_), .B1(KEYINPUT57), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n338_), .A2(new_n650_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n832_), .A2(new_n332_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n834_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n332_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n854_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n841_), .B1(new_n351_), .B2(new_n345_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n660_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n853_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n850_), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n236_), .B1(new_n852_), .B2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n313_), .A2(new_n651_), .A3(new_n355_), .A4(new_n354_), .ZN(new_n866_));
  AND2_X1   g665(.A1(KEYINPUT118), .A2(KEYINPUT54), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(KEYINPUT118), .A2(KEYINPUT54), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n866_), .B1(new_n869_), .B2(new_n867_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n865_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n579_), .A2(new_n481_), .A3(new_n611_), .A4(new_n634_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n851_), .A2(new_n876_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n847_), .B(KEYINPUT121), .C1(KEYINPUT57), .C2(new_n850_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n864_), .A3(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n871_), .B1(new_n879_), .B2(new_n237_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n873_), .A2(KEYINPUT59), .ZN(new_n881_));
  OAI22_X1  g680(.A1(new_n874_), .A2(new_n875_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G113gat), .B1(new_n882_), .B2(new_n651_), .ZN(new_n883_));
  INV_X1    g682(.A(G113gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n874_), .A2(new_n884_), .A3(new_n650_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1340gat));
  OAI21_X1  g685(.A(G120gat), .B1(new_n882_), .B2(new_n358_), .ZN(new_n887_));
  INV_X1    g686(.A(G120gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n358_), .B2(KEYINPUT60), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n874_), .B(new_n889_), .C1(KEYINPUT60), .C2(new_n888_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n887_), .A2(new_n890_), .ZN(G1341gat));
  OAI21_X1  g690(.A(G127gat), .B1(new_n882_), .B2(new_n237_), .ZN(new_n892_));
  INV_X1    g691(.A(G127gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n874_), .A2(new_n893_), .A3(new_n236_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1342gat));
  OAI21_X1  g694(.A(G134gat), .B1(new_n882_), .B2(new_n702_), .ZN(new_n896_));
  INV_X1    g695(.A(G134gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n874_), .A2(new_n897_), .A3(new_n661_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1343gat));
  NAND2_X1  g698(.A1(new_n868_), .A2(new_n870_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n851_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n236_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n691_), .A2(new_n611_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n481_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n676_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n902_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n650_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g707(.A1(new_n902_), .A2(new_n357_), .A3(new_n905_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT123), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n902_), .A2(new_n911_), .A3(new_n357_), .A4(new_n905_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT122), .B(G148gat), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n910_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n910_), .B2(new_n912_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1345gat));
  NAND2_X1  g715(.A1(new_n906_), .A2(new_n236_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT61), .B(G155gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1346gat));
  NAND3_X1  g718(.A1(new_n902_), .A2(new_n708_), .A3(new_n905_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G162gat), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n902_), .A2(new_n422_), .A3(new_n661_), .A4(new_n905_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n921_), .A2(KEYINPUT124), .A3(new_n922_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n579_), .A2(new_n481_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n691_), .A2(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(KEYINPUT125), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n746_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n851_), .A2(new_n876_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n236_), .B1(new_n932_), .B2(new_n878_), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n650_), .B(new_n931_), .C1(new_n933_), .C2(new_n871_), .ZN(new_n934_));
  OAI211_X1 g733(.A(KEYINPUT62), .B(G169gat), .C1(new_n934_), .C2(KEYINPUT22), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  INV_X1    g735(.A(new_n934_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT22), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n373_), .B1(new_n937_), .B2(new_n936_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n935_), .B1(new_n939_), .B2(new_n940_), .ZN(G1348gat));
  INV_X1    g740(.A(new_n931_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n880_), .A2(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(G176gat), .B1(new_n943_), .B2(new_n357_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n872_), .A2(new_n942_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n358_), .A2(new_n374_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n944_), .B1(new_n945_), .B2(new_n946_), .ZN(G1349gat));
  AOI21_X1  g746(.A(G183gat), .B1(new_n945_), .B2(new_n236_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n237_), .A2(new_n522_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n948_), .B1(new_n943_), .B2(new_n949_), .ZN(G1350gat));
  INV_X1    g749(.A(new_n943_), .ZN(new_n951_));
  OAI21_X1  g750(.A(G190gat), .B1(new_n951_), .B2(new_n702_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n943_), .A2(new_n523_), .A3(new_n661_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1351gat));
  NAND2_X1  g753(.A1(new_n903_), .A2(new_n928_), .ZN(new_n955_));
  OAI21_X1  g754(.A(KEYINPUT126), .B1(new_n872_), .B2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957_));
  INV_X1    g756(.A(new_n955_), .ZN(new_n958_));
  OAI211_X1 g757(.A(new_n957_), .B(new_n958_), .C1(new_n865_), .C2(new_n871_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n956_), .A2(new_n959_), .ZN(new_n960_));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960_), .B2(new_n650_), .ZN(new_n961_));
  AOI211_X1 g760(.A(new_n484_), .B(new_n651_), .C1(new_n956_), .C2(new_n959_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1352gat));
  INV_X1    g762(.A(new_n959_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n957_), .B1(new_n902_), .B2(new_n958_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n357_), .B1(new_n964_), .B2(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n966_), .A2(new_n967_), .A3(G204gat), .ZN(new_n968_));
  OAI211_X1 g767(.A(new_n960_), .B(new_n357_), .C1(KEYINPUT127), .C2(new_n487_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1353gat));
  OR2_X1    g769(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n971_), .B1(new_n960_), .B2(new_n236_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(KEYINPUT63), .B(G211gat), .ZN(new_n973_));
  AOI211_X1 g772(.A(new_n237_), .B(new_n973_), .C1(new_n956_), .C2(new_n959_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n972_), .A2(new_n974_), .ZN(G1354gat));
  NAND3_X1  g774(.A1(new_n960_), .A2(new_n496_), .A3(new_n661_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n702_), .B1(new_n956_), .B2(new_n959_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n496_), .B2(new_n977_), .ZN(G1355gat));
endmodule


