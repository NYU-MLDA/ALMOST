//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  INV_X1    g000(.A(G36gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G29gat), .ZN(new_n203_));
  INV_X1    g002(.A(G29gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G36gat), .ZN(new_n205_));
  INV_X1    g004(.A(G50gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G43gat), .ZN(new_n207_));
  INV_X1    g006(.A(G43gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G50gat), .ZN(new_n209_));
  AND4_X1   g008(.A1(new_n203_), .A2(new_n205_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n203_), .A2(new_n205_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT15), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(G1gat), .B2(G8gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT71), .A2(G15gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT71), .A2(G15gat), .ZN(new_n219_));
  INV_X1    g018(.A(G22gat), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT71), .ZN(new_n222_));
  INV_X1    g021(.A(G15gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(G22gat), .B1(new_n224_), .B2(new_n217_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n216_), .B1(new_n221_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G1gat), .B(G8gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n220_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n224_), .A2(G22gat), .A3(new_n217_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n227_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n216_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n228_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n213_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n228_), .A2(new_n212_), .A3(new_n233_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G113gat), .B(G141gat), .Z(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT79), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G169gat), .B(G197gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n240_), .B(new_n241_), .Z(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n210_), .A2(new_n211_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n234_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT76), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n237_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n248_), .B1(new_n237_), .B2(new_n247_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n246_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n232_), .B1(new_n231_), .B2(new_n216_), .ZN(new_n252_));
  AOI211_X1 g051(.A(new_n215_), .B(new_n227_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n252_), .A2(new_n253_), .A3(new_n245_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT76), .B1(new_n254_), .B2(KEYINPUT75), .ZN(new_n255_));
  INV_X1    g054(.A(new_n246_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n237_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n251_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n236_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n244_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AOI211_X1 g060(.A(KEYINPUT77), .B(new_n236_), .C1(new_n251_), .C2(new_n258_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n238_), .B(new_n243_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT80), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n249_), .A2(new_n250_), .A3(new_n246_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n256_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n260_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT77), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n259_), .A2(new_n244_), .A3(new_n260_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n271_), .A2(KEYINPUT80), .A3(new_n238_), .A4(new_n243_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n265_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n238_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT78), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OAI211_X1 g075(.A(KEYINPUT78), .B(new_n238_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n242_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT81), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(KEYINPUT24), .A3(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT83), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT25), .B(G183gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT26), .B(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT23), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n289_), .B(new_n295_), .C1(KEYINPUT24), .C2(new_n286_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT22), .B(G169gat), .ZN(new_n297_));
  INV_X1    g096(.A(G176gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(KEYINPUT84), .Z(new_n300_));
  OAI21_X1  g099(.A(new_n294_), .B1(G183gat), .B2(G190gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n287_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n296_), .A2(KEYINPUT85), .A3(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G227gat), .A2(G233gat), .ZN(new_n308_));
  INV_X1    g107(.A(G71gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(G99gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n307_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n314_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G15gat), .B(G43gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT86), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT30), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G127gat), .B(G134gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G113gat), .B(G120gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n320_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n315_), .A2(new_n324_), .A3(new_n316_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G211gat), .B(G218gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(G197gat), .B(G204gat), .Z(new_n331_));
  INV_X1    g130(.A(KEYINPUT90), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G204gat), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n334_), .A2(G197gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT21), .B1(new_n335_), .B2(KEYINPUT90), .ZN(new_n336_));
  OAI221_X1 g135(.A(new_n330_), .B1(KEYINPUT21), .B2(new_n331_), .C1(new_n333_), .C2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n330_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(KEYINPUT21), .A3(new_n331_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n342_));
  NAND3_X1  g141(.A1(new_n286_), .A2(new_n287_), .A3(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n295_), .B(new_n343_), .C1(new_n286_), .C2(new_n342_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n301_), .A2(new_n287_), .A3(new_n299_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n340_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n346_), .A2(KEYINPUT93), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(KEYINPUT93), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT19), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT20), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n348_), .A3(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n341_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n305_), .A2(new_n340_), .A3(new_n306_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n340_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n344_), .A2(new_n345_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n351_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n350_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT18), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND3_X1  g163(.A1(new_n354_), .A2(new_n360_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT96), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n346_), .A2(KEYINPUT20), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n350_), .B1(new_n341_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n350_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n355_), .A2(new_n371_), .A3(new_n358_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n364_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n368_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n354_), .A2(new_n360_), .A3(KEYINPUT96), .A4(new_n364_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n367_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n341_), .A2(new_n353_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n371_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n374_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n365_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n368_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G78gat), .B(G106gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT3), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT2), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT89), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394_));
  OR2_X1    g193(.A1(G155gat), .A2(G162gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(KEYINPUT1), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n395_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n394_), .A2(KEYINPUT1), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n397_), .B(new_n389_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n401_), .B(KEYINPUT88), .Z(new_n402_));
  NAND2_X1  g201(.A1(new_n396_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT29), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n356_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(G228gat), .A3(G233gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G228gat), .A2(G233gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n356_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n386_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n408_), .A3(new_n386_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n403_), .A2(KEYINPUT29), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G22gat), .B(G50gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT28), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n413_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT91), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n416_), .B1(new_n409_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n412_), .A2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n410_), .A2(new_n417_), .A3(new_n411_), .A4(new_n416_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(G85gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT0), .B(G57gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  OR2_X1    g224(.A1(new_n403_), .A2(new_n323_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n403_), .A2(new_n323_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(KEYINPUT4), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT94), .B1(new_n427_), .B2(KEYINPUT4), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT94), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n403_), .A2(new_n432_), .A3(new_n433_), .A4(new_n323_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .A4(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n426_), .A2(new_n427_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n429_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n425_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n437_), .A3(new_n425_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n421_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n384_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT95), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n444_), .B1(new_n373_), .B2(new_n446_), .ZN(new_n447_));
  AOI211_X1 g246(.A(KEYINPUT95), .B(new_n445_), .C1(new_n370_), .C2(new_n372_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n354_), .A2(new_n360_), .A3(new_n445_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n435_), .A2(new_n425_), .A3(new_n437_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(new_n438_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n425_), .B1(new_n436_), .B2(new_n430_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n428_), .A2(new_n434_), .A3(new_n431_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n454_), .B1(new_n455_), .B2(new_n430_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n435_), .A2(new_n437_), .A3(KEYINPUT33), .A4(new_n425_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n456_), .A2(new_n365_), .A3(new_n457_), .A4(new_n380_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n451_), .A2(KEYINPUT33), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n421_), .B1(new_n453_), .B2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n329_), .B1(new_n443_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n441_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n326_), .A2(new_n463_), .A3(new_n327_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n419_), .A2(new_n420_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT97), .B1(new_n383_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT97), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n421_), .A2(new_n377_), .A3(new_n467_), .A4(new_n382_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n464_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n282_), .B1(new_n462_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT66), .ZN(new_n471_));
  INV_X1    g270(.A(G57gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(G64gat), .ZN(new_n473_));
  INV_X1    g272(.A(G64gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(G57gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n471_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT11), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(G57gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(G64gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(KEYINPUT66), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(new_n477_), .A3(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G71gat), .B(G78gat), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT67), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n476_), .A2(new_n480_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(KEYINPUT11), .ZN(new_n486_));
  AOI211_X1 g285(.A(KEYINPUT67), .B(new_n477_), .C1(new_n476_), .C2(new_n480_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n483_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n478_), .A2(new_n479_), .A3(KEYINPUT66), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT66), .B1(new_n478_), .B2(new_n479_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT11), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT67), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n485_), .A2(new_n484_), .A3(KEYINPUT11), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n252_), .A2(new_n253_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G231gat), .A2(G233gat), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT74), .B(KEYINPUT17), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n498_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G127gat), .B(G155gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G183gat), .B(G211gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n502_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n502_), .A2(new_n508_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n499_), .A2(new_n501_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT73), .B(KEYINPUT17), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G232gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT34), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT35), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n517_), .B(KEYINPUT69), .Z(new_n518_));
  NOR2_X1   g317(.A1(new_n516_), .A2(KEYINPUT35), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G85gat), .B(G92gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT6), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(G99gat), .A3(G106gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  AOI211_X1 g328(.A(KEYINPUT8), .B(new_n520_), .C1(new_n524_), .C2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT8), .ZN(new_n531_));
  INV_X1    g330(.A(new_n523_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(new_n532_), .A3(new_n521_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n520_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n531_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT65), .B(G92gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT64), .B(G85gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT9), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(G85gat), .ZN(new_n540_));
  INV_X1    g339(.A(G92gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT9), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n539_), .A2(new_n542_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT10), .B(G99gat), .Z(new_n544_));
  INV_X1    g343(.A(G106gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n529_), .ZN(new_n547_));
  OAI22_X1  g346(.A1(new_n530_), .A2(new_n535_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n519_), .B1(new_n213_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n548_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n212_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n518_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(KEYINPUT36), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n549_), .A2(new_n551_), .A3(new_n518_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n553_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT37), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(new_n558_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n556_), .B(KEYINPUT36), .Z(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT70), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n553_), .A2(KEYINPUT70), .A3(new_n558_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n562_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n559_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n563_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(G230gat), .A2(G233gat), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n495_), .B2(new_n550_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n488_), .A2(new_n548_), .A3(new_n494_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n488_), .A2(new_n548_), .A3(new_n494_), .A4(KEYINPUT12), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n495_), .A2(new_n550_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n573_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n579_), .A2(KEYINPUT68), .A3(new_n571_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT68), .B1(new_n579_), .B2(new_n571_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n577_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT5), .ZN(new_n584_));
  XOR2_X1   g383(.A(G176gat), .B(G204gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n586_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n587_), .A2(KEYINPUT13), .A3(new_n588_), .ZN(new_n592_));
  AND4_X1   g391(.A1(new_n514_), .A2(new_n570_), .A3(new_n591_), .A4(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n470_), .A2(KEYINPUT98), .A3(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT98), .B1(new_n470_), .B2(new_n594_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(G1gat), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n441_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT38), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n462_), .A2(new_n469_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n568_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n591_), .A2(new_n592_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n273_), .A2(new_n278_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT99), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(new_n514_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n603_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n598_), .B1(new_n609_), .B2(new_n441_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT100), .Z(new_n611_));
  NAND2_X1  g410(.A1(new_n600_), .A2(new_n611_), .ZN(G1324gat));
  NOR2_X1   g411(.A1(new_n384_), .A2(G8gat), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n595_), .A2(new_n596_), .A3(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT101), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n603_), .A2(new_n383_), .A3(new_n608_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n616_), .A2(G8gat), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n616_), .B2(G8gat), .ZN(new_n621_));
  OAI22_X1  g420(.A1(new_n620_), .A2(new_n621_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n615_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n615_), .B2(new_n622_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1325gat));
  NAND3_X1  g425(.A1(new_n597_), .A2(new_n223_), .A3(new_n329_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n609_), .A2(new_n329_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n628_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT41), .B1(new_n628_), .B2(G15gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n627_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT104), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n633_), .B(new_n627_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1326gat));
  AOI21_X1  g434(.A(new_n220_), .B1(new_n609_), .B2(new_n465_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT42), .Z(new_n637_));
  NAND3_X1  g436(.A1(new_n597_), .A2(new_n220_), .A3(new_n465_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1327gat));
  INV_X1    g438(.A(new_n514_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n602_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n470_), .A2(new_n604_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n441_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n607_), .A2(new_n640_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n570_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n462_), .B2(new_n469_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT43), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n648_), .B(new_n645_), .C1(new_n462_), .C2(new_n469_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n644_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(KEYINPUT44), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n649_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n644_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(KEYINPUT44), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n650_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n651_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n463_), .A2(new_n204_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n643_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  NAND3_X1  g459(.A1(new_n642_), .A2(new_n202_), .A3(new_n383_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT45), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n383_), .B1(new_n650_), .B2(KEYINPUT44), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n662_), .B1(new_n664_), .B2(new_n202_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT46), .B(new_n662_), .C1(new_n664_), .C2(new_n202_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  XNOR2_X1  g468(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n328_), .A2(new_n208_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n673_), .B(new_n651_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G43gat), .B1(new_n642_), .B2(new_n329_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n658_), .A2(new_n672_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n675_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n678_), .A3(new_n670_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1330gat));
  AOI21_X1  g479(.A(G50gat), .B1(new_n642_), .B2(new_n465_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n421_), .A2(new_n206_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n658_), .B2(new_n682_), .ZN(G1331gat));
  INV_X1    g482(.A(new_n604_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(new_n640_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n603_), .A2(new_n281_), .A3(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(G57gat), .A3(new_n441_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT108), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n601_), .A2(new_n279_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n685_), .A2(new_n570_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n472_), .B1(new_n692_), .B2(new_n463_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n694_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n688_), .A2(new_n695_), .A3(new_n696_), .ZN(G1332gat));
  AOI21_X1  g496(.A(new_n474_), .B1(new_n686_), .B2(new_n383_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT48), .Z(new_n699_));
  INV_X1    g498(.A(new_n692_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(new_n474_), .A3(new_n383_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1333gat));
  AOI21_X1  g501(.A(new_n309_), .B1(new_n686_), .B2(new_n329_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT49), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n700_), .A2(new_n309_), .A3(new_n329_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1334gat));
  INV_X1    g505(.A(G78gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n686_), .B2(new_n465_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT50), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n700_), .A2(new_n707_), .A3(new_n465_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n684_), .A2(new_n641_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n689_), .A2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n540_), .B1(new_n713_), .B2(new_n463_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT109), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n684_), .A2(new_n514_), .A3(new_n279_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n441_), .A2(new_n537_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(G1336gat));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n383_), .A3(new_n536_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n541_), .B1(new_n713_), .B2(new_n384_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1337gat));
  AND2_X1   g522(.A1(new_n718_), .A2(new_n329_), .ZN(new_n724_));
  INV_X1    g523(.A(G99gat), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n689_), .A2(new_n329_), .A3(new_n544_), .A4(new_n712_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n726_), .A2(new_n727_), .A3(KEYINPUT111), .A4(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n728_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n731_), .A2(new_n733_), .A3(new_n735_), .ZN(G1338gat));
  NAND3_X1  g535(.A1(new_n652_), .A2(new_n465_), .A3(new_n716_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT113), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n718_), .A2(new_n739_), .A3(new_n465_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n738_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n689_), .A2(new_n545_), .A3(new_n465_), .A4(new_n712_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT112), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n421_), .B(new_n717_), .C1(new_n647_), .C2(new_n649_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n545_), .B1(new_n745_), .B2(new_n739_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT52), .B1(new_n746_), .B2(new_n738_), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT53), .B1(new_n744_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n740_), .A2(G106gat), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n745_), .A2(new_n739_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n741_), .A4(new_n743_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n748_), .A2(new_n754_), .ZN(G1339gat));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n281_), .A2(new_n756_), .A3(new_n593_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n281_), .B2(new_n593_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n577_), .A2(KEYINPUT55), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n572_), .A2(new_n575_), .A3(new_n761_), .A4(new_n576_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n575_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n571_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n763_), .A2(new_n764_), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n764_), .B1(new_n763_), .B2(new_n766_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n586_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT56), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT56), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n586_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n279_), .A2(new_n587_), .A3(new_n770_), .A4(new_n772_), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n236_), .B(new_n254_), .C1(new_n213_), .C2(new_n234_), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n243_), .B(new_n774_), .C1(new_n259_), .C2(new_n236_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n265_), .B2(new_n272_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n589_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n602_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n770_), .A2(new_n776_), .A3(new_n587_), .A4(new_n772_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n570_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n772_), .A2(new_n587_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n780_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n783_), .A2(new_n776_), .A3(new_n770_), .A4(new_n784_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n778_), .A2(KEYINPUT57), .B1(new_n781_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n776_), .A2(new_n589_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n763_), .A2(new_n766_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT114), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n763_), .A2(new_n764_), .A3(new_n766_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n771_), .B1(new_n793_), .B2(new_n586_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n782_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n789_), .B1(new_n795_), .B2(new_n279_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n787_), .B(new_n788_), .C1(new_n796_), .C2(new_n602_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT115), .B1(new_n778_), .B2(KEYINPUT57), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n786_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n759_), .B1(new_n799_), .B2(new_n640_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n466_), .A2(new_n468_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(new_n441_), .A3(new_n329_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G113gat), .B1(new_n803_), .B2(new_n279_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT117), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT59), .B1(new_n800_), .B2(new_n802_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT118), .B(KEYINPUT59), .C1(new_n800_), .C2(new_n802_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n770_), .A2(new_n587_), .A3(new_n772_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n777_), .B1(new_n811_), .B2(new_n605_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT57), .A3(new_n568_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n779_), .A2(new_n780_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n785_), .A2(new_n814_), .A3(new_n645_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n778_), .A2(KEYINPUT57), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n640_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n758_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n281_), .A2(new_n756_), .A3(new_n593_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n801_), .A2(new_n823_), .A3(new_n441_), .A4(new_n329_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT119), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n822_), .A2(new_n828_), .A3(new_n825_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n810_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n282_), .A2(G113gat), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT120), .Z(new_n833_));
  AOI21_X1  g632(.A(new_n805_), .B1(new_n831_), .B2(new_n833_), .ZN(G1340gat));
  INV_X1    g633(.A(G120gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n684_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n810_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT60), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT121), .B1(new_n838_), .B2(G120gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(G120gat), .B1(new_n604_), .B2(new_n838_), .ZN(new_n840_));
  MUX2_X1   g639(.A(new_n839_), .B(KEYINPUT121), .S(new_n840_), .Z(new_n841_));
  NAND2_X1  g640(.A1(new_n803_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT122), .B1(new_n837_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n828_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n846_));
  AOI211_X1 g645(.A(KEYINPUT119), .B(new_n824_), .C1(new_n818_), .C2(new_n821_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n604_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n845_), .B(new_n842_), .C1(new_n849_), .C2(new_n835_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n844_), .A2(new_n850_), .ZN(G1341gat));
  INV_X1    g650(.A(G127gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n803_), .A2(new_n852_), .A3(new_n514_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n810_), .A2(new_n514_), .A3(new_n830_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n852_), .ZN(G1342gat));
  INV_X1    g654(.A(G134gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n803_), .A2(new_n856_), .A3(new_n602_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n810_), .A2(new_n645_), .A3(new_n830_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n856_), .ZN(G1343gat));
  INV_X1    g658(.A(new_n800_), .ZN(new_n860_));
  NOR4_X1   g659(.A1(new_n329_), .A2(new_n383_), .A3(new_n463_), .A4(new_n421_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n279_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n604_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n863_), .A2(new_n514_), .A3(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n862_), .B2(new_n640_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  AOI21_X1  g673(.A(G162gat), .B1(new_n863_), .B2(new_n602_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n645_), .A2(G162gat), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(KEYINPUT125), .Z(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n863_), .B2(new_n877_), .ZN(G1347gat));
  AOI21_X1  g677(.A(new_n465_), .B1(new_n818_), .B2(new_n821_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n384_), .A2(new_n464_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G169gat), .B1(new_n881_), .B2(new_n605_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT127), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n883_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n886_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n882_), .A2(new_n883_), .A3(new_n888_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n879_), .A2(new_n297_), .A3(new_n279_), .A4(new_n880_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n889_), .A3(new_n890_), .ZN(G1348gat));
  NAND3_X1  g690(.A1(new_n879_), .A2(new_n604_), .A3(new_n880_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n800_), .A2(new_n465_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n880_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n894_), .A2(new_n298_), .A3(new_n684_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n892_), .A2(new_n298_), .B1(new_n893_), .B2(new_n895_), .ZN(G1349gat));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n640_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G183gat), .B1(new_n893_), .B2(new_n897_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n894_), .A2(new_n290_), .A3(new_n640_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n879_), .B2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n881_), .B2(new_n570_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n602_), .A2(new_n291_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n881_), .B2(new_n902_), .ZN(G1351gat));
  AND3_X1   g702(.A1(new_n442_), .A2(new_n328_), .A3(new_n383_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n860_), .A2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n279_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g707(.A1(new_n905_), .A2(new_n684_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n334_), .ZN(G1353gat));
  NAND2_X1  g709(.A1(new_n906_), .A2(new_n514_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  AND2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n911_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n911_), .B2(new_n912_), .ZN(G1354gat));
  OR3_X1    g714(.A1(new_n905_), .A2(G218gat), .A3(new_n568_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G218gat), .B1(new_n905_), .B2(new_n570_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1355gat));
endmodule


