//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT8), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT64), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  AND2_X1   g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n206_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G85gat), .B(G92gat), .Z(new_n215_));
  AOI21_X1  g014(.A(new_n204_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n204_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n212_), .A2(new_n213_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n207_), .A2(KEYINPUT64), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT65), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n206_), .B1(new_n219_), .B2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n217_), .B1(new_n226_), .B2(KEYINPUT66), .ZN(new_n227_));
  INV_X1    g026(.A(new_n206_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n218_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n223_), .A2(KEYINPUT65), .A3(new_n224_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n216_), .B1(new_n227_), .B2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n219_), .A2(new_n225_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT10), .B(G99gat), .ZN(new_n238_));
  OAI221_X1 g037(.A(new_n236_), .B1(KEYINPUT9), .B2(new_n237_), .C1(G106gat), .C2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n235_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n203_), .B1(new_n234_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n216_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n204_), .B(new_n215_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n226_), .A2(KEYINPUT66), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n240_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(KEYINPUT67), .A3(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G57gat), .B(G64gat), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n248_), .A2(KEYINPUT11), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(KEYINPUT11), .ZN(new_n250_));
  XOR2_X1   g049(.A(G71gat), .B(G78gat), .Z(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n250_), .A2(new_n251_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT12), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n241_), .A2(new_n247_), .A3(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n227_), .A2(new_n233_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n240_), .B1(new_n260_), .B2(new_n242_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n261_), .B2(new_n254_), .ZN(new_n262_));
  AND2_X1   g061(.A1(G230gat), .A2(G233gat), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n261_), .B2(new_n254_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n261_), .A2(new_n254_), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n234_), .A2(new_n255_), .A3(new_n240_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n263_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G120gat), .B(G148gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT5), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G176gat), .B(G204gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n271_), .B(new_n272_), .Z(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT69), .B1(new_n269_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275_));
  INV_X1    g074(.A(new_n273_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n265_), .A2(new_n268_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n269_), .A2(new_n273_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(KEYINPUT70), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT70), .B1(new_n278_), .B2(new_n279_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n202_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n282_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(KEYINPUT13), .A3(new_n280_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT71), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(KEYINPUT72), .A3(new_n290_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G43gat), .B(G50gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT15), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n241_), .A2(new_n247_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT35), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G232gat), .A2(G233gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n261_), .A2(new_n299_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n305_), .A2(new_n302_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n301_), .A2(new_n306_), .A3(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G190gat), .B(G218gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT74), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G134gat), .B(G162gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT36), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT75), .Z(new_n318_));
  NAND3_X1  g117(.A1(new_n309_), .A2(new_n311_), .A3(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n319_), .A2(KEYINPUT76), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n315_), .B(new_n316_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT77), .ZN(new_n322_));
  INV_X1    g121(.A(new_n311_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n310_), .B1(new_n301_), .B2(new_n306_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT78), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(KEYINPUT76), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT78), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n328_), .B(new_n322_), .C1(new_n323_), .C2(new_n324_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n320_), .A2(new_n326_), .A3(new_n327_), .A4(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT37), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n319_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n332_), .A2(KEYINPUT37), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G15gat), .B(G22gat), .ZN(new_n335_));
  INV_X1    g134(.A(G1gat), .ZN(new_n336_));
  INV_X1    g135(.A(G8gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT14), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G1gat), .B(G8gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(new_n254_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G231gat), .A2(G233gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G127gat), .B(G155gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G183gat), .B(G211gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT17), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n349_), .B(KEYINPUT17), .Z(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n344_), .B2(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n353_), .B(KEYINPUT80), .Z(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n334_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n341_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n300_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT82), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G229gat), .A2(G233gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n341_), .A2(new_n299_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(KEYINPUT81), .B1(new_n341_), .B2(new_n299_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n341_), .A2(new_n299_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n360_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G113gat), .B(G141gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G169gat), .B(G197gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OR3_X1    g170(.A1(new_n362_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n362_), .B2(new_n367_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G127gat), .B(G134gat), .Z(new_n376_));
  XOR2_X1   g175(.A(G113gat), .B(G120gat), .Z(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT31), .Z(new_n379_));
  NAND2_X1  g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT23), .ZN(new_n381_));
  OR2_X1    g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT84), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n385_), .A3(new_n382_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT83), .B(G169gat), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n388_));
  OR3_X1    g187(.A1(new_n387_), .A2(KEYINPUT22), .A3(G176gat), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n384_), .A2(new_n386_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT25), .B(G183gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT26), .B(G190gat), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G169gat), .ZN(new_n395_));
  INV_X1    g194(.A(G176gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n394_), .B(new_n381_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n390_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G43gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n400_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(G15gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT30), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n403_), .B(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n379_), .B1(new_n408_), .B2(KEYINPUT85), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(KEYINPUT85), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G8gat), .B(G36gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT18), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G64gat), .B(G92gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n413_), .B(new_n414_), .Z(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G226gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT19), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT20), .ZN(new_n420_));
  XOR2_X1   g219(.A(G197gat), .B(G204gat), .Z(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT93), .ZN(new_n422_));
  XOR2_X1   g221(.A(G211gat), .B(G218gat), .Z(new_n423_));
  XNOR2_X1  g222(.A(G197gat), .B(G204gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT93), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n422_), .A2(KEYINPUT21), .A3(new_n423_), .A4(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n421_), .A2(KEYINPUT21), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT92), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n421_), .A2(KEYINPUT21), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n431_), .A2(new_n423_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n428_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT22), .B(G169gat), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n397_), .B1(new_n435_), .B2(new_n396_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT96), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n437_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n383_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n399_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n420_), .B1(new_n434_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n433_), .A2(new_n399_), .A3(new_n390_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n419_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n433_), .A2(new_n399_), .A3(new_n440_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n431_), .A2(new_n423_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n429_), .A2(KEYINPUT92), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n429_), .A2(KEYINPUT92), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n400_), .B1(new_n449_), .B2(new_n428_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n445_), .A2(new_n450_), .A3(KEYINPUT20), .A4(new_n419_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n416_), .B1(new_n444_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n441_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n443_), .B(KEYINPUT20), .C1(new_n433_), .C2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n418_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(new_n415_), .A3(new_n451_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G29gat), .ZN(new_n459_));
  INV_X1    g258(.A(G85gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT0), .B(G57gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G141gat), .A2(G148gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT3), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G141gat), .A2(G148gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT2), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n465_), .A2(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n470_), .A2(new_n471_), .ZN(new_n473_));
  OAI221_X1 g272(.A(new_n469_), .B1(new_n466_), .B2(new_n465_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n475_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G155gat), .B(G162gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(new_n477_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n467_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(new_n465_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n483_), .B(new_n484_), .C1(new_n478_), .C2(KEYINPUT1), .ZN(new_n485_));
  INV_X1    g284(.A(new_n378_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n481_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n477_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n480_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n485_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n378_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G225gat), .A2(G233gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n464_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT98), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(KEYINPUT98), .B(new_n464_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n493_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT97), .B1(new_n491_), .B2(KEYINPUT4), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n487_), .A2(new_n491_), .A3(KEYINPUT4), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT97), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT4), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n490_), .A2(new_n501_), .A3(new_n502_), .A4(new_n378_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n496_), .B(new_n497_), .C1(new_n498_), .C2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n498_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n492_), .A2(new_n493_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n464_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n458_), .B(new_n505_), .C1(KEYINPUT33), .C2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n508_), .A2(KEYINPUT33), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n506_), .A2(new_n464_), .A3(new_n507_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n511_), .A2(new_n508_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n445_), .A2(new_n450_), .A3(KEYINPUT20), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n418_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n442_), .A2(new_n419_), .A3(new_n443_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n444_), .A2(new_n452_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n415_), .A2(KEYINPUT32), .ZN(new_n518_));
  MUX2_X1   g317(.A(new_n516_), .B(new_n517_), .S(new_n518_), .Z(new_n519_));
  OAI22_X1  g318(.A1(new_n509_), .A2(new_n510_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G22gat), .B(G50gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT89), .B1(new_n490_), .B2(KEYINPUT29), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT29), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n481_), .A2(new_n524_), .A3(new_n525_), .A4(new_n485_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT91), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n523_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n522_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n532_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(new_n521_), .A3(new_n530_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G78gat), .B(G106gat), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n490_), .A2(KEYINPUT29), .ZN(new_n538_));
  INV_X1    g337(.A(G228gat), .ZN(new_n539_));
  INV_X1    g338(.A(G233gat), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n434_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n538_), .B2(new_n434_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n537_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n545_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(new_n543_), .A3(new_n536_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n533_), .A2(new_n535_), .A3(new_n546_), .A4(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n533_), .A2(new_n535_), .ZN(new_n551_));
  OAI22_X1  g350(.A1(new_n544_), .A2(new_n545_), .B1(KEYINPUT94), .B2(new_n537_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n537_), .A2(KEYINPUT94), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(new_n543_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT95), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n551_), .A2(new_n558_), .A3(new_n555_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n550_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n520_), .A2(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n551_), .A2(new_n558_), .A3(new_n555_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n558_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n549_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT27), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n517_), .B2(new_n415_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n516_), .A2(new_n416_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n453_), .A2(new_n457_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n566_), .A2(new_n567_), .B1(new_n568_), .B2(new_n565_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(new_n512_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n411_), .B1(new_n561_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n411_), .A2(new_n512_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n569_), .B(new_n549_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT99), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n557_), .A2(new_n559_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(KEYINPUT99), .A3(new_n549_), .A4(new_n569_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n572_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  NOR4_X1   g378(.A1(new_n296_), .A2(new_n356_), .A3(new_n375_), .A4(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n512_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n336_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT38), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n288_), .A2(new_n290_), .A3(new_n374_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n355_), .B(new_n332_), .C1(new_n571_), .C2(new_n578_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n336_), .B1(new_n588_), .B2(new_n581_), .ZN(new_n589_));
  OR3_X1    g388(.A1(new_n584_), .A2(new_n585_), .A3(new_n589_), .ZN(G1324gat));
  INV_X1    g389(.A(new_n569_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n337_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT39), .Z(new_n593_));
  NAND3_X1  g392(.A1(new_n580_), .A2(new_n337_), .A3(new_n591_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(G1325gat));
  NAND3_X1  g396(.A1(new_n580_), .A2(new_n405_), .A3(new_n411_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n405_), .B1(new_n588_), .B2(new_n411_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT41), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(G1326gat));
  INV_X1    g400(.A(G22gat), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n588_), .B2(new_n564_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT42), .Z(new_n604_));
  NAND3_X1  g403(.A1(new_n580_), .A2(new_n602_), .A3(new_n564_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(G1327gat));
  INV_X1    g405(.A(new_n586_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n579_), .A2(new_n355_), .A3(new_n332_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(G29gat), .B1(new_n610_), .B2(new_n581_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT43), .B1(new_n579_), .B2(new_n334_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n334_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n613_), .B(new_n614_), .C1(new_n571_), .C2(new_n578_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n616_), .A2(new_n586_), .A3(new_n355_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(KEYINPUT44), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(KEYINPUT44), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n581_), .A2(G29gat), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n611_), .B1(new_n620_), .B2(new_n621_), .ZN(G1328gat));
  OR2_X1    g421(.A1(new_n569_), .A2(G36gat), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n609_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT45), .Z(new_n625_));
  NAND3_X1  g424(.A1(new_n618_), .A2(new_n591_), .A3(new_n619_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(G36gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT101), .B(KEYINPUT46), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n628_), .B(new_n630_), .ZN(G1329gat));
  NAND3_X1  g430(.A1(new_n620_), .A2(G43gat), .A3(new_n411_), .ZN(new_n632_));
  AOI21_X1  g431(.A(G43gat), .B1(new_n610_), .B2(new_n411_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT102), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n632_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1330gat));
  NAND2_X1  g437(.A1(new_n620_), .A2(new_n564_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G50gat), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n560_), .A2(G50gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT104), .Z(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n609_), .B2(new_n642_), .ZN(G1331gat));
  NOR3_X1   g442(.A1(new_n295_), .A2(new_n374_), .A3(new_n587_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G57gat), .B1(new_n645_), .B2(new_n512_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n334_), .A2(new_n355_), .A3(new_n375_), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n579_), .B(new_n647_), .C1(new_n288_), .C2(new_n290_), .ZN(new_n648_));
  INV_X1    g447(.A(G57gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n581_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(new_n650_), .ZN(G1332gat));
  INV_X1    g450(.A(G64gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n644_), .B2(new_n591_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT48), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n648_), .A2(new_n652_), .A3(new_n591_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1333gat));
  INV_X1    g455(.A(G71gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n648_), .A2(new_n657_), .A3(new_n411_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n644_), .A2(new_n411_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT49), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n660_), .A3(G71gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n659_), .B2(G71gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT105), .B(new_n658_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1334gat));
  INV_X1    g467(.A(G78gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n644_), .B2(new_n564_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT50), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n648_), .A2(new_n669_), .A3(new_n564_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1335gat));
  NAND4_X1  g472(.A1(new_n293_), .A2(new_n294_), .A3(new_n375_), .A4(new_n608_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n675_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G85gat), .B1(new_n678_), .B2(new_n581_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n354_), .A2(new_n375_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n612_), .A2(new_n682_), .A3(new_n615_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT108), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n687_), .B(new_n681_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n686_), .A2(KEYINPUT109), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT109), .B1(new_n686_), .B2(new_n688_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n512_), .A2(new_n460_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n679_), .B1(new_n691_), .B2(new_n692_), .ZN(G1336gat));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n591_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G92gat), .ZN(new_n696_));
  INV_X1    g495(.A(G92gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n591_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n694_), .B1(new_n696_), .B2(new_n700_), .ZN(new_n701_));
  AOI211_X1 g500(.A(KEYINPUT110), .B(new_n699_), .C1(new_n695_), .C2(G92gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1337gat));
  INV_X1    g502(.A(new_n238_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n678_), .A2(new_n704_), .A3(new_n411_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n686_), .A2(new_n411_), .A3(new_n688_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G99gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g508(.A(G106gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n678_), .A2(new_n710_), .A3(new_n564_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n616_), .A2(new_n560_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n681_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G106gat), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT52), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT111), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n714_), .B(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(KEYINPUT111), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n711_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT53), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT53), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n711_), .B(new_n721_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1339gat));
  INV_X1    g522(.A(KEYINPUT117), .ZN(new_n724_));
  XOR2_X1   g523(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT113), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n647_), .A2(new_n286_), .A3(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n726_), .A2(KEYINPUT113), .ZN(new_n730_));
  OAI22_X1  g529(.A1(new_n647_), .A2(new_n286_), .B1(new_n730_), .B2(new_n728_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n278_), .A2(new_n374_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735_));
  INV_X1    g534(.A(new_n267_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n258_), .A2(new_n736_), .A3(new_n262_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n265_), .A2(KEYINPUT55), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n258_), .A2(new_n262_), .A3(new_n264_), .A4(new_n739_), .ZN(new_n740_));
  AOI221_X4 g539(.A(new_n735_), .B1(new_n737_), .B2(new_n263_), .C1(new_n738_), .C2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n740_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n737_), .A2(new_n263_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT114), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n273_), .B1(new_n741_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT56), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(KEYINPUT56), .B(new_n273_), .C1(new_n741_), .C2(new_n744_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n734_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n359_), .A2(new_n366_), .A3(new_n361_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n370_), .B1(new_n365_), .B2(new_n360_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n372_), .A2(KEYINPUT115), .A3(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT115), .B1(new_n372_), .B2(new_n752_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n284_), .B2(new_n280_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n332_), .B1(new_n749_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT57), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n759_), .B(new_n332_), .C1(new_n749_), .C2(new_n756_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n755_), .B1(new_n274_), .B2(new_n277_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n742_), .A2(new_n743_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n735_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n742_), .A2(KEYINPUT114), .A3(new_n743_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n273_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n748_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n761_), .B(KEYINPUT58), .C1(new_n766_), .C2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n761_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n334_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n758_), .A2(new_n760_), .B1(new_n768_), .B2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n355_), .B1(new_n772_), .B2(KEYINPUT116), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n768_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n734_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n776_));
  OAI22_X1  g575(.A1(new_n281_), .A2(new_n282_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n759_), .B1(new_n778_), .B2(new_n332_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n760_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n774_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n733_), .B1(new_n773_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n575_), .A2(new_n577_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n581_), .A3(new_n411_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n724_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT116), .B(new_n774_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n354_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n772_), .A2(KEYINPUT116), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n732_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n786_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(KEYINPUT117), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n374_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(G113gat), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT118), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n794_), .A2(new_n798_), .A3(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n781_), .A2(new_n354_), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT59), .B(new_n786_), .C1(new_n800_), .C2(new_n732_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n791_), .A2(new_n792_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(KEYINPUT59), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n375_), .A2(new_n795_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n797_), .A2(new_n799_), .B1(new_n803_), .B2(new_n804_), .ZN(G1340gat));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806_));
  INV_X1    g605(.A(G120gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n803_), .B2(new_n296_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT60), .ZN(new_n809_));
  AOI21_X1  g608(.A(G120gat), .B1(new_n291_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n809_), .B2(G120gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n787_), .A2(new_n793_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n806_), .B1(new_n808_), .B2(new_n813_), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n295_), .B(new_n801_), .C1(new_n802_), .C2(KEYINPUT59), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT119), .B(new_n812_), .C1(new_n815_), .C2(new_n807_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1341gat));
  AND2_X1   g616(.A1(new_n787_), .A2(new_n793_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G127gat), .B1(new_n818_), .B2(new_n355_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n355_), .A2(G127gat), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT120), .Z(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n803_), .B2(new_n821_), .ZN(G1342gat));
  INV_X1    g621(.A(G134gat), .ZN(new_n823_));
  INV_X1    g622(.A(new_n332_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n818_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n803_), .A2(new_n613_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n823_), .ZN(G1343gat));
  NOR2_X1   g626(.A1(new_n784_), .A2(new_n411_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n560_), .A2(new_n512_), .A3(new_n591_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n374_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n296_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g633(.A1(new_n828_), .A2(new_n829_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n354_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT61), .B(G155gat), .Z(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1346gat));
  OAI21_X1  g637(.A(G162gat), .B1(new_n835_), .B2(new_n334_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n332_), .A2(G162gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n835_), .B2(new_n840_), .ZN(G1347gat));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n800_), .A2(new_n732_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n411_), .A2(new_n512_), .A3(new_n591_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT121), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n564_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n374_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n374_), .A3(new_n435_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT62), .B1(new_n848_), .B2(G169gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n842_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n848_), .A2(G169gat), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n856_), .A2(KEYINPUT122), .A3(new_n850_), .A4(new_n849_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(G1348gat));
  AOI21_X1  g657(.A(G176gat), .B1(new_n847_), .B2(new_n291_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT123), .B1(new_n784_), .B2(new_n564_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n791_), .A2(new_n861_), .A3(new_n560_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n295_), .A2(new_n396_), .A3(new_n845_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT124), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n863_), .A2(new_n867_), .A3(new_n864_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n859_), .B1(new_n866_), .B2(new_n868_), .ZN(G1349gat));
  NAND2_X1  g668(.A1(new_n843_), .A2(new_n846_), .ZN(new_n870_));
  OR3_X1    g669(.A1(new_n870_), .A2(new_n354_), .A3(new_n392_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n845_), .A2(new_n354_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n871_), .B1(new_n874_), .B2(G183gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT125), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n871_), .B(new_n877_), .C1(new_n874_), .C2(G183gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n870_), .B2(new_n334_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n824_), .A2(new_n393_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT126), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n870_), .B2(new_n882_), .ZN(G1351gat));
  NOR3_X1   g682(.A1(new_n560_), .A2(new_n581_), .A3(new_n569_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n828_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n374_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n296_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g688(.A(new_n354_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n885_), .A2(new_n890_), .ZN(new_n891_));
  OR2_X1    g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1354gat));
  INV_X1    g692(.A(new_n885_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G218gat), .B1(new_n894_), .B2(new_n334_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n332_), .A2(G218gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n894_), .B2(new_n896_), .ZN(G1355gat));
endmodule


