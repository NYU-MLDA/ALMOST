//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G231gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT79), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n208_), .B(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G71gat), .B(G78gat), .Z(new_n212_));
  INV_X1    g011(.A(G57gat), .ZN(new_n213_));
  INV_X1    g012(.A(G64gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G57gat), .A2(G64gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n216_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT70), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT69), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT69), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT70), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(G57gat), .A2(G64gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G57gat), .A2(G64gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT11), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n219_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n220_), .A2(new_n225_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(new_n230_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n218_), .A4(new_n212_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n211_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT16), .B(G183gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G211gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(G127gat), .B(G155gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT17), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n241_), .A2(new_n242_), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n237_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n237_), .A2(new_n243_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n246_), .A2(KEYINPUT80), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(KEYINPUT80), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n245_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G43gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G169gat), .ZN(new_n255_));
  INV_X1    g054(.A(G176gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(KEYINPUT24), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n257_), .A2(KEYINPUT24), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G190gat), .ZN(new_n262_));
  OR3_X1    g061(.A1(new_n262_), .A2(KEYINPUT82), .A3(KEYINPUT26), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT25), .B(G183gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT26), .B1(new_n262_), .B2(KEYINPUT82), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n259_), .A2(new_n261_), .A3(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT22), .B(G169gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n256_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n269_), .B(new_n260_), .C1(new_n254_), .C2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT83), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n273_), .A2(new_n274_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278_));
  INV_X1    g077(.A(G15gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n276_), .A2(new_n277_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n272_), .B(KEYINPUT83), .Z(new_n283_));
  INV_X1    g082(.A(new_n274_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n282_), .B1(new_n285_), .B2(new_n275_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n251_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n280_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n251_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n285_), .A2(new_n275_), .A3(new_n282_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G127gat), .B(G134gat), .Z(new_n293_));
  XOR2_X1   g092(.A(G113gat), .B(G120gat), .Z(new_n294_));
  OR2_X1    g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n294_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT85), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT31), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT86), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n292_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT86), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n287_), .A2(new_n304_), .A3(new_n301_), .A4(new_n291_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G78gat), .B(G106gat), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT3), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT2), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(KEYINPUT1), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n311_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT89), .B1(new_n323_), .B2(KEYINPUT29), .ZN(new_n324_));
  XOR2_X1   g123(.A(G197gat), .B(G204gat), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT21), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n325_), .A2(KEYINPUT21), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n324_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n335_), .B(KEYINPUT88), .Z(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n324_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n308_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT91), .Z(new_n341_));
  OR2_X1    g140(.A1(new_n323_), .A2(KEYINPUT29), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G22gat), .B(G50gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT28), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n342_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n338_), .A2(new_n308_), .A3(new_n339_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT92), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n341_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT93), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n347_), .B1(new_n340_), .B2(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n338_), .A2(KEYINPUT93), .A3(new_n308_), .A4(new_n339_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n345_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n349_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n306_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n303_), .A2(new_n305_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(new_n354_), .A3(new_n349_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n317_), .A2(new_n322_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n295_), .A2(new_n297_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n323_), .A2(new_n300_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT4), .ZN(new_n365_));
  INV_X1    g164(.A(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n365_), .B1(KEYINPUT4), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(G225gat), .A3(G233gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n362_), .A2(new_n369_), .A3(new_n363_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT0), .B(G57gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G85gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(G1gat), .B(G29gat), .Z(new_n374_));
  XOR2_X1   g173(.A(new_n373_), .B(new_n374_), .Z(new_n375_));
  NAND2_X1  g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n368_), .A2(new_n370_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT26), .B(G190gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n264_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n261_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT94), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n259_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n271_), .B(KEYINPUT95), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n333_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n388_), .B(KEYINPUT20), .C1(new_n283_), .C2(new_n333_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G8gat), .B(G36gat), .Z(new_n393_));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n395_), .B(new_n396_), .Z(new_n397_));
  NAND2_X1  g196(.A1(new_n283_), .A2(new_n333_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n333_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n391_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n398_), .A2(new_n400_), .A3(KEYINPUT20), .A4(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n392_), .A2(new_n397_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT27), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n389_), .A2(new_n391_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(new_n271_), .A3(new_n385_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n398_), .A2(KEYINPUT20), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n391_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n397_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n404_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT98), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT27), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n392_), .A2(new_n402_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n414_), .A2(new_n397_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n403_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n413_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT98), .B1(new_n404_), .B2(new_n409_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n412_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n359_), .A2(new_n380_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n367_), .A2(new_n369_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n364_), .B(KEYINPUT97), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n422_), .B(new_n375_), .C1(new_n369_), .C2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n378_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT33), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n415_), .A2(new_n416_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n378_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n426_), .B(new_n427_), .C1(KEYINPUT33), .C2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n397_), .A2(KEYINPUT32), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n414_), .A2(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n405_), .A2(new_n408_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n379_), .B(new_n431_), .C1(new_n432_), .C2(new_n430_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n306_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n355_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n421_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT76), .B(G43gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G50gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(G29gat), .B(G36gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT15), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(KEYINPUT66), .B(G106gat), .Z(new_n443_));
  INV_X1    g242(.A(G99gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT10), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT10), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(G99gat), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n445_), .A2(new_n447_), .A3(KEYINPUT65), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT65), .B1(new_n445_), .B2(new_n447_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n443_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(G85gat), .ZN(new_n451_));
  INV_X1    g250(.A(G92gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT67), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT9), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT9), .ZN(new_n455_));
  OAI211_X1 g254(.A(KEYINPUT67), .B(new_n455_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n454_), .B(new_n456_), .C1(G85gat), .C2(G92gat), .ZN(new_n457_));
  AND3_X1   g256(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n450_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT8), .ZN(new_n462_));
  XOR2_X1   g261(.A(G85gat), .B(G92gat), .Z(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  INV_X1    g263(.A(G106gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n444_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT68), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n467_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n444_), .B(new_n465_), .C1(new_n471_), .C2(KEYINPUT68), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(KEYINPUT68), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n462_), .B(new_n463_), .C1(new_n470_), .C2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n460_), .A2(new_n468_), .A3(new_n473_), .A4(new_n472_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n462_), .B1(new_n477_), .B2(new_n463_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n461_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT77), .B1(new_n442_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G232gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT34), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(KEYINPUT35), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n440_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(new_n442_), .B2(new_n480_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(KEYINPUT35), .A3(new_n483_), .A4(new_n481_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G190gat), .B(G218gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G134gat), .ZN(new_n492_));
  INV_X1    g291(.A(G162gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(KEYINPUT36), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n483_), .A2(KEYINPUT35), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(KEYINPUT36), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n490_), .A2(new_n497_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n487_), .A2(new_n489_), .A3(new_n498_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n501_), .A2(KEYINPUT78), .A3(new_n496_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT78), .B1(new_n501_), .B2(new_n496_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n500_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT100), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT72), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n463_), .B1(new_n470_), .B2(new_n474_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT8), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n475_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n236_), .B1(new_n510_), .B2(new_n461_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n507_), .B1(new_n511_), .B2(KEYINPUT12), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n232_), .A2(new_n235_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n479_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT12), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(KEYINPUT72), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n479_), .A2(KEYINPUT12), .A3(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT71), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT71), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n479_), .A2(new_n513_), .A3(new_n519_), .A4(KEYINPUT12), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n512_), .A2(new_n516_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G230gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT64), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(new_n479_), .B2(new_n513_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT73), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n527_), .B(new_n524_), .C1(new_n479_), .C2(new_n513_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n521_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n480_), .A2(new_n236_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n514_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n523_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT74), .B(G204gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G120gat), .B(G148gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT5), .B(G176gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n530_), .A2(new_n533_), .A3(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(KEYINPUT75), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT75), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n534_), .A2(new_n544_), .A3(new_n539_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(KEYINPUT13), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT13), .B1(new_n543_), .B2(new_n545_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n208_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n440_), .B(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n440_), .A2(new_n550_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n442_), .B2(new_n550_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n554_), .B1(new_n556_), .B2(new_n553_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G169gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(G197gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n557_), .B(new_n560_), .Z(new_n561_));
  NOR2_X1   g360(.A1(new_n549_), .A2(new_n561_), .ZN(new_n562_));
  AND4_X1   g361(.A1(new_n249_), .A2(new_n436_), .A3(new_n506_), .A4(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT101), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n202_), .B1(new_n564_), .B2(new_n379_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT102), .Z(new_n566_));
  AOI21_X1  g365(.A(new_n419_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n567_), .A2(new_n380_), .B1(new_n434_), .B2(new_n355_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n561_), .B(KEYINPUT81), .Z(new_n569_));
  NOR3_X1   g368(.A1(new_n568_), .A2(new_n549_), .A3(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n504_), .B(KEYINPUT37), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n249_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(new_n202_), .A3(new_n379_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT38), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT103), .Z(new_n578_));
  NOR2_X1   g377(.A1(new_n575_), .A2(new_n576_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT99), .Z(new_n580_));
  NAND3_X1  g379(.A1(new_n566_), .A2(new_n578_), .A3(new_n580_), .ZN(G1324gat));
  AOI21_X1  g380(.A(new_n204_), .B1(new_n563_), .B2(new_n419_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT39), .Z(new_n583_));
  NAND3_X1  g382(.A1(new_n574_), .A2(new_n204_), .A3(new_n419_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g385(.A1(new_n574_), .A2(new_n279_), .A3(new_n306_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n564_), .A2(new_n306_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n588_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT41), .B1(new_n588_), .B2(G15gat), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n587_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT104), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(KEYINPUT104), .B(new_n587_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(G1326gat));
  INV_X1    g394(.A(G22gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n355_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n564_), .B2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT42), .Z(new_n599_));
  NAND3_X1  g398(.A1(new_n574_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(G1327gat));
  INV_X1    g400(.A(new_n249_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n568_), .A2(KEYINPUT43), .A3(new_n571_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT43), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n504_), .B(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n604_), .B1(new_n436_), .B2(new_n606_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n602_), .B(new_n562_), .C1(new_n603_), .C2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT44), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT43), .B1(new_n568_), .B2(new_n571_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n436_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n613_), .A2(KEYINPUT44), .A3(new_n602_), .A4(new_n562_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G29gat), .B1(new_n615_), .B2(new_n380_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n506_), .A2(new_n249_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n570_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n619_), .A2(G29gat), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n616_), .B1(new_n380_), .B2(new_n620_), .ZN(G1328gat));
  INV_X1    g420(.A(KEYINPUT107), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT46), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n610_), .A2(new_n419_), .A3(new_n614_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT105), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n610_), .A2(new_n628_), .A3(new_n419_), .A4(new_n614_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(G36gat), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT106), .ZN(new_n631_));
  INV_X1    g430(.A(G36gat), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n618_), .A2(new_n631_), .A3(new_n632_), .A4(new_n419_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n570_), .A2(new_n632_), .A3(new_n617_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT106), .B1(new_n634_), .B2(new_n420_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n633_), .A2(KEYINPUT45), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT45), .B1(new_n633_), .B2(new_n635_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AOI211_X1 g437(.A(new_n624_), .B(new_n625_), .C1(new_n630_), .C2(new_n638_), .ZN(new_n639_));
  AND4_X1   g438(.A1(new_n622_), .A2(new_n630_), .A3(new_n623_), .A4(new_n638_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1329gat));
  OAI21_X1  g440(.A(G43gat), .B1(new_n615_), .B2(new_n357_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n357_), .A2(G43gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n642_), .B1(new_n619_), .B2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g444(.A(G50gat), .B1(new_n615_), .B2(new_n355_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n355_), .A2(G50gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n619_), .B2(new_n647_), .ZN(G1331gat));
  INV_X1    g447(.A(new_n549_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n602_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n436_), .A2(new_n506_), .A3(new_n569_), .A4(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT109), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(G57gat), .A3(new_n379_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(KEYINPUT110), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n573_), .A2(new_n549_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT108), .ZN(new_n656_));
  INV_X1    g455(.A(new_n561_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n568_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n213_), .B1(new_n659_), .B2(new_n380_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n653_), .A2(KEYINPUT110), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n654_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT111), .ZN(G1332gat));
  INV_X1    g462(.A(new_n659_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n214_), .A3(new_n419_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n652_), .A2(new_n419_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G64gat), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT112), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(KEYINPUT112), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(KEYINPUT48), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT48), .B1(new_n668_), .B2(new_n669_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n665_), .B1(new_n670_), .B2(new_n671_), .ZN(G1333gat));
  INV_X1    g471(.A(G71gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n652_), .B2(new_n306_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT49), .Z(new_n675_));
  NAND3_X1  g474(.A1(new_n664_), .A2(new_n673_), .A3(new_n306_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1334gat));
  INV_X1    g476(.A(G78gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n652_), .B2(new_n597_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT50), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n664_), .A2(new_n678_), .A3(new_n597_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1335gat));
  AND3_X1   g481(.A1(new_n658_), .A2(new_n549_), .A3(new_n617_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n451_), .A3(new_n379_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n649_), .A2(new_n249_), .A3(new_n657_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n613_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT113), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT114), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(KEYINPUT114), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(new_n379_), .A3(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n684_), .B1(new_n690_), .B2(new_n451_), .ZN(G1336gat));
  NAND3_X1  g490(.A1(new_n683_), .A2(new_n452_), .A3(new_n419_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n688_), .A2(new_n419_), .A3(new_n689_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n452_), .ZN(G1337gat));
  OAI211_X1 g493(.A(new_n683_), .B(new_n306_), .C1(new_n449_), .C2(new_n448_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n687_), .A2(new_n306_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(G99gat), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g498(.A(KEYINPUT53), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n683_), .A2(new_n443_), .A3(new_n597_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n613_), .A2(new_n597_), .A3(new_n685_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT52), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(G106gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n702_), .B2(G106gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT115), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n706_), .A2(KEYINPUT115), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n700_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n709_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(KEYINPUT53), .A3(new_n707_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1339gat));
  NAND3_X1  g512(.A1(new_n573_), .A2(new_n649_), .A3(new_n569_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT54), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT54), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n573_), .A2(new_n716_), .A3(new_n649_), .A4(new_n569_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT57), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n551_), .A2(new_n552_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n556_), .B2(new_n552_), .ZN(new_n720_));
  MUX2_X1   g519(.A(new_n557_), .B(new_n720_), .S(new_n560_), .Z(new_n721_));
  NAND3_X1  g520(.A1(new_n543_), .A2(new_n545_), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT55), .B1(new_n521_), .B2(new_n529_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n512_), .A2(new_n516_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n518_), .A2(new_n520_), .ZN(new_n726_));
  AND4_X1   g525(.A1(KEYINPUT55), .A2(new_n529_), .A3(new_n725_), .A4(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n726_), .A3(new_n531_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT116), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT116), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n725_), .A2(new_n726_), .A3(new_n731_), .A4(new_n531_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n730_), .A2(new_n523_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n728_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT56), .B1(new_n734_), .B2(new_n539_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT56), .ZN(new_n736_));
  AOI211_X1 g535(.A(new_n736_), .B(new_n541_), .C1(new_n728_), .C2(new_n733_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT117), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n561_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n542_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n735_), .B2(KEYINPUT117), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n723_), .B1(new_n740_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n504_), .B(KEYINPUT100), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n718_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n735_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n737_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n739_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(new_n657_), .A3(new_n742_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n722_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n506_), .A3(KEYINPUT57), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n746_), .A2(new_n747_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(new_n542_), .A3(new_n721_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT58), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n752_), .A2(KEYINPUT58), .A3(new_n542_), .A4(new_n721_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n606_), .A3(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n745_), .A2(new_n751_), .A3(new_n757_), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n715_), .A2(new_n717_), .B1(new_n758_), .B2(new_n602_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n356_), .A2(new_n419_), .A3(new_n380_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G113gat), .B1(new_n762_), .B2(new_n657_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n715_), .A2(new_n717_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n758_), .A2(KEYINPUT118), .A3(new_n602_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT118), .B1(new_n758_), .B2(new_n602_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT59), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n760_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT59), .B1(new_n759_), .B2(new_n761_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n569_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n763_), .B1(new_n772_), .B2(G113gat), .ZN(G1340gat));
  XOR2_X1   g572(.A(KEYINPUT119), .B(G120gat), .Z(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n771_), .B2(new_n649_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n774_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n649_), .B2(KEYINPUT60), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n762_), .B(new_n777_), .C1(KEYINPUT60), .C2(new_n776_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n775_), .A2(new_n778_), .ZN(G1341gat));
  AOI21_X1  g578(.A(G127gat), .B1(new_n762_), .B2(new_n249_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n769_), .A2(G127gat), .A3(new_n770_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n249_), .ZN(G1342gat));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n769_), .A2(new_n606_), .A3(new_n770_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(G134gat), .ZN(new_n785_));
  NOR4_X1   g584(.A1(new_n759_), .A2(G134gat), .A3(new_n506_), .A4(new_n761_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n783_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT120), .B(new_n786_), .C1(new_n784_), .C2(G134gat), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1343gat));
  NOR2_X1   g589(.A1(new_n759_), .A2(new_n358_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n419_), .A2(new_n380_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(new_n561_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g594(.A1(new_n793_), .A2(new_n649_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g596(.A1(new_n793_), .A2(new_n602_), .ZN(new_n798_));
  XOR2_X1   g597(.A(KEYINPUT61), .B(G155gat), .Z(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(G1346gat));
  NOR3_X1   g599(.A1(new_n793_), .A2(new_n493_), .A3(new_n571_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n791_), .A2(new_n744_), .A3(new_n792_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n493_), .B2(new_n802_), .ZN(G1347gat));
  XNOR2_X1  g602(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(KEYINPUT122), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(KEYINPUT122), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n420_), .A2(new_n379_), .A3(new_n356_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n767_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n561_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n807_), .B(new_n808_), .C1(new_n811_), .C2(new_n255_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n268_), .ZN(new_n813_));
  OAI211_X1 g612(.A(G169gat), .B(new_n806_), .C1(new_n810_), .C2(new_n561_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(new_n813_), .A3(new_n814_), .ZN(G1348gat));
  INV_X1    g614(.A(new_n809_), .ZN(new_n816_));
  NOR4_X1   g615(.A1(new_n759_), .A2(new_n256_), .A3(new_n649_), .A4(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n256_), .B1(new_n810_), .B2(new_n649_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n819_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n817_), .B1(new_n820_), .B2(new_n821_), .ZN(G1349gat));
  NOR3_X1   g621(.A1(new_n759_), .A2(new_n602_), .A3(new_n816_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT125), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(G183gat), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n824_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n602_), .A2(new_n264_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n767_), .A2(KEYINPUT124), .A3(new_n809_), .A4(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT124), .ZN(new_n831_));
  INV_X1    g630(.A(new_n829_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n810_), .B2(new_n832_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n828_), .A2(new_n830_), .A3(new_n833_), .ZN(G1350gat));
  OAI21_X1  g633(.A(G190gat), .B1(new_n810_), .B2(new_n571_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n744_), .A2(new_n381_), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT126), .Z(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n810_), .B2(new_n837_), .ZN(G1351gat));
  NOR2_X1   g637(.A1(new_n420_), .A2(new_n379_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n791_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n561_), .ZN(new_n841_));
  XOR2_X1   g640(.A(new_n841_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n649_), .ZN(new_n843_));
  INV_X1    g642(.A(G204gat), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(KEYINPUT127), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n843_), .B(new_n845_), .Z(G1353gat));
  NOR2_X1   g645(.A1(new_n840_), .A2(new_n602_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n847_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT63), .B(G211gat), .Z(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n847_), .B2(new_n849_), .ZN(G1354gat));
  NOR2_X1   g649(.A1(new_n840_), .A2(new_n506_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(G218gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n840_), .A2(new_n571_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(G218gat), .B2(new_n853_), .ZN(G1355gat));
endmodule


