//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_;
  XNOR2_X1  g000(.A(KEYINPUT75), .B(G43gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT31), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT23), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT73), .B(KEYINPUT23), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(new_n205_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n208_), .B2(KEYINPUT74), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n209_), .B1(KEYINPUT74), .B2(new_n208_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OR3_X1    g012(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G169gat), .B(G176gat), .Z(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(KEYINPUT24), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n210_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n205_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT23), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(new_n207_), .B2(new_n219_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(G169gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT30), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G227gat), .A2(G233gat), .ZN(new_n228_));
  INV_X1    g027(.A(G15gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(G71gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G99gat), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234_));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT76), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n234_), .A2(new_n235_), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  NAND2_X1  g038(.A1(new_n227_), .A2(new_n232_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n233_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n239_), .B1(new_n233_), .B2(new_n240_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n204_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(new_n241_), .A3(new_n203_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT77), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(G155gat), .B2(G162gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G141gat), .A2(G148gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n255_), .A2(KEYINPUT2), .ZN(new_n256_));
  OR2_X1    g055(.A1(G141gat), .A2(G148gat), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT3), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(KEYINPUT3), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n258_), .B(new_n259_), .C1(new_n255_), .C2(KEYINPUT2), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n252_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT29), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT1), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n257_), .B(new_n253_), .C1(new_n251_), .C2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT28), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G22gat), .B(G50gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT79), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT79), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT80), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G197gat), .B(G204gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT21), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n279_), .B(new_n280_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT81), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G228gat), .A2(G233gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n261_), .A2(new_n265_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT29), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G78gat), .B(G106gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT82), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n290_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(G228gat), .A3(G233gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n295_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n293_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n275_), .A2(new_n276_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n296_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n292_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n291_), .B2(new_n295_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n301_), .A2(new_n273_), .A3(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n248_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G226gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT19), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n210_), .B1(G183gat), .B2(G190gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n310_), .A2(new_n224_), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT83), .B(KEYINPUT24), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n313_), .A2(G169gat), .A3(G176gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n216_), .ZN(new_n315_));
  AND4_X1   g114(.A1(new_n221_), .A2(new_n314_), .A3(new_n213_), .A4(new_n315_), .ZN(new_n316_));
  NOR4_X1   g115(.A1(new_n311_), .A2(new_n283_), .A3(new_n285_), .A4(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n317_), .A2(KEYINPUT85), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT20), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n287_), .B2(new_n226_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(new_n317_), .B2(KEYINPUT85), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n309_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n311_), .A2(new_n316_), .ZN(new_n323_));
  OR3_X1    g122(.A1(new_n323_), .A2(KEYINPUT84), .A3(new_n286_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n287_), .A2(new_n226_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(new_n319_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT84), .B1(new_n323_), .B2(new_n286_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n324_), .A2(new_n326_), .A3(new_n308_), .A4(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n322_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT18), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n333_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n322_), .A2(new_n335_), .A3(new_n328_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT86), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(G85gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT0), .B(G57gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n239_), .A2(new_n289_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n289_), .B1(new_n238_), .B2(new_n236_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT4), .ZN(new_n348_));
  XOR2_X1   g147(.A(KEYINPUT88), .B(KEYINPUT4), .Z(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT89), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n345_), .A2(KEYINPUT89), .A3(new_n349_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(KEYINPUT87), .A2(new_n348_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n348_), .A2(KEYINPUT87), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n344_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n344_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n347_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n343_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT33), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n354_), .A2(new_n355_), .A3(new_n344_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n343_), .B1(new_n347_), .B2(new_n357_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n359_), .A2(new_n360_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n334_), .A2(KEYINPUT86), .A3(new_n336_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n339_), .A2(new_n361_), .A3(new_n364_), .A4(new_n365_), .ZN(new_n366_));
  OR3_X1    g165(.A1(new_n356_), .A2(new_n343_), .A3(new_n358_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n359_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n324_), .A2(new_n326_), .A3(new_n309_), .A4(new_n327_), .ZN(new_n369_));
  AOI211_X1 g168(.A(new_n319_), .B(new_n317_), .C1(new_n226_), .C2(new_n287_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n309_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(KEYINPUT32), .A3(new_n333_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n333_), .A2(KEYINPUT32), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n329_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT90), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n329_), .A2(KEYINPUT90), .A3(new_n373_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n368_), .A2(new_n372_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n306_), .B1(new_n366_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n247_), .A2(new_n305_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n244_), .B(new_n246_), .C1(new_n300_), .C2(new_n304_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n368_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n329_), .B2(new_n333_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n371_), .A2(new_n335_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n337_), .A2(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n379_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G29gat), .B(G36gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G43gat), .B(G50gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT15), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G15gat), .B(G22gat), .ZN(new_n393_));
  INV_X1    g192(.A(G1gat), .ZN(new_n394_));
  INV_X1    g193(.A(G8gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT14), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G1gat), .B(G8gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n392_), .A2(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n389_), .B(new_n390_), .Z(new_n401_));
  OR2_X1    g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G229gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT72), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT70), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n402_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT71), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n399_), .A2(new_n401_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n407_), .B1(new_n412_), .B2(new_n404_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G113gat), .B(G141gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G169gat), .B(G197gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n414_), .B(new_n415_), .Z(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n407_), .B(new_n416_), .C1(new_n412_), .C2(new_n404_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n388_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT65), .B(KEYINPUT12), .ZN(new_n423_));
  INV_X1    g222(.A(G85gat), .ZN(new_n424_));
  INV_X1    g223(.A(G92gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT9), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G85gat), .A2(G92gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT64), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n426_), .B(new_n427_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n426_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n428_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G99gat), .A2(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT6), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(G99gat), .A3(G106gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n438_));
  INV_X1    g237(.A(G106gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n431_), .A2(new_n432_), .A3(new_n437_), .A4(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n426_), .A2(new_n428_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n434_), .A2(new_n436_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT7), .ZN(new_n447_));
  INV_X1    g246(.A(G99gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n439_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n445_), .B1(new_n446_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT8), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n437_), .A2(new_n450_), .A3(new_n449_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT8), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n445_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n443_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G57gat), .B(G64gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G71gat), .B(G78gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(KEYINPUT11), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  INV_X1    g260(.A(G64gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G57gat), .ZN(new_n463_));
  INV_X1    g262(.A(G57gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(G64gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n465_), .A3(KEYINPUT11), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n458_), .A2(KEYINPUT11), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n460_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n423_), .B1(new_n457_), .B2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n449_), .A2(new_n450_), .ZN(new_n471_));
  AOI211_X1 g270(.A(KEYINPUT8), .B(new_n444_), .C1(new_n471_), .C2(new_n437_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n455_), .B1(new_n454_), .B2(new_n445_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n442_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n469_), .ZN(new_n475_));
  OR2_X1    g274(.A1(KEYINPUT65), .A2(KEYINPUT12), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n442_), .B(new_n469_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G230gat), .A2(G233gat), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n478_), .A2(KEYINPUT66), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT66), .B1(new_n478_), .B2(new_n479_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n470_), .B(new_n477_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n479_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n457_), .A2(new_n469_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n478_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G120gat), .B(G148gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT5), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G176gat), .B(G204gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT67), .Z(new_n494_));
  OR2_X1    g293(.A1(new_n487_), .A2(new_n492_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT13), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n497_), .A2(KEYINPUT68), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(KEYINPUT68), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n496_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n496_), .A2(new_n499_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G232gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT34), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(KEYINPUT35), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n392_), .B2(new_n474_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n506_), .B1(new_n401_), .B2(new_n474_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(KEYINPUT35), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G190gat), .B(G218gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G134gat), .B(G162gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(KEYINPUT36), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n512_), .B(KEYINPUT36), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT37), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n399_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(new_n475_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G127gat), .B(G155gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT16), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G183gat), .B(G211gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n527_), .A2(KEYINPUT69), .ZN(new_n528_));
  OR3_X1    g327(.A1(new_n522_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n527_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n522_), .B(new_n530_), .C1(new_n526_), .C2(new_n528_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n518_), .A2(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n502_), .A2(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n422_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n368_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n535_), .A2(G1gat), .A3(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n388_), .A2(new_n517_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n500_), .A2(new_n501_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n421_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n502_), .A2(KEYINPUT92), .A3(new_n420_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n532_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n540_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(G1gat), .B1(new_n547_), .B2(new_n536_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n539_), .A2(new_n548_), .ZN(G1324gat));
  INV_X1    g348(.A(new_n386_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n395_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT93), .B1(new_n535_), .B2(new_n551_), .ZN(new_n552_));
  OR4_X1    g351(.A1(KEYINPUT93), .A2(new_n422_), .A3(new_n534_), .A4(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(G8gat), .B1(new_n547_), .B2(new_n386_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT39), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI211_X1 g356(.A(KEYINPUT39), .B(G8gat), .C1(new_n547_), .C2(new_n386_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT40), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(G1325gat));
  OAI21_X1  g360(.A(G15gat), .B1(new_n547_), .B2(new_n248_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT41), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n247_), .A2(new_n229_), .ZN(new_n566_));
  OAI22_X1  g365(.A1(new_n564_), .A2(new_n565_), .B1(new_n535_), .B2(new_n566_), .ZN(G1326gat));
  OAI21_X1  g366(.A(G22gat), .B1(new_n547_), .B2(new_n305_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n568_), .A2(KEYINPUT42), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(KEYINPUT42), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n305_), .A2(G22gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT94), .ZN(new_n572_));
  OAI22_X1  g371(.A1(new_n569_), .A2(new_n570_), .B1(new_n535_), .B2(new_n572_), .ZN(G1327gat));
  INV_X1    g372(.A(new_n517_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n545_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n502_), .A2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n421_), .B(new_n576_), .C1(new_n379_), .C2(new_n387_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(G29gat), .B1(new_n578_), .B2(new_n368_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n518_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n379_), .B2(new_n387_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT43), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT43), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n583_), .B(new_n580_), .C1(new_n379_), .C2(new_n387_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n543_), .A2(new_n544_), .A3(new_n532_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(KEYINPUT95), .A2(KEYINPUT44), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n585_), .A2(new_n588_), .A3(new_n586_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n368_), .A2(G29gat), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n579_), .B1(new_n592_), .B2(new_n593_), .ZN(G1328gat));
  INV_X1    g393(.A(KEYINPUT45), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n386_), .A2(G36gat), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n578_), .A2(KEYINPUT97), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n599_));
  INV_X1    g398(.A(new_n596_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n599_), .B1(new_n577_), .B2(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n597_), .A2(new_n598_), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n598_), .B1(new_n597_), .B2(new_n601_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n595_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n597_), .A2(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT96), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n597_), .A2(new_n598_), .A3(new_n601_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(KEYINPUT45), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n386_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n609_));
  INV_X1    g408(.A(G36gat), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n604_), .B(new_n608_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT46), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n591_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n588_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n550_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(G36gat), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n617_), .A2(KEYINPUT46), .A3(new_n604_), .A4(new_n608_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n618_), .ZN(G1329gat));
  NOR3_X1   g418(.A1(new_n577_), .A2(G43gat), .A3(new_n248_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n248_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n622_));
  INV_X1    g421(.A(G43gat), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n621_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT98), .B(KEYINPUT47), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n621_), .B(new_n625_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1330gat));
  INV_X1    g428(.A(new_n305_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G50gat), .B1(new_n578_), .B2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(G50gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n592_), .B2(new_n632_), .ZN(G1331gat));
  NAND2_X1  g432(.A1(new_n420_), .A2(new_n532_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n542_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(KEYINPUT100), .B(G57gat), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n540_), .A2(new_n368_), .A3(new_n635_), .A4(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT101), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n388_), .A2(new_n420_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n542_), .A2(new_n533_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n642_), .A2(KEYINPUT99), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(KEYINPUT99), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n368_), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n638_), .B1(new_n645_), .B2(new_n464_), .ZN(G1332gat));
  NAND2_X1  g445(.A1(new_n540_), .A2(new_n635_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G64gat), .B1(new_n647_), .B2(new_n386_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT102), .B(KEYINPUT48), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n642_), .A2(new_n462_), .A3(new_n550_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1333gat));
  OAI21_X1  g451(.A(G71gat), .B1(new_n647_), .B2(new_n248_), .ZN(new_n653_));
  XOR2_X1   g452(.A(KEYINPUT103), .B(KEYINPUT49), .Z(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n248_), .A2(G71gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n641_), .B2(new_n656_), .ZN(G1334gat));
  OAI21_X1  g456(.A(G78gat), .B1(new_n647_), .B2(new_n305_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT50), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n305_), .A2(G78gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n641_), .B2(new_n660_), .ZN(G1335gat));
  NOR2_X1   g460(.A1(new_n542_), .A2(new_n575_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n639_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n424_), .A3(new_n368_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n502_), .A2(new_n545_), .A3(new_n420_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(new_n368_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n665_), .B1(new_n668_), .B2(new_n424_), .ZN(G1336gat));
  NAND3_X1  g468(.A1(new_n664_), .A2(new_n425_), .A3(new_n550_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n667_), .A2(new_n550_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n425_), .ZN(G1337gat));
  AND4_X1   g471(.A1(new_n247_), .A2(new_n664_), .A3(new_n438_), .A4(new_n440_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT51), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(KEYINPUT104), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n448_), .B1(new_n667_), .B2(new_n247_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n673_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1338gat));
  NOR3_X1   g478(.A1(new_n663_), .A2(G106gat), .A3(new_n305_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681_));
  INV_X1    g480(.A(new_n666_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n585_), .A2(new_n630_), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n683_), .B2(G106gat), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT52), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n680_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  AOI211_X1 g485(.A(new_n305_), .B(new_n666_), .C1(new_n582_), .C2(new_n584_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT105), .B1(new_n687_), .B2(new_n439_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(new_n681_), .A3(G106gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(KEYINPUT52), .A3(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT106), .B(KEYINPUT53), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n686_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n686_), .B2(new_n690_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1339gat));
  NOR2_X1   g493(.A1(new_n403_), .A2(KEYINPUT115), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n403_), .A2(KEYINPUT115), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n405_), .ZN(new_n697_));
  OAI221_X1 g496(.A(new_n417_), .B1(new_n695_), .B2(new_n697_), .C1(new_n412_), .C2(new_n405_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n494_), .A2(new_n698_), .A3(new_n419_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n470_), .A2(new_n478_), .A3(new_n477_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT111), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT111), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n470_), .A2(new_n477_), .A3(new_n702_), .A4(new_n478_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n483_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n482_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT55), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n482_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n482_), .B2(new_n709_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n705_), .B(new_n707_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT112), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n482_), .A2(new_n709_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT110), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n482_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI22_X1  g516(.A1(new_n704_), .A2(new_n483_), .B1(new_n706_), .B2(KEYINPUT55), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n717_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n713_), .A2(KEYINPUT56), .A3(new_n491_), .A4(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n492_), .B1(new_n712_), .B2(KEYINPUT112), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT56), .B1(new_n723_), .B2(new_n720_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n699_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT58), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n518_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n699_), .B(KEYINPUT58), .C1(new_n722_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n494_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n420_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n713_), .A2(new_n491_), .A3(new_n720_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT56), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n734_), .A2(KEYINPUT114), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n733_), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n721_), .A2(KEYINPUT114), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n735_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n731_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n496_), .A2(new_n419_), .A3(new_n698_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n574_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n729_), .B1(new_n742_), .B2(KEYINPUT57), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT57), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n744_), .B(new_n574_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n545_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n518_), .B1(new_n634_), .B2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n748_), .B2(new_n634_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n542_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT108), .B(KEYINPUT54), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n751_), .B(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n747_), .A2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n550_), .A2(new_n536_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n380_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT116), .Z(new_n759_));
  NOR2_X1   g558(.A1(new_n755_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT59), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n745_), .B1(new_n743_), .B2(KEYINPUT117), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT117), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n729_), .B(new_n763_), .C1(new_n742_), .C2(KEYINPUT57), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n532_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n765_), .A2(new_n754_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n759_), .A2(KEYINPUT59), .ZN(new_n767_));
  OAI22_X1  g566(.A1(new_n760_), .A2(new_n761_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G113gat), .B1(new_n768_), .B2(new_n420_), .ZN(new_n769_));
  INV_X1    g568(.A(G113gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n760_), .A2(new_n770_), .A3(new_n421_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1340gat));
  OAI21_X1  g571(.A(G120gat), .B1(new_n768_), .B2(new_n542_), .ZN(new_n773_));
  INV_X1    g572(.A(G120gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n542_), .B2(KEYINPUT60), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n760_), .B(new_n775_), .C1(KEYINPUT60), .C2(new_n774_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1341gat));
  NOR3_X1   g576(.A1(new_n755_), .A2(new_n545_), .A3(new_n759_), .ZN(new_n778_));
  OR3_X1    g577(.A1(new_n778_), .A2(KEYINPUT118), .A3(G127gat), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n532_), .A2(G127gat), .ZN(new_n780_));
  OAI221_X1 g579(.A(new_n780_), .B1(new_n766_), .B2(new_n767_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT118), .B1(new_n778_), .B2(G127gat), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n779_), .A2(new_n781_), .A3(new_n782_), .ZN(G1342gat));
  OAI21_X1  g582(.A(G134gat), .B1(new_n768_), .B2(new_n518_), .ZN(new_n784_));
  INV_X1    g583(.A(G134gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n760_), .A2(new_n785_), .A3(new_n574_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1343gat));
  XNOR2_X1  g586(.A(new_n751_), .B(new_n752_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n746_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n381_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n756_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(new_n420_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g592(.A1(new_n791_), .A2(new_n542_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT119), .B(G148gat), .Z(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(G1345gat));
  OAI21_X1  g595(.A(KEYINPUT120), .B1(new_n791_), .B2(new_n545_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n381_), .B1(new_n788_), .B2(new_n746_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n532_), .A4(new_n756_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT61), .B(G155gat), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n797_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1346gat));
  INV_X1    g603(.A(G162gat), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n791_), .A2(new_n805_), .A3(new_n518_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n791_), .B2(new_n517_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n808_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n806_), .B1(new_n809_), .B2(new_n810_), .ZN(G1347gat));
  NOR2_X1   g610(.A1(new_n386_), .A2(new_n368_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n757_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n420_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n765_), .B2(new_n754_), .ZN(new_n815_));
  XOR2_X1   g614(.A(KEYINPUT22), .B(G169gat), .Z(new_n816_));
  OR2_X1    g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT62), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT122), .B(new_n814_), .C1(new_n765_), .C2(new_n754_), .ZN(new_n821_));
  AND4_X1   g620(.A1(new_n818_), .A2(new_n820_), .A3(G169gat), .A4(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(G169gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n818_), .B1(new_n824_), .B2(new_n821_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n817_), .B1(new_n822_), .B2(new_n825_), .ZN(G1348gat));
  INV_X1    g625(.A(new_n813_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n789_), .A2(G176gat), .A3(new_n502_), .A4(new_n827_), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT123), .Z(new_n829_));
  NOR2_X1   g628(.A1(new_n766_), .A2(new_n813_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G176gat), .B1(new_n830_), .B2(new_n502_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1349gat));
  NOR3_X1   g631(.A1(new_n755_), .A2(new_n545_), .A3(new_n813_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n833_), .A2(KEYINPUT124), .ZN(new_n834_));
  AOI21_X1  g633(.A(G183gat), .B1(new_n833_), .B2(KEYINPUT124), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n545_), .A2(new_n211_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n834_), .A2(new_n835_), .B1(new_n830_), .B2(new_n836_), .ZN(G1350gat));
  NAND2_X1  g636(.A1(new_n830_), .A2(new_n580_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G190gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n830_), .A2(new_n212_), .A3(new_n574_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1351gat));
  OAI211_X1 g640(.A(new_n790_), .B(new_n812_), .C1(new_n747_), .C2(new_n754_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n421_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n502_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g646(.A(new_n545_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT125), .B1(new_n842_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT125), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n798_), .A2(new_n851_), .A3(new_n812_), .A4(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1354gat));
  XNOR2_X1  g654(.A(KEYINPUT127), .B(G218gat), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n842_), .A2(new_n518_), .A3(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n843_), .A2(KEYINPUT126), .A3(new_n574_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n842_), .B2(new_n517_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n857_), .B1(new_n861_), .B2(new_n856_), .ZN(G1355gat));
endmodule


