//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_;
  XNOR2_X1  g000(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n204_), .A2(new_n205_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n203_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n204_), .A2(new_n205_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(new_n202_), .A3(new_n206_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n212_), .B(G15gat), .Z(new_n213_));
  INV_X1    g012(.A(G71gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G227gat), .A2(G233gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n216_), .B(KEYINPUT30), .Z(new_n217_));
  XNOR2_X1  g016(.A(new_n215_), .B(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT79), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n223_), .A2(new_n222_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT79), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n224_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT26), .B(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n237_), .B1(new_n238_), .B2(G183gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT25), .B(G183gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n236_), .B(new_n239_), .C1(new_n240_), .C2(new_n237_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n229_), .B1(G183gat), .B2(G190gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n243_));
  AOI21_X1  g042(.A(G176gat), .B1(new_n243_), .B2(KEYINPUT22), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G169gat), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n235_), .A2(new_n241_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT81), .B(G43gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT31), .ZN(new_n248_));
  INV_X1    g047(.A(G99gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n246_), .B(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n218_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n218_), .A2(new_n251_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G78gat), .B(G106gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT88), .Z(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G197gat), .B(G204gat), .Z(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT21), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G197gat), .B(G204gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT21), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G211gat), .ZN(new_n263_));
  INV_X1    g062(.A(G218gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G211gat), .A2(G218gat), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n259_), .A2(KEYINPUT87), .A3(new_n262_), .A4(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n265_), .A2(new_n266_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT87), .ZN(new_n270_));
  OAI211_X1 g069(.A(KEYINPUT21), .B(new_n258_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G141gat), .A2(G148gat), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT85), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n273_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT84), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n280_), .A2(new_n283_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n273_), .B(KEYINPUT3), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n284_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n275_), .A2(new_n276_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n282_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n272_), .B1(new_n290_), .B2(KEYINPUT29), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G228gat), .A2(G233gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n268_), .A2(new_n271_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n285_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n287_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n289_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n296_), .A2(new_n297_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n294_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n292_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n257_), .B1(new_n293_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT91), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n291_), .A2(new_n292_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n300_), .A2(new_n301_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n256_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n307_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(KEYINPUT91), .A3(new_n257_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(new_n290_), .B2(KEYINPUT29), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G22gat), .B(G50gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n311_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n298_), .A2(new_n299_), .A3(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n312_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n313_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n305_), .A2(new_n308_), .A3(new_n310_), .A4(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT89), .B1(new_n309_), .B2(new_n257_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n318_), .B1(new_n321_), .B2(new_n308_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n308_), .A2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n320_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n303_), .A2(new_n323_), .A3(new_n308_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n318_), .ZN(new_n327_));
  AND4_X1   g126(.A1(new_n320_), .A2(new_n326_), .A3(new_n324_), .A4(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n319_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G1gat), .B(G29gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G85gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT0), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G57gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n296_), .A2(new_n297_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n334_), .A2(new_n211_), .A3(new_n209_), .A4(new_n282_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n275_), .A2(new_n278_), .ZN(new_n336_));
  OR2_X1    g135(.A1(G141gat), .A2(G148gat), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n336_), .A2(new_n281_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n289_), .B1(new_n295_), .B2(new_n287_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n212_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G225gat), .A2(G233gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n335_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n333_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n335_), .A2(new_n340_), .A3(KEYINPUT4), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n290_), .A2(new_n346_), .A3(new_n212_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n341_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT97), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT97), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n345_), .A2(new_n350_), .A3(new_n341_), .A4(new_n347_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n344_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT98), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G64gat), .B(G92gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n221_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT22), .B(G169gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT93), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n361_), .B(new_n242_), .C1(new_n363_), .C2(G176gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n233_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n224_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT92), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n240_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n236_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n365_), .B(new_n366_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n272_), .A2(new_n364_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT20), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT94), .B1(new_n246_), .B2(new_n272_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n232_), .A2(new_n234_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n366_), .A3(new_n241_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n242_), .A2(new_n245_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT94), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n294_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n372_), .B1(new_n373_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT19), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n364_), .A2(new_n370_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n294_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n246_), .A2(new_n272_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(KEYINPUT20), .A4(new_n382_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n360_), .B1(new_n383_), .B2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n359_), .B(new_n387_), .C1(new_n380_), .C2(new_n382_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(KEYINPUT96), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT96), .ZN(new_n392_));
  INV_X1    g191(.A(new_n382_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n373_), .A2(new_n379_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(new_n372_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n359_), .B1(new_n395_), .B2(new_n387_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n390_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n392_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n333_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n341_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n342_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n399_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT33), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT33), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n404_), .B(new_n399_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n354_), .A2(new_n391_), .A3(new_n398_), .A4(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n383_), .B2(new_n388_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT99), .ZN(new_n410_));
  OR3_X1    g209(.A1(new_n400_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n402_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n380_), .A2(new_n393_), .ZN(new_n413_));
  AND4_X1   g212(.A1(KEYINPUT20), .A2(new_n385_), .A3(new_n393_), .A4(new_n386_), .ZN(new_n414_));
  OAI211_X1 g213(.A(KEYINPUT32), .B(new_n360_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n416_), .B(new_n408_), .C1(new_n383_), .C2(new_n388_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n410_), .A2(new_n412_), .A3(new_n415_), .A4(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n329_), .B1(new_n407_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n319_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n326_), .A2(new_n324_), .A3(new_n327_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT90), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n322_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT27), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n359_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n389_), .A2(new_n427_), .A3(KEYINPUT27), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n424_), .A2(new_n429_), .A3(new_n412_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n254_), .B1(new_n419_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n429_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n424_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n412_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n252_), .A2(new_n434_), .A3(new_n253_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n431_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT12), .ZN(new_n439_));
  INV_X1    g238(.A(G85gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(KEYINPUT9), .ZN(new_n441_));
  INV_X1    g240(.A(G92gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT65), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT65), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G92gat), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n441_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT9), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(G85gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(G92gat), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT66), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n446_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n440_), .A2(G92gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n442_), .A2(G85gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT9), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n441_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT66), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G99gat), .A2(G106gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G106gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT10), .B(G99gat), .Z(new_n463_));
  AOI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n448_), .A2(new_n449_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(new_n249_), .A3(new_n462_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n465_), .B1(new_n461_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT8), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT8), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n472_), .B(new_n465_), .C1(new_n461_), .C2(new_n469_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n458_), .A2(new_n464_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT11), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n477_), .A2(new_n478_), .A3(G78gat), .ZN(new_n479_));
  INV_X1    g278(.A(G78gat), .ZN(new_n480_));
  OR2_X1    g279(.A1(KEYINPUT67), .A2(G71gat), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n481_), .B2(new_n476_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n475_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(G78gat), .B1(new_n477_), .B2(new_n478_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n480_), .A3(new_n476_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n485_), .A3(KEYINPUT11), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G57gat), .B(G64gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n487_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n489_), .A2(new_n484_), .A3(KEYINPUT11), .A4(new_n485_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n439_), .B1(new_n474_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G230gat), .A2(G233gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT64), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n474_), .B2(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n471_), .A2(new_n473_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n451_), .B1(new_n446_), .B2(new_n450_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n455_), .A2(KEYINPUT66), .A3(new_n456_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n464_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n488_), .A2(new_n490_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT12), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n492_), .A2(new_n496_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT69), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT68), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n474_), .B2(new_n491_), .ZN(new_n508_));
  AND4_X1   g307(.A1(new_n507_), .A2(new_n491_), .A3(new_n497_), .A4(new_n500_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n501_), .A2(new_n502_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT68), .B1(new_n501_), .B2(new_n502_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n474_), .A2(new_n507_), .A3(new_n491_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT69), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n505_), .B1(new_n515_), .B2(new_n495_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G120gat), .B(G148gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT5), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(G176gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(G204gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n520_), .ZN(new_n525_));
  AOI211_X1 g324(.A(new_n525_), .B(new_n505_), .C1(new_n515_), .C2(new_n495_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT13), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n515_), .A2(new_n495_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(new_n504_), .A3(new_n520_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT13), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n529_), .B(new_n530_), .C1(new_n516_), .C2(new_n523_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G1gat), .A2(G8gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT14), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT74), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n536_), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT75), .ZN(new_n543_));
  XOR2_X1   g342(.A(G1gat), .B(G8gat), .Z(new_n544_));
  INV_X1    g343(.A(KEYINPUT75), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n539_), .A2(new_n545_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n543_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G29gat), .B(G36gat), .ZN(new_n549_));
  INV_X1    g348(.A(G50gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(G43gat), .ZN(new_n551_));
  INV_X1    g350(.A(G43gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(G50gat), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT71), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n549_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n552_), .A2(G50gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n550_), .A2(G43gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT71), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n549_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n557_), .A2(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n547_), .A2(new_n548_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n544_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n536_), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT74), .B1(new_n536_), .B2(KEYINPUT14), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n545_), .B1(new_n570_), .B2(new_n540_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n546_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n567_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n543_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n566_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n535_), .B1(new_n565_), .B2(new_n575_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n557_), .A2(KEYINPUT15), .A3(new_n563_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT15), .B1(new_n557_), .B2(new_n563_), .ZN(new_n578_));
  OAI22_X1  g377(.A1(new_n547_), .A2(new_n548_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(new_n566_), .A3(new_n574_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n534_), .B(KEYINPUT77), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G113gat), .B(G141gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n219_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(G197gat), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n576_), .A2(new_n583_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n576_), .B2(new_n583_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n533_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n438_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n491_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT76), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n547_), .A2(new_n548_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n598_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT16), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(G183gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(new_n263_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT17), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n599_), .A2(new_n609_), .A3(new_n600_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(G134gat), .ZN(new_n613_));
  INV_X1    g412(.A(G162gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT34), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n501_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(KEYINPUT72), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n474_), .A2(new_n566_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n620_), .B2(KEYINPUT72), .ZN(new_n623_));
  OAI211_X1 g422(.A(KEYINPUT35), .B(new_n619_), .C1(new_n621_), .C2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n619_), .B(KEYINPUT35), .Z(new_n625_));
  NAND3_X1  g424(.A1(new_n620_), .A2(new_n622_), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n617_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n615_), .A2(new_n616_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n624_), .A2(new_n616_), .A3(new_n615_), .A4(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT73), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT37), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n629_), .A2(new_n630_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n611_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n593_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT100), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n640_), .A2(G1gat), .A3(new_n434_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT101), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n631_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n611_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n593_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n434_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT38), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n642_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n641_), .A2(new_n651_), .A3(KEYINPUT38), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n644_), .A2(new_n650_), .A3(new_n652_), .ZN(G1324gat));
  OAI21_X1  g452(.A(G8gat), .B1(new_n647_), .B2(new_n432_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT39), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n432_), .A2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n640_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  NOR3_X1   g458(.A1(new_n640_), .A2(G15gat), .A3(new_n254_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(KEYINPUT104), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(KEYINPUT104), .ZN(new_n662_));
  OAI21_X1  g461(.A(G15gat), .B1(new_n647_), .B2(new_n254_), .ZN(new_n663_));
  XOR2_X1   g462(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT41), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n663_), .B(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(new_n662_), .A3(new_n666_), .ZN(G1326gat));
  OAI21_X1  g466(.A(G22gat), .B1(new_n647_), .B2(new_n424_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n424_), .A2(G22gat), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT106), .Z(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n640_), .B2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(new_n611_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n631_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n593_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(G29gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n412_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT44), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n635_), .A2(new_n637_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT43), .B(new_n682_), .C1(new_n431_), .C2(new_n437_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n629_), .A2(new_n630_), .A3(new_n636_), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n629_), .A2(new_n630_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(KEYINPUT107), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n431_), .B2(new_n437_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT108), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n684_), .A2(new_n685_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n687_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n682_), .A2(KEYINPUT107), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n252_), .A2(new_n253_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n398_), .A2(new_n391_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n349_), .A2(new_n351_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n344_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n353_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AOI211_X1 g500(.A(KEYINPUT98), .B(new_n344_), .C1(new_n349_), .C2(new_n351_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n406_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n418_), .B1(new_n698_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n424_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n329_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n697_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n696_), .B1(new_n707_), .B2(new_n436_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(KEYINPUT43), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n683_), .B1(new_n692_), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n592_), .B1(new_n679_), .B2(KEYINPUT44), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(new_n674_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n681_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n683_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n708_), .A2(new_n709_), .A3(KEYINPUT43), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n709_), .B1(new_n708_), .B2(KEYINPUT43), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n680_), .A3(new_n713_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n434_), .B1(new_n715_), .B2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n678_), .B1(new_n721_), .B2(new_n677_), .ZN(G1328gat));
  INV_X1    g521(.A(G36gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n676_), .A2(new_n723_), .A3(new_n429_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT45), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n432_), .B1(new_n715_), .B2(new_n720_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n723_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n725_), .B(KEYINPUT46), .C1(new_n723_), .C2(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1329gat));
  NAND3_X1  g530(.A1(new_n676_), .A2(new_n552_), .A3(new_n697_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n254_), .B1(new_n715_), .B2(new_n720_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n552_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n734_), .B(new_n736_), .ZN(G1330gat));
  NAND3_X1  g536(.A1(new_n676_), .A2(new_n550_), .A3(new_n329_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n715_), .A2(new_n720_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n329_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n740_), .A2(KEYINPUT111), .A3(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT111), .B1(new_n740_), .B2(G50gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(G1331gat));
  INV_X1    g542(.A(new_n591_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n532_), .A2(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n438_), .A2(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(new_n638_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G57gat), .B1(new_n747_), .B2(new_n412_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n646_), .ZN(new_n749_));
  INV_X1    g548(.A(G57gat), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n434_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1332gat));
  OAI21_X1  g551(.A(G64gat), .B1(new_n749_), .B2(new_n432_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT48), .ZN(new_n754_));
  INV_X1    g553(.A(G64gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n747_), .A2(new_n755_), .A3(new_n429_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1333gat));
  OAI21_X1  g556(.A(G71gat), .B1(new_n749_), .B2(new_n254_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT49), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n747_), .A2(new_n214_), .A3(new_n697_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1334gat));
  OAI21_X1  g560(.A(G78gat), .B1(new_n749_), .B2(new_n424_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT50), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n747_), .A2(new_n480_), .A3(new_n329_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1335gat));
  NAND2_X1  g564(.A1(new_n746_), .A2(new_n675_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT112), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n746_), .A2(new_n768_), .A3(new_n675_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G85gat), .B1(new_n770_), .B2(new_n412_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(KEYINPUT113), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n771_), .A2(KEYINPUT113), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n719_), .A2(new_n611_), .A3(new_n745_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n434_), .A2(new_n440_), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n772_), .B(new_n773_), .C1(new_n774_), .C2(new_n775_), .ZN(G1336gat));
  AOI21_X1  g575(.A(G92gat), .B1(new_n770_), .B2(new_n429_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n429_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n774_), .B2(new_n778_), .ZN(G1337gat));
  AOI21_X1  g578(.A(new_n249_), .B1(new_n774_), .B2(new_n697_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n770_), .A2(new_n463_), .A3(new_n697_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT114), .ZN(new_n782_));
  OR3_X1    g581(.A1(new_n780_), .A2(new_n782_), .A3(KEYINPUT51), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT51), .B1(new_n780_), .B2(new_n782_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1338gat));
  NAND3_X1  g584(.A1(new_n770_), .A2(new_n462_), .A3(new_n329_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n719_), .A2(new_n329_), .A3(new_n611_), .A4(new_n745_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n787_), .A2(new_n788_), .A3(G106gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n787_), .B2(G106gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n793_), .B(new_n786_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n508_), .A2(new_n509_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n492_), .A2(new_n503_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n495_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n504_), .A2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n492_), .A2(new_n496_), .A3(KEYINPUT55), .A4(new_n503_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n801_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n798_), .B(KEYINPUT56), .C1(new_n805_), .C2(new_n522_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n582_), .B1(new_n565_), .B2(new_n575_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n586_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n588_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT116), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n588_), .A2(new_n809_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n529_), .A2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n806_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n805_), .A2(new_n522_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n522_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n798_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT58), .B1(new_n816_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n797_), .B1(new_n822_), .B2(new_n682_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n816_), .A2(KEYINPUT58), .A3(new_n821_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n522_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n522_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n826_), .A2(new_n827_), .A3(KEYINPUT118), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n817_), .A2(KEYINPUT118), .A3(new_n818_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n516_), .A2(new_n520_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n825_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n693_), .A3(KEYINPUT119), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n823_), .A2(new_n824_), .A3(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n814_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n744_), .B(new_n529_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n814_), .C1(new_n524_), .C2(new_n526_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n631_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(KEYINPUT57), .A3(new_n631_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n840_), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n631_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n834_), .A2(new_n843_), .A3(new_n846_), .A4(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n611_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n674_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n532_), .A2(new_n591_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT115), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n638_), .A2(new_n853_), .A3(new_n591_), .A4(new_n532_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n852_), .A2(KEYINPUT54), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT54), .B1(new_n852_), .B2(new_n854_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n849_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n433_), .A2(new_n434_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n697_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT59), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n858_), .A2(new_n862_), .A3(new_n697_), .A4(new_n859_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n744_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G113gat), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n591_), .A2(G113gat), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n860_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n796_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  AOI211_X1 g668(.A(KEYINPUT121), .B(new_n867_), .C1(new_n864_), .C2(G113gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1340gat));
  INV_X1    g670(.A(new_n860_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT122), .B(G120gat), .Z(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n532_), .B2(KEYINPUT60), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(KEYINPUT60), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(KEYINPUT123), .B2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n872_), .B(new_n876_), .C1(KEYINPUT123), .C2(new_n874_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n861_), .A2(new_n863_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n532_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n877_), .B1(new_n879_), .B2(new_n873_), .ZN(G1341gat));
  NAND2_X1  g679(.A1(new_n674_), .A2(G127gat), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n860_), .A2(new_n611_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(G127gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT124), .B1(new_n882_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886_));
  OAI221_X1 g685(.A(new_n886_), .B1(G127gat), .B2(new_n883_), .C1(new_n878_), .C2(new_n881_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1342gat));
  AOI21_X1  g687(.A(G134gat), .B1(new_n872_), .B2(new_n645_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n878_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n693_), .A2(G134gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(G1343gat));
  NAND3_X1  g691(.A1(new_n858_), .A2(new_n329_), .A3(new_n432_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n893_), .A2(new_n434_), .A3(new_n697_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n744_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n533_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n674_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1346gat));
  AOI21_X1  g700(.A(G162gat), .B1(new_n894_), .B2(new_n645_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n689_), .A2(new_n614_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n894_), .B2(new_n903_), .ZN(G1347gat));
  AOI21_X1  g703(.A(new_n412_), .B1(new_n849_), .B2(new_n857_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n254_), .A2(new_n329_), .A3(new_n432_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n744_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G169gat), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n912_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n909_), .A2(G169gat), .A3(new_n914_), .A4(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n913_), .B(new_n916_), .C1(new_n363_), .C2(new_n909_), .ZN(G1348gat));
  NOR2_X1   g716(.A1(new_n907_), .A2(new_n532_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n220_), .ZN(G1349gat));
  NAND2_X1  g718(.A1(new_n908_), .A2(new_n674_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G183gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(new_n920_), .B2(new_n368_), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n908_), .A2(new_n236_), .A3(new_n645_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G190gat), .B1(new_n907_), .B2(new_n682_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1351gat));
  NOR2_X1   g724(.A1(new_n424_), .A2(new_n432_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n905_), .A2(new_n254_), .A3(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n744_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n533_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n263_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n928_), .A2(new_n674_), .A3(new_n934_), .A4(new_n935_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n933_), .B(new_n263_), .C1(new_n927_), .C2(new_n611_), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n936_), .B2(new_n938_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1354gat));
  NOR3_X1   g740(.A1(new_n927_), .A2(new_n264_), .A3(new_n682_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n928_), .A2(new_n645_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n264_), .B2(new_n943_), .ZN(G1355gat));
endmodule


