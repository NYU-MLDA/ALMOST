//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n962_, new_n963_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n996_, new_n997_, new_n998_;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(KEYINPUT84), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211_));
  NOR3_X1   g010(.A1(new_n211_), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT85), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(KEYINPUT84), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n211_), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .A4(new_n208_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT82), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT82), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n219_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT86), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT86), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n227_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n224_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n207_), .B1(new_n218_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n222_), .A2(KEYINPUT82), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n220_), .A2(G141gat), .A3(G148gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n209_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n204_), .B1(new_n206_), .B2(KEYINPUT1), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n240_), .B2(KEYINPUT83), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT83), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n242_), .B(new_n204_), .C1(new_n206_), .C2(KEYINPUT1), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n238_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AND4_X1   g044(.A1(new_n203_), .A2(new_n232_), .A3(new_n233_), .A4(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n230_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(new_n236_), .B2(new_n219_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n248_), .A2(new_n213_), .A3(new_n229_), .A4(new_n217_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n244_), .B1(new_n249_), .B2(new_n207_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n203_), .B1(new_n250_), .B2(new_n233_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G22gat), .B(G50gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n246_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n232_), .A2(new_n233_), .A3(new_n245_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT28), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n203_), .A3(new_n233_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n202_), .B1(new_n254_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n253_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(new_n257_), .A3(new_n252_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT88), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G228gat), .A2(G233gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n233_), .B1(new_n232_), .B2(new_n245_), .ZN(new_n268_));
  INV_X1    g067(.A(G197gat), .ZN(new_n269_));
  INV_X1    g068(.A(G204gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G197gat), .A2(G204gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT21), .A3(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT21), .ZN(new_n276_));
  INV_X1    g075(.A(new_n272_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G197gat), .A2(G204gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n265_), .B2(new_n264_), .ZN(new_n282_));
  OAI21_X1  g081(.A(G78gat), .B1(new_n268_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n282_), .ZN(new_n284_));
  INV_X1    g083(.A(G78gat), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n284_), .B(new_n285_), .C1(new_n250_), .C2(new_n233_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n283_), .A2(G106gat), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(G106gat), .B1(new_n283_), .B2(new_n286_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n267_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n283_), .A2(new_n286_), .ZN(new_n290_));
  INV_X1    g089(.A(G106gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n283_), .A2(G106gat), .A3(new_n286_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n266_), .A3(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n263_), .B1(new_n289_), .B2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT88), .B1(new_n260_), .B2(new_n261_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n289_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT98), .ZN(new_n299_));
  INV_X1    g098(.A(G134gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G127gat), .ZN(new_n301_));
  INV_X1    g100(.A(G127gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G134gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G120gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G113gat), .ZN(new_n306_));
  INV_X1    g105(.A(G113gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G120gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n301_), .A2(new_n303_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AOI211_X1 g112(.A(new_n313_), .B(new_n244_), .C1(new_n249_), .C2(new_n207_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT80), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n315_), .A3(new_n311_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n304_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n317_), .A2(KEYINPUT80), .A3(new_n306_), .A4(new_n308_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n232_), .B2(new_n245_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT4), .B1(new_n314_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n232_), .A2(new_n245_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n319_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n321_), .A2(new_n323_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G1gat), .B(G29gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G57gat), .B(G85gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n232_), .A2(new_n245_), .A3(new_n312_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n323_), .B1(new_n326_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n329_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n329_), .B2(new_n338_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n299_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n329_), .A2(new_n338_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n334_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n329_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(KEYINPUT98), .A3(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G8gat), .B(G36gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT18), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n352_));
  AND2_X1   g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT90), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G183gat), .ZN(new_n357_));
  INV_X1    g156(.A(G190gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT23), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(G183gat), .A3(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(KEYINPUT25), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G183gat), .ZN(new_n365_));
  AND2_X1   g164(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n363_), .B(new_n365_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT24), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT91), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT24), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n373_), .B2(KEYINPUT24), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n369_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT92), .B1(new_n372_), .B2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n376_), .A2(new_n369_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n375_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n359_), .A2(new_n361_), .B1(new_n370_), .B2(new_n369_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT92), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .A4(new_n368_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n378_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n357_), .A2(new_n358_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n362_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G169gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT22), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT22), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G169gat), .ZN(new_n391_));
  INV_X1    g190(.A(G176gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n387_), .A2(new_n373_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n385_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n281_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT20), .ZN(new_n397_));
  INV_X1    g196(.A(new_n369_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT24), .A3(new_n373_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n362_), .A2(new_n399_), .A3(new_n371_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n363_), .A2(new_n365_), .ZN(new_n401_));
  AND2_X1   g200(.A1(KEYINPUT77), .A2(G190gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(KEYINPUT77), .A2(G190gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT26), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n367_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n401_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n400_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n403_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(KEYINPUT77), .A2(G190gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n357_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n362_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT79), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT78), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n393_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT22), .B(G169gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(KEYINPUT78), .A3(new_n392_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n411_), .A2(new_n412_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n402_), .A2(new_n403_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n418_), .A2(new_n357_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n419_), .A2(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n407_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n275_), .A2(new_n280_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n397_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n356_), .B1(new_n396_), .B2(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n385_), .A2(new_n422_), .A3(new_n394_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n417_), .A2(new_n420_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n404_), .A2(new_n405_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n382_), .B(new_n399_), .C1(new_n427_), .C2(new_n401_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n422_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n354_), .A2(new_n397_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n425_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n351_), .B1(new_n424_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT78), .B1(new_n415_), .B2(new_n392_), .ZN(new_n435_));
  AND4_X1   g234(.A1(KEYINPUT78), .A2(new_n389_), .A3(new_n391_), .A4(new_n392_), .ZN(new_n436_));
  OAI22_X1  g235(.A1(new_n419_), .A2(KEYINPUT79), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n373_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n428_), .B(new_n422_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT20), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n422_), .B1(new_n385_), .B2(new_n394_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n355_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n385_), .A2(new_n422_), .A3(new_n394_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(new_n430_), .C1(new_n422_), .C2(new_n421_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n444_), .A3(new_n350_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n433_), .A2(new_n434_), .A3(new_n445_), .ZN(new_n446_));
  AOI211_X1 g245(.A(new_n434_), .B(new_n350_), .C1(new_n442_), .C2(new_n444_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT27), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n396_), .A2(new_n423_), .A3(new_n356_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n422_), .B(new_n394_), .C1(new_n377_), .C2(new_n372_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT20), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n354_), .B1(new_n453_), .B2(new_n429_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n351_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(KEYINPUT27), .A3(new_n445_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n450_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n298_), .B1(new_n346_), .B2(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n260_), .A2(KEYINPUT88), .A3(new_n261_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(new_n296_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n287_), .A2(new_n288_), .A3(new_n267_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n266_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n289_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n455_), .A2(KEYINPUT32), .A3(new_n350_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n350_), .A2(KEYINPUT32), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n442_), .A2(new_n444_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT97), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n442_), .A2(new_n444_), .A3(KEYINPUT97), .A4(new_n468_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n467_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n343_), .A2(new_n344_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT95), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n476_), .B1(new_n340_), .B2(KEYINPUT33), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT4), .B1(new_n324_), .B2(new_n325_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n336_), .B1(new_n250_), .B2(new_n319_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n480_), .B2(KEYINPUT4), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n337_), .B1(new_n481_), .B2(new_n323_), .ZN(new_n482_));
  OAI211_X1 g281(.A(KEYINPUT95), .B(new_n478_), .C1(new_n482_), .C2(new_n335_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n340_), .A2(KEYINPUT33), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n323_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n480_), .A2(new_n486_), .ZN(new_n489_));
  OAI221_X1 g288(.A(new_n335_), .B1(new_n481_), .B2(new_n323_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n445_), .A2(new_n434_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n350_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n485_), .B(new_n490_), .C1(new_n493_), .C2(new_n447_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n466_), .B(new_n475_), .C1(new_n484_), .C2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n319_), .B(KEYINPUT31), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G227gat), .A2(G233gat), .ZN(new_n497_));
  INV_X1    g296(.A(G15gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT30), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G71gat), .B(G99gat), .ZN(new_n502_));
  INV_X1    g301(.A(G43gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n421_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n421_), .A2(new_n505_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n501_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(new_n500_), .A3(new_n506_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT81), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n496_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n513_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n509_), .A2(new_n511_), .A3(KEYINPUT81), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n514_), .B1(new_n517_), .B2(new_n496_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n459_), .A2(new_n495_), .A3(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n298_), .A2(new_n458_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n346_), .A2(new_n518_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT13), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n525_));
  INV_X1    g324(.A(G85gat), .ZN(new_n526_));
  INV_X1    g325(.A(G92gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT64), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n528_), .B(new_n529_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n530_), .A2(new_n531_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT6), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT6), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(G99gat), .A3(G106gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT10), .B(G99gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n539_), .B1(new_n540_), .B2(G106gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT65), .B1(new_n534_), .B2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n545_), .A2(new_n291_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT65), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n546_), .B(new_n547_), .C1(new_n533_), .C2(new_n532_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n542_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n528_), .A2(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n536_), .A2(new_n538_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553_));
  INV_X1    g352(.A(G99gat), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n291_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n551_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT8), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT8), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n560_), .B(new_n551_), .C1(new_n552_), .C2(new_n557_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n549_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G57gat), .B(G64gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT11), .ZN(new_n565_));
  XOR2_X1   g364(.A(G71gat), .B(G78gat), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n564_), .A2(KEYINPUT11), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n565_), .A2(new_n566_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n525_), .B1(new_n563_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n563_), .A2(new_n571_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n542_), .A2(new_n548_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n570_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(KEYINPUT66), .A3(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n573_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT67), .B(KEYINPUT12), .Z(new_n581_));
  NAND2_X1  g380(.A1(new_n573_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT67), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n563_), .B(new_n571_), .C1(new_n583_), .C2(KEYINPUT12), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n579_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n582_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G120gat), .B(G148gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT5), .ZN(new_n588_));
  XOR2_X1   g387(.A(G176gat), .B(G204gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT68), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n580_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n580_), .B2(new_n586_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n524_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n580_), .A2(new_n586_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n591_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n580_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(KEYINPUT13), .A3(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n594_), .A2(new_n599_), .A3(KEYINPUT69), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT69), .B1(new_n594_), .B2(new_n599_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(G36gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(G29gat), .ZN(new_n604_));
  INV_X1    g403(.A(G29gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G36gat), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(G50gat), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(G43gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n503_), .A2(G50gat), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n604_), .A2(new_n606_), .A3(new_n609_), .A4(new_n610_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT75), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G1gat), .B(G8gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT73), .ZN(new_n617_));
  INV_X1    g416(.A(G22gat), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n498_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G15gat), .A2(G22gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G1gat), .A2(G8gat), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n619_), .A2(new_n620_), .B1(KEYINPUT14), .B2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n617_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n615_), .B(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G229gat), .A2(G233gat), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n615_), .A2(new_n623_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n612_), .A2(new_n613_), .A3(KEYINPUT15), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT15), .B1(new_n612_), .B2(new_n613_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n623_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n628_), .A2(new_n625_), .A3(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G113gat), .B(G141gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G169gat), .B(G197gat), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n634_), .B(new_n635_), .Z(new_n636_));
  NAND3_X1  g435(.A1(new_n627_), .A2(new_n633_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT76), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n627_), .A2(new_n633_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(new_n636_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n602_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n523_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT37), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT72), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(KEYINPUT72), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT71), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT70), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n549_), .A2(new_n562_), .A3(new_n614_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n631_), .B1(new_n549_), .B2(new_n562_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n549_), .A2(new_n562_), .A3(new_n614_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT35), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n654_), .B(new_n655_), .C1(new_n631_), .C2(new_n574_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n657_));
  NAND2_X1  g456(.A1(G232gat), .A2(G233gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n653_), .A2(new_n656_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n659_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n650_), .B(new_n661_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n649_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(G190gat), .B(G218gat), .Z(new_n664_));
  XNOR2_X1  g463(.A(G134gat), .B(G162gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT36), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n667_), .A2(KEYINPUT36), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n663_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n670_), .ZN(new_n672_));
  AOI221_X4 g471(.A(new_n649_), .B1(new_n672_), .B2(new_n668_), .C1(new_n660_), .C2(new_n662_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n647_), .B(new_n648_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n669_), .A2(new_n670_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n663_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n673_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n677_), .A2(KEYINPUT72), .A3(new_n646_), .A4(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(G231gat), .A2(G233gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n575_), .B(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n623_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(G127gat), .B(G155gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT16), .ZN(new_n686_));
  XOR2_X1   g485(.A(G183gat), .B(G211gat), .Z(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n684_), .A2(KEYINPUT17), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT74), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n684_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(KEYINPUT17), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n693_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n690_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n680_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n645_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n346_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n698_), .A2(G1gat), .A3(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT38), .ZN(new_n701_));
  INV_X1    g500(.A(new_n518_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n477_), .A2(new_n483_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n446_), .A2(new_n448_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n485_), .A4(new_n490_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n464_), .A2(new_n465_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  AOI22_X1  g506(.A1(new_n707_), .A2(new_n459_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n671_), .A2(new_n673_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n696_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n644_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n346_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n700_), .B1(G1gat), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT38), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n701_), .B1(new_n716_), .B2(new_n717_), .ZN(G1324gat));
  INV_X1    g517(.A(new_n698_), .ZN(new_n719_));
  INV_X1    g518(.A(G8gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n458_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n458_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n713_), .A2(new_n722_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n723_), .A2(KEYINPUT99), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT39), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n720_), .B1(new_n723_), .B2(KEYINPUT99), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n721_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT40), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(KEYINPUT40), .B(new_n721_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1325gat));
  AOI21_X1  g532(.A(new_n498_), .B1(new_n714_), .B2(new_n702_), .ZN(new_n734_));
  XOR2_X1   g533(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n735_));
  OR2_X1    g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n719_), .A2(new_n498_), .A3(new_n702_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n735_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(G1326gat));
  XNOR2_X1  g538(.A(new_n298_), .B(KEYINPUT101), .ZN(new_n740_));
  OAI21_X1  g539(.A(G22gat), .B1(new_n713_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT42), .ZN(new_n742_));
  INV_X1    g541(.A(new_n740_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n719_), .A2(new_n618_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT102), .Z(G1327gat));
  NOR2_X1   g545(.A1(new_n712_), .A2(new_n709_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n645_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G29gat), .B1(new_n749_), .B2(new_n346_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n696_), .B(new_n642_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT103), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n674_), .A2(new_n679_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT43), .B1(new_n708_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n523_), .A2(new_n755_), .A3(new_n680_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n752_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT105), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n751_), .B(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n755_), .B1(new_n523_), .B2(new_n680_), .ZN(new_n762_));
  AOI211_X1 g561(.A(KEYINPUT43), .B(new_n753_), .C1(new_n519_), .C2(new_n522_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n765_));
  INV_X1    g564(.A(new_n758_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n757_), .A2(KEYINPUT44), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n759_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n699_), .A2(new_n605_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n750_), .B1(new_n770_), .B2(new_n771_), .ZN(G1328gat));
  NOR3_X1   g571(.A1(new_n748_), .A2(G36gat), .A3(new_n722_), .ZN(new_n773_));
  XOR2_X1   g572(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT108), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n773_), .B(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n759_), .A2(new_n767_), .A3(new_n458_), .A4(new_n768_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT106), .ZN(new_n778_));
  OAI21_X1  g577(.A(G36gat), .B1(new_n777_), .B2(KEYINPUT106), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(KEYINPUT46), .B(new_n776_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1329gat));
  OAI21_X1  g583(.A(G43gat), .B1(new_n769_), .B2(new_n518_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n749_), .A2(new_n503_), .A3(new_n702_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(G1330gat));
  AOI21_X1  g588(.A(G50gat), .B1(new_n749_), .B2(new_n743_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n466_), .A2(new_n608_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n770_), .B2(new_n791_), .ZN(G1331gat));
  INV_X1    g591(.A(new_n602_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n708_), .A2(new_n642_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n697_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(G57gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n346_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n793_), .A2(new_n642_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n711_), .A2(new_n712_), .A3(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(new_n346_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n798_), .B1(new_n801_), .B2(new_n797_), .ZN(G1332gat));
  INV_X1    g601(.A(G64gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n800_), .B2(new_n458_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n796_), .A2(new_n803_), .A3(new_n458_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1333gat));
  INV_X1    g607(.A(G71gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n800_), .B2(new_n702_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n702_), .A2(new_n809_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n795_), .B2(new_n813_), .ZN(G1334gat));
  AOI21_X1  g613(.A(new_n285_), .B1(new_n800_), .B2(new_n743_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT50), .Z(new_n816_));
  NAND3_X1  g615(.A1(new_n796_), .A2(new_n285_), .A3(new_n743_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(G1335gat));
  NAND2_X1  g617(.A1(new_n794_), .A2(new_n747_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n526_), .B1(new_n819_), .B2(new_n699_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT111), .Z(new_n821_));
  NAND2_X1  g620(.A1(new_n799_), .A2(new_n696_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n346_), .A2(G85gat), .ZN(new_n824_));
  XOR2_X1   g623(.A(new_n824_), .B(KEYINPUT112), .Z(new_n825_));
  AOI21_X1  g624(.A(new_n821_), .B1(new_n823_), .B2(new_n825_), .ZN(G1336gat));
  AND2_X1   g625(.A1(new_n823_), .A2(new_n458_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n458_), .A2(new_n527_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n827_), .A2(new_n527_), .B1(new_n819_), .B2(new_n828_), .ZN(G1337gat));
  AND2_X1   g628(.A1(new_n823_), .A2(new_n702_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n702_), .A2(new_n545_), .ZN(new_n831_));
  OAI22_X1  g630(.A1(new_n830_), .A2(new_n554_), .B1(new_n819_), .B2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g632(.A1(new_n794_), .A2(new_n291_), .A3(new_n298_), .A4(new_n747_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n823_), .A2(new_n298_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G106gat), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT113), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n838_), .A3(G106gat), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n837_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n834_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT53), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n845_), .B(new_n834_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1339gat));
  NAND4_X1  g646(.A1(new_n697_), .A2(new_n643_), .A3(new_n599_), .A4(new_n594_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n586_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n586_), .B2(new_n852_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n586_), .A2(new_n852_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n582_), .A2(new_n572_), .A3(new_n584_), .A4(new_n576_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n579_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .A4(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n590_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n858_), .A2(KEYINPUT56), .A3(new_n590_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n859_), .A2(KEYINPUT118), .A3(new_n860_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n628_), .A2(new_n626_), .A3(new_n632_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n624_), .A2(new_n625_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n867_), .A2(new_n636_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n639_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n595_), .A2(new_n590_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n864_), .A2(new_n865_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n864_), .A2(KEYINPUT58), .A3(new_n871_), .A4(new_n865_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n680_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT119), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n869_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n858_), .B2(new_n590_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n860_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n863_), .A2(KEYINPUT117), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n860_), .A2(KEYINPUT117), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n882_), .B(new_n883_), .C1(new_n881_), .C2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n642_), .B1(new_n595_), .B2(new_n590_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n879_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n878_), .B1(new_n888_), .B2(new_n710_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n882_), .A2(new_n883_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n881_), .A2(new_n884_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n886_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT57), .B(new_n709_), .C1(new_n892_), .C2(new_n879_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n874_), .A2(new_n894_), .A3(new_n680_), .A4(new_n875_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n877_), .A2(new_n889_), .A3(new_n893_), .A4(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n850_), .B1(new_n896_), .B2(new_n696_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n520_), .A2(new_n346_), .A3(new_n702_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT59), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n893_), .A2(new_n889_), .A3(new_n876_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n696_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n850_), .B1(new_n901_), .B2(KEYINPUT120), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n900_), .A2(new_n903_), .A3(new_n696_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n902_), .A2(new_n904_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n898_), .A2(KEYINPUT59), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n642_), .B(new_n899_), .C1(new_n905_), .C2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G113gat), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n897_), .A2(new_n898_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n307_), .A3(new_n642_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1340gat));
  OAI211_X1 g710(.A(new_n602_), .B(new_n899_), .C1(new_n905_), .C2(new_n906_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G120gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n305_), .B1(new_n793_), .B2(KEYINPUT60), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n909_), .B(new_n914_), .C1(KEYINPUT60), .C2(new_n305_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1341gat));
  OAI211_X1 g715(.A(new_n712_), .B(new_n899_), .C1(new_n905_), .C2(new_n906_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G127gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n909_), .A2(new_n302_), .A3(new_n712_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1342gat));
  OAI211_X1 g719(.A(new_n680_), .B(new_n899_), .C1(new_n905_), .C2(new_n906_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(G134gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n909_), .A2(new_n300_), .A3(new_n710_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1343gat));
  NOR2_X1   g723(.A1(new_n702_), .A2(new_n466_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n925_), .A2(new_n346_), .A3(new_n722_), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT121), .Z(new_n927_));
  NOR2_X1   g726(.A1(new_n897_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n642_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n602_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g731(.A1(new_n928_), .A2(new_n712_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT61), .B(G155gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1346gat));
  AOI21_X1  g734(.A(G162gat), .B1(new_n928_), .B2(new_n710_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n680_), .A2(G162gat), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT122), .Z(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n928_), .B2(new_n938_), .ZN(G1347gat));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n521_), .A2(new_n458_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n743_), .A2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  AOI211_X1 g742(.A(new_n643_), .B(new_n943_), .C1(new_n902_), .C2(new_n904_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n940_), .B1(new_n944_), .B2(new_n388_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n902_), .A2(new_n904_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n942_), .ZN(new_n947_));
  OAI211_X1 g746(.A(KEYINPUT62), .B(G169gat), .C1(new_n947_), .C2(new_n643_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n944_), .A2(new_n415_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n945_), .A2(new_n948_), .A3(new_n949_), .ZN(G1348gat));
  AOI21_X1  g749(.A(new_n943_), .B1(new_n902_), .B2(new_n904_), .ZN(new_n951_));
  AOI21_X1  g750(.A(G176gat), .B1(new_n951_), .B2(new_n602_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n897_), .A2(new_n298_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n793_), .A2(new_n392_), .A3(new_n941_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n952_), .B1(new_n953_), .B2(new_n954_), .ZN(G1349gat));
  AND3_X1   g754(.A1(new_n951_), .A2(new_n401_), .A3(new_n712_), .ZN(new_n956_));
  NOR4_X1   g755(.A1(new_n897_), .A2(new_n298_), .A3(new_n696_), .A4(new_n941_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n958_));
  OR2_X1    g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(G183gat), .B1(new_n957_), .B2(new_n958_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n956_), .B1(new_n959_), .B2(new_n960_), .ZN(G1350gat));
  OAI21_X1  g760(.A(G190gat), .B1(new_n947_), .B2(new_n753_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n710_), .B1(new_n367_), .B2(new_n366_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n962_), .B1(new_n947_), .B2(new_n963_), .ZN(G1351gat));
  XNOR2_X1  g763(.A(KEYINPUT126), .B(G197gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n896_), .A2(new_n696_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n850_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n925_), .A2(new_n699_), .ZN(new_n969_));
  OR2_X1    g768(.A1(new_n969_), .A2(KEYINPUT124), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(KEYINPUT124), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n970_), .A2(new_n458_), .A3(new_n971_), .ZN(new_n972_));
  INV_X1    g771(.A(new_n972_), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n968_), .A2(KEYINPUT125), .A3(new_n973_), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n975_), .B1(new_n897_), .B2(new_n972_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n974_), .A2(new_n976_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n965_), .B1(new_n977_), .B2(new_n642_), .ZN(new_n978_));
  AND2_X1   g777(.A1(new_n269_), .A2(KEYINPUT126), .ZN(new_n979_));
  AOI211_X1 g778(.A(new_n643_), .B(new_n979_), .C1(new_n974_), .C2(new_n976_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n978_), .A2(new_n980_), .ZN(G1352gat));
  AOI21_X1  g780(.A(KEYINPUT125), .B1(new_n968_), .B2(new_n973_), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n897_), .A2(new_n975_), .A3(new_n972_), .ZN(new_n983_));
  OAI21_X1  g782(.A(new_n602_), .B1(new_n982_), .B2(new_n983_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n984_), .A2(G204gat), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n977_), .A2(new_n270_), .A3(new_n602_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n985_), .A2(new_n986_), .ZN(G1353gat));
  NOR2_X1   g786(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(KEYINPUT127), .ZN(new_n989_));
  AOI21_X1  g788(.A(new_n696_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n989_), .B1(new_n977_), .B2(new_n990_), .ZN(new_n991_));
  INV_X1    g790(.A(new_n989_), .ZN(new_n992_));
  INV_X1    g791(.A(new_n990_), .ZN(new_n993_));
  AOI211_X1 g792(.A(new_n992_), .B(new_n993_), .C1(new_n974_), .C2(new_n976_), .ZN(new_n994_));
  NOR2_X1   g793(.A1(new_n991_), .A2(new_n994_), .ZN(G1354gat));
  INV_X1    g794(.A(G218gat), .ZN(new_n996_));
  NAND3_X1  g795(.A1(new_n977_), .A2(new_n996_), .A3(new_n710_), .ZN(new_n997_));
  AOI21_X1  g796(.A(new_n753_), .B1(new_n974_), .B2(new_n976_), .ZN(new_n998_));
  OAI21_X1  g797(.A(new_n997_), .B1(new_n996_), .B2(new_n998_), .ZN(G1355gat));
endmodule


