//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n952_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT86), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n202_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n204_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT96), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT88), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n216_));
  OR2_X1    g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n212_), .A2(KEYINPUT88), .A3(KEYINPUT1), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n226_), .A2(new_n228_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n217_), .A2(new_n212_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n224_), .A2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n210_), .B1(new_n211_), .B2(new_n234_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n219_), .A2(new_n223_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n205_), .A2(new_n209_), .A3(new_n236_), .A4(KEYINPUT96), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(KEYINPUT4), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G225gat), .A2(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n210_), .A2(new_n241_), .A3(new_n234_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n235_), .A2(new_n239_), .A3(new_n237_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G57gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n243_), .A2(new_n251_), .A3(new_n244_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT98), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT98), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n255_), .A3(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G176gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT85), .ZN(new_n259_));
  INV_X1    g058(.A(G169gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(KEYINPUT22), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT22), .B(G169gat), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n258_), .B(new_n261_), .C1(new_n262_), .C2(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT23), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(new_n265_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n263_), .B(new_n264_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT25), .B(G183gat), .ZN(new_n273_));
  INV_X1    g072(.A(G190gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT81), .B1(new_n274_), .B2(KEYINPUT26), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G190gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT81), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT82), .B1(new_n276_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G183gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT25), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT25), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G183gat), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n275_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT82), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT81), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n277_), .A2(G190gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n287_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n260_), .A3(new_n258_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT83), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(KEYINPUT23), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n266_), .A2(KEYINPUT83), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n265_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n265_), .A2(KEYINPUT23), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n295_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n281_), .A2(new_n292_), .B1(new_n302_), .B2(KEYINPUT84), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n266_), .A2(KEYINPUT83), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n296_), .A2(KEYINPUT23), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n304_), .A2(new_n305_), .B1(G183gat), .B2(G190gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n294_), .B1(new_n306_), .B2(new_n300_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT84), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n260_), .A2(new_n258_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n293_), .B1(G169gat), .B2(G176gat), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n307_), .A2(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n272_), .B1(new_n303_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G71gat), .B(G99gat), .ZN(new_n313_));
  INV_X1    g112(.A(G43gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n312_), .B(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n316_), .A2(new_n210_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n210_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G227gat), .A2(G233gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n319_), .B(G15gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT30), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT31), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OR3_X1    g122(.A1(new_n317_), .A2(new_n318_), .A3(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n323_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n257_), .A2(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G78gat), .B(G106gat), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G22gat), .B(G50gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n236_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n236_), .B2(new_n333_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n331_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT28), .B1(new_n234_), .B2(KEYINPUT29), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n236_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n330_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n339_), .A3(KEYINPUT92), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT91), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n236_), .A2(new_n333_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT89), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G211gat), .B(G218gat), .ZN(new_n345_));
  OR2_X1    g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT21), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n344_), .B(new_n345_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G218gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G211gat), .ZN(new_n352_));
  INV_X1    g151(.A(G211gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G218gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n354_), .A3(new_n344_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n355_), .A2(KEYINPUT21), .A3(new_n346_), .A4(new_n347_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n348_), .A2(new_n345_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n342_), .B1(new_n343_), .B2(new_n362_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n356_), .A2(new_n350_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n341_), .B(KEYINPUT91), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n364_), .B(new_n365_), .C1(new_n333_), .C2(new_n236_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n329_), .B1(new_n340_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT92), .B1(new_n336_), .B2(new_n339_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n340_), .A2(new_n367_), .A3(new_n329_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n370_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n340_), .A2(new_n329_), .A3(new_n367_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n373_), .B1(new_n374_), .B2(new_n368_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT18), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT19), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n287_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n276_), .A2(new_n280_), .A3(KEYINPUT82), .ZN(new_n386_));
  OAI22_X1  g185(.A1(new_n385_), .A2(new_n386_), .B1(new_n308_), .B2(new_n307_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n310_), .A2(new_n309_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(new_n302_), .B2(KEYINPUT84), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n271_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n384_), .B1(new_n390_), .B2(new_n364_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n267_), .B(new_n294_), .C1(new_n268_), .C2(new_n265_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(G183gat), .B(G190gat), .C1(new_n297_), .C2(new_n298_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n395_), .A2(KEYINPUT93), .A3(new_n267_), .A4(new_n294_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n289_), .A2(new_n290_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n397_), .A2(new_n273_), .B1(new_n310_), .B2(new_n309_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  OAI22_X1  g198(.A1(new_n306_), .A2(new_n300_), .B1(G183gat), .B2(G190gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n262_), .A2(KEYINPUT94), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n260_), .A2(KEYINPUT22), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT22), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(G169gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n402_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n401_), .A2(new_n406_), .A3(new_n258_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n400_), .A2(new_n407_), .A3(new_n264_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n399_), .A2(new_n362_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n383_), .B1(new_n391_), .B2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n362_), .B(new_n271_), .C1(new_n387_), .C2(new_n389_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n399_), .A2(new_n408_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n364_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(KEYINPUT20), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n414_), .A2(new_n382_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n380_), .B1(new_n410_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n382_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n380_), .ZN(new_n418_));
  OAI211_X1 g217(.A(KEYINPUT20), .B(new_n383_), .C1(new_n312_), .C2(new_n362_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT95), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n409_), .A2(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n399_), .A2(new_n362_), .A3(new_n408_), .A4(KEYINPUT95), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n417_), .B(new_n418_), .C1(new_n419_), .C2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n416_), .A2(KEYINPUT27), .A3(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n419_), .A2(new_n423_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n384_), .B1(new_n412_), .B2(new_n364_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n383_), .B1(new_n427_), .B2(new_n411_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n380_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n424_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT27), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT99), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT99), .ZN(new_n433_));
  AOI211_X1 g232(.A(new_n433_), .B(KEYINPUT27), .C1(new_n429_), .C2(new_n424_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n376_), .B(new_n425_), .C1(new_n432_), .C2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT100), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n426_), .A2(new_n428_), .A3(new_n380_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n391_), .A2(new_n383_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n418_), .B1(new_n438_), .B2(new_n417_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n431_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n433_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n430_), .A2(KEYINPUT99), .A3(new_n431_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT100), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n376_), .A4(new_n425_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n327_), .B1(new_n436_), .B2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n324_), .A2(KEYINPUT87), .A3(new_n325_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT87), .B1(new_n324_), .B2(new_n325_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n254_), .A2(new_n256_), .B1(new_n375_), .B2(new_n372_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n443_), .A2(new_n450_), .A3(new_n425_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n418_), .A2(KEYINPUT32), .ZN(new_n452_));
  OR3_X1    g251(.A1(new_n426_), .A2(new_n428_), .A3(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n452_), .B1(new_n410_), .B2(new_n415_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n253_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n238_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n235_), .A2(new_n240_), .A3(new_n237_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n458_), .A2(new_n249_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n252_), .A2(new_n456_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n243_), .A2(KEYINPUT33), .A3(new_n251_), .A4(new_n244_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT97), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n455_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n376_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n449_), .B1(new_n451_), .B2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n446_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT6), .ZN(new_n469_));
  INV_X1    g268(.A(G85gat), .ZN(new_n470_));
  INV_X1    g269(.A(G92gat), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT9), .ZN(new_n472_));
  XOR2_X1   g271(.A(G85gat), .B(G92gat), .Z(new_n473_));
  AOI21_X1  g272(.A(new_n472_), .B1(new_n473_), .B2(KEYINPUT9), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT10), .B(G99gat), .Z(new_n475_));
  INV_X1    g274(.A(G106gat), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n475_), .A2(KEYINPUT65), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT65), .B1(new_n475_), .B2(new_n476_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n469_), .B(new_n474_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(G99gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(new_n476_), .A3(KEYINPUT67), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT67), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(G99gat), .B2(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT7), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT68), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT66), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n481_), .A2(new_n483_), .A3(new_n490_), .A4(new_n484_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n486_), .A2(new_n489_), .A3(new_n469_), .A4(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n473_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n492_), .B2(new_n473_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n479_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT71), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G29gat), .B(G36gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT74), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n499_), .A2(KEYINPUT74), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n501_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G29gat), .B(G36gat), .Z(new_n506_));
  INV_X1    g305(.A(KEYINPUT74), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n503_), .B1(new_n508_), .B2(new_n500_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n498_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(KEYINPUT15), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n515_), .B(new_n479_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n497_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT35), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n520_), .A2(new_n521_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT76), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n496_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n511_), .A2(new_n512_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n525_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n517_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n523_), .A2(new_n524_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n517_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G190gat), .B(G218gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G134gat), .B(G162gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n537_), .A2(KEYINPUT36), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT75), .B1(new_n533_), .B2(new_n534_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n537_), .A2(KEYINPUT36), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n539_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT75), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n517_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n531_), .B1(new_n517_), .B2(new_n529_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n544_), .B(new_n542_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT37), .B1(new_n543_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n545_), .A2(new_n546_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n550_), .A2(new_n541_), .B1(new_n551_), .B2(new_n538_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n547_), .ZN(new_n554_));
  INV_X1    g353(.A(G1gat), .ZN(new_n555_));
  INV_X1    g354(.A(G8gat), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT77), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT77), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n559_), .B(KEYINPUT14), .C1(new_n555_), .C2(new_n556_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(G1gat), .B(G8gat), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n558_), .A2(new_n563_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT11), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT69), .B(G71gat), .Z(new_n573_));
  INV_X1    g372(.A(G78gat), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n571_), .A2(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(KEYINPUT69), .A2(G71gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(KEYINPUT69), .A2(G71gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(G78gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n570_), .A2(KEYINPUT11), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT70), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT70), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n570_), .A2(new_n582_), .A3(KEYINPUT11), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n575_), .A2(new_n579_), .A3(new_n581_), .A4(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n583_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n576_), .A2(new_n574_), .A3(new_n577_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n579_), .B(new_n586_), .C1(KEYINPUT11), .C2(new_n570_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n569_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G127gat), .B(G155gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT16), .ZN(new_n593_));
  XOR2_X1   g392(.A(G183gat), .B(G211gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n590_), .A2(new_n591_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(KEYINPUT17), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n590_), .B2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n549_), .A2(new_n554_), .A3(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n467_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n589_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n497_), .A2(KEYINPUT12), .A3(new_n601_), .A4(new_n516_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT64), .Z(new_n604_));
  OAI211_X1 g403(.A(new_n589_), .B(new_n479_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT12), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n496_), .A2(new_n601_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(new_n604_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT72), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n607_), .A2(new_n605_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(new_n604_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT72), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n602_), .A2(new_n608_), .A3(new_n613_), .A4(new_n604_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT5), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n610_), .A2(new_n612_), .A3(new_n614_), .A4(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(KEYINPUT13), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT80), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n505_), .A2(new_n509_), .A3(new_n498_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT15), .B1(new_n511_), .B2(new_n512_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n567_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT78), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G229gat), .A2(G233gat), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n511_), .A2(new_n565_), .A3(new_n566_), .A4(new_n512_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .A4(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT79), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G169gat), .B(G197gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n510_), .A2(new_n513_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n630_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n631_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  AOI22_X1  g439(.A1(new_n511_), .A2(new_n512_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n638_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT78), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n632_), .B(new_n636_), .C1(new_n640_), .C2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n628_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n527_), .A2(new_n567_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n631_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n629_), .B1(new_n648_), .B2(new_n638_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n636_), .B1(new_n650_), .B2(new_n632_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n625_), .B1(new_n645_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n632_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n636_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(KEYINPUT80), .A3(new_n644_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT13), .B1(new_n620_), .B2(new_n622_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n624_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n600_), .A2(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n661_), .A2(G1gat), .A3(new_n257_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT38), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(KEYINPUT38), .ZN(new_n664_));
  INV_X1    g463(.A(new_n327_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n425_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n444_), .B1(new_n667_), .B2(new_n376_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n435_), .A2(KEYINPUT100), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n451_), .A2(new_n465_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n449_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n543_), .A2(new_n548_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n659_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n623_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n598_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n677_), .A2(new_n658_), .A3(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n674_), .A2(new_n675_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G1gat), .B1(new_n680_), .B2(new_n257_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n663_), .A2(new_n664_), .A3(new_n681_), .ZN(G1324gat));
  OAI21_X1  g481(.A(G8gat), .B1(new_n680_), .B2(new_n667_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT101), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(KEYINPUT101), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(KEYINPUT39), .A3(new_n685_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n685_), .A2(KEYINPUT39), .ZN(new_n687_));
  INV_X1    g486(.A(new_n667_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n600_), .A2(new_n556_), .A3(new_n660_), .A4(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n686_), .A2(new_n687_), .A3(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n686_), .A2(new_n687_), .A3(new_n689_), .A4(new_n691_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1325gat));
  OAI21_X1  g494(.A(G15gat), .B1(new_n680_), .B2(new_n672_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n697_), .ZN(new_n699_));
  OR3_X1    g498(.A1(new_n661_), .A2(G15gat), .A3(new_n672_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(G1326gat));
  OAI21_X1  g500(.A(G22gat), .B1(new_n680_), .B2(new_n376_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT42), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n376_), .A2(G22gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n661_), .B2(new_n704_), .ZN(G1327gat));
  NOR2_X1   g504(.A1(new_n675_), .A2(new_n598_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n674_), .A2(KEYINPUT105), .A3(new_n660_), .A4(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n660_), .B(new_n706_), .C1(new_n446_), .C2(new_n466_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n257_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G29gat), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n549_), .A2(new_n554_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n549_), .A2(new_n554_), .A3(KEYINPUT104), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n718_), .B(new_n719_), .C1(new_n446_), .C2(new_n466_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n716_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n720_), .A2(KEYINPUT43), .B1(new_n674_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n660_), .A2(new_n678_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n715_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n725_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n719_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT104), .B1(new_n549_), .B2(new_n554_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n721_), .B1(new_n674_), .B2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n467_), .A2(new_n722_), .ZN(new_n732_));
  OAI211_X1 g531(.A(KEYINPUT44), .B(new_n727_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n726_), .A2(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n713_), .A2(G29gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n714_), .B1(new_n734_), .B2(new_n735_), .ZN(G1328gat));
  NAND3_X1  g535(.A1(new_n726_), .A2(new_n688_), .A3(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G36gat), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n667_), .A2(G36gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n707_), .A2(new_n710_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT106), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n707_), .A2(new_n710_), .A3(new_n743_), .A4(new_n739_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n741_), .A2(new_n742_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n742_), .B1(new_n741_), .B2(new_n744_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n738_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT107), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT108), .Z(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n747_), .A2(new_n751_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n738_), .B(new_n750_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1329gat));
  AOI21_X1  g553(.A(new_n314_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n726_), .A2(new_n733_), .A3(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n726_), .A2(new_n733_), .A3(KEYINPUT109), .A4(new_n755_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n314_), .B1(new_n711_), .B2(new_n672_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .A4(new_n762_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1330gat));
  INV_X1    g565(.A(new_n376_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G50gat), .B1(new_n712_), .B2(new_n767_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n767_), .A2(G50gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n734_), .B2(new_n769_), .ZN(G1331gat));
  INV_X1    g569(.A(new_n677_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n657_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n674_), .A2(new_n772_), .A3(new_n598_), .A4(new_n675_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G57gat), .B1(new_n773_), .B2(new_n257_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n600_), .A2(new_n772_), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n257_), .A2(G57gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n774_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT111), .ZN(G1332gat));
  OAI21_X1  g577(.A(G64gat), .B1(new_n773_), .B2(new_n667_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT48), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n667_), .A2(G64gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n775_), .B2(new_n781_), .ZN(G1333gat));
  OAI21_X1  g581(.A(G71gat), .B1(new_n773_), .B2(new_n672_), .ZN(new_n783_));
  XOR2_X1   g582(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n672_), .A2(G71gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n775_), .B2(new_n786_), .ZN(G1334gat));
  OAI21_X1  g586(.A(G78gat), .B1(new_n773_), .B2(new_n376_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT50), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n767_), .A2(new_n574_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n789_), .B1(new_n775_), .B2(new_n790_), .ZN(G1335gat));
  NOR3_X1   g590(.A1(new_n467_), .A2(new_n598_), .A3(new_n675_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n772_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n470_), .A3(new_n713_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n772_), .A2(new_n678_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n720_), .A2(KEYINPUT43), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n674_), .A2(new_n723_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n724_), .A2(KEYINPUT113), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n802_), .A2(new_n257_), .A3(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n795_), .B1(new_n804_), .B2(new_n470_), .ZN(G1336gat));
  NAND3_X1  g604(.A1(new_n794_), .A2(new_n471_), .A3(new_n688_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n802_), .A2(new_n667_), .A3(new_n803_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n471_), .ZN(G1337gat));
  NAND2_X1  g607(.A1(new_n326_), .A2(new_n475_), .ZN(new_n809_));
  OR3_X1    g608(.A1(new_n793_), .A2(KEYINPUT114), .A3(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT114), .B1(new_n793_), .B2(new_n809_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n802_), .A2(new_n672_), .A3(new_n803_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n480_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  OAI221_X1 g617(.A(new_n812_), .B1(new_n815_), .B2(new_n816_), .C1(new_n813_), .C2(new_n480_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1338gat));
  NAND3_X1  g619(.A1(new_n794_), .A2(new_n476_), .A3(new_n767_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n796_), .A2(new_n376_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n800_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n824_), .B2(G106gat), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT52), .B(new_n476_), .C1(new_n800_), .C2(new_n823_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n821_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g627(.A1(new_n624_), .A2(new_n657_), .A3(new_n659_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n549_), .A2(new_n554_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .A4(new_n598_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n676_), .A2(new_n658_), .A3(new_n623_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT54), .B1(new_n833_), .B2(new_n599_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n628_), .A2(new_n638_), .A3(new_n631_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n654_), .B1(new_n648_), .B2(new_n630_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n651_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n657_), .A2(new_n622_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n610_), .A2(new_n844_), .A3(new_n614_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n604_), .B1(new_n602_), .B2(new_n608_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n602_), .A2(new_n604_), .A3(new_n608_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(KEYINPUT55), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n619_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n843_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n621_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n851_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n842_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n675_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n837_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n855_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n657_), .B(new_n622_), .C1(new_n854_), .C2(new_n851_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT57), .B(new_n675_), .C1(new_n861_), .C2(new_n842_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n854_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n622_), .A2(new_n840_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n854_), .B2(new_n865_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n863_), .B(new_n864_), .C1(new_n867_), .C2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n716_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n850_), .A2(KEYINPUT56), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n866_), .A3(new_n868_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n864_), .B1(new_n873_), .B2(new_n863_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n858_), .B(new_n862_), .C1(new_n871_), .C2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n836_), .B1(new_n875_), .B2(new_n678_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n713_), .B(new_n326_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT118), .Z(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n876_), .A2(new_n879_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n876_), .A2(new_n879_), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n657_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G113gat), .ZN(new_n886_));
  INV_X1    g685(.A(new_n880_), .ZN(new_n887_));
  OR3_X1    g686(.A1(new_n887_), .A2(G113gat), .A3(new_n658_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1340gat));
  INV_X1    g688(.A(G120gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n771_), .B2(KEYINPUT60), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n880_), .B(new_n891_), .C1(KEYINPUT60), .C2(new_n890_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n883_), .A2(new_n677_), .A3(new_n884_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n890_), .ZN(G1341gat));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895_));
  INV_X1    g694(.A(G127gat), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n895_), .B(new_n896_), .C1(new_n887_), .C2(new_n678_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n883_), .A2(G127gat), .A3(new_n598_), .A4(new_n884_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n876_), .A2(new_n879_), .A3(new_n678_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT120), .B1(new_n899_), .B2(G127gat), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n897_), .A2(new_n898_), .A3(new_n900_), .ZN(G1342gat));
  AOI21_X1  g700(.A(G134gat), .B1(new_n880_), .B2(new_n857_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n883_), .A2(new_n884_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n716_), .A2(G134gat), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT121), .Z(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n903_), .B2(new_n905_), .ZN(G1343gat));
  NAND3_X1  g705(.A1(new_n672_), .A2(new_n767_), .A3(new_n713_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n688_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n876_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n657_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n677_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n598_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT61), .B(G155gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1346gat));
  NOR3_X1   g716(.A1(new_n876_), .A2(new_n675_), .A3(new_n909_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(G162gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n875_), .A2(new_n678_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n835_), .ZN(new_n921_));
  AND4_X1   g720(.A1(G162gat), .A2(new_n921_), .A3(new_n730_), .A4(new_n908_), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT122), .B1(new_n919_), .B2(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n910_), .A2(G162gat), .A3(new_n730_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n924_), .B(new_n925_), .C1(G162gat), .C2(new_n918_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n923_), .A2(new_n926_), .ZN(G1347gat));
  NOR3_X1   g726(.A1(new_n672_), .A2(new_n713_), .A3(new_n667_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n657_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT123), .Z(new_n930_));
  NAND3_X1  g729(.A1(new_n921_), .A2(new_n930_), .A3(new_n376_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n931_), .A2(new_n932_), .A3(G169gat), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n931_), .B2(G169gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n921_), .A2(new_n376_), .A3(new_n928_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n657_), .A2(new_n406_), .A3(new_n401_), .ZN(new_n936_));
  OAI22_X1  g735(.A1(new_n933_), .A2(new_n934_), .B1(new_n935_), .B2(new_n936_), .ZN(G1348gat));
  NOR2_X1   g736(.A1(new_n935_), .A2(new_n771_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n258_), .ZN(G1349gat));
  NOR3_X1   g738(.A1(new_n935_), .A2(new_n273_), .A3(new_n678_), .ZN(new_n940_));
  OR2_X1    g739(.A1(new_n935_), .A2(new_n678_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n282_), .B2(new_n941_), .ZN(G1350gat));
  NOR3_X1   g741(.A1(new_n675_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n921_), .A2(new_n376_), .A3(new_n928_), .A4(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n928_), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n876_), .A2(new_n767_), .A3(new_n830_), .A4(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n944_), .B1(new_n946_), .B2(new_n274_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(KEYINPUT124), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n949_), .B(new_n944_), .C1(new_n946_), .C2(new_n274_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n950_), .ZN(G1351gat));
  NOR4_X1   g750(.A1(new_n449_), .A2(new_n667_), .A3(new_n376_), .A4(new_n713_), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n921_), .A2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(new_n657_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g754(.A1(new_n921_), .A2(new_n952_), .ZN(new_n956_));
  OAI22_X1  g755(.A1(new_n956_), .A2(new_n771_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n957_));
  NAND2_X1  g756(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n958_));
  XOR2_X1   g757(.A(new_n958_), .B(KEYINPUT126), .Z(new_n959_));
  INV_X1    g758(.A(new_n959_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n957_), .B(new_n960_), .ZN(G1353gat));
  AND3_X1   g760(.A1(new_n921_), .A2(new_n598_), .A3(new_n952_), .ZN(new_n962_));
  XOR2_X1   g761(.A(KEYINPUT63), .B(G211gat), .Z(new_n963_));
  AOI21_X1  g762(.A(KEYINPUT127), .B1(new_n962_), .B2(new_n963_), .ZN(new_n964_));
  NAND4_X1  g763(.A1(new_n921_), .A2(new_n598_), .A3(new_n952_), .A4(new_n963_), .ZN(new_n965_));
  OR2_X1    g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n962_), .B2(new_n966_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n964_), .B1(KEYINPUT127), .B2(new_n967_), .ZN(G1354gat));
  NAND3_X1  g767(.A1(new_n953_), .A2(new_n351_), .A3(new_n857_), .ZN(new_n969_));
  OAI21_X1  g768(.A(G218gat), .B1(new_n956_), .B2(new_n830_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1355gat));
endmodule


