//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G85gat), .ZN(new_n204_));
  INV_X1    g003(.A(G92gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT6), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n212_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n208_), .B1(new_n215_), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT8), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT10), .B(G99gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n210_), .B1(G106gat), .B2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n206_), .B1(KEYINPUT9), .B2(new_n207_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT67), .ZN(new_n231_));
  XOR2_X1   g030(.A(G71gat), .B(G78gat), .Z(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(KEYINPUT11), .B2(new_n229_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n233_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n228_), .A2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n227_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n203_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n239_), .A2(KEYINPUT68), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(KEYINPUT68), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT12), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n236_), .B2(KEYINPUT70), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n226_), .B(KEYINPUT69), .ZN(new_n244_));
  INV_X1    g043(.A(new_n220_), .ZN(new_n245_));
  OAI221_X1 g044(.A(new_n243_), .B1(KEYINPUT70), .B2(new_n236_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n238_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n242_), .B1(new_n228_), .B2(new_n236_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n246_), .A2(new_n202_), .A3(new_n247_), .A4(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n240_), .A2(new_n241_), .A3(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G120gat), .B(G148gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT5), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G176gat), .B(G204gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT72), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n254_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT71), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT13), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n256_), .A2(KEYINPUT13), .A3(new_n258_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT73), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT80), .ZN(new_n265_));
  XOR2_X1   g064(.A(G190gat), .B(G218gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT75), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G134gat), .B(G162gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT36), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n244_), .A2(new_n245_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G29gat), .B(G36gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT74), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G43gat), .B(G50gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT15), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n272_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G232gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT34), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n281_), .A2(KEYINPUT35), .ZN(new_n282_));
  INV_X1    g081(.A(new_n276_), .ZN(new_n283_));
  OAI22_X1  g082(.A1(new_n227_), .A2(new_n283_), .B1(KEYINPUT35), .B2(new_n281_), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n279_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n282_), .B1(new_n279_), .B2(new_n284_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n271_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n269_), .A2(new_n270_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n288_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT37), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT76), .B1(new_n287_), .B2(new_n288_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT37), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT77), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n291_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n291_), .B1(new_n298_), .B2(new_n295_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G231gat), .A2(G233gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n302_), .B(KEYINPUT79), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n236_), .B(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G1gat), .B(G8gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT78), .ZN(new_n306_));
  INV_X1    g105(.A(G15gat), .ZN(new_n307_));
  INV_X1    g106(.A(G22gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G15gat), .A2(G22gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G1gat), .A2(G8gat), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n309_), .A2(new_n310_), .B1(KEYINPUT14), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n306_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n304_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G127gat), .B(G155gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT16), .ZN(new_n317_));
  XOR2_X1   g116(.A(G183gat), .B(G211gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(KEYINPUT70), .A3(KEYINPUT17), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n321_), .B1(KEYINPUT17), .B2(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n314_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n265_), .B1(new_n301_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n295_), .A2(new_n298_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n291_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n291_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(KEYINPUT80), .A3(new_n325_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n264_), .A2(new_n327_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT101), .ZN(new_n335_));
  INV_X1    g134(.A(G169gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT22), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT22), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(G169gat), .ZN(new_n339_));
  INV_X1    g138(.A(G176gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT99), .ZN(new_n344_));
  INV_X1    g143(.A(G183gat), .ZN(new_n345_));
  INV_X1    g144(.A(G190gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT86), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(KEYINPUT86), .A2(G183gat), .A3(G190gat), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT23), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(KEYINPUT23), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n347_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT99), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n341_), .A2(new_n356_), .A3(new_n342_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n344_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n345_), .A2(KEYINPUT25), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n346_), .A2(KEYINPUT26), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT26), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(G190gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G183gat), .ZN(new_n364_));
  AND4_X1   g163(.A1(new_n359_), .A2(new_n360_), .A3(new_n362_), .A4(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT24), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n342_), .A2(KEYINPUT24), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n366_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(KEYINPUT86), .A2(G183gat), .A3(G190gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT86), .B1(G183gat), .B2(G190gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT23), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n348_), .A2(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n358_), .A2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G211gat), .B(G218gat), .Z(new_n380_));
  OR2_X1    g179(.A1(KEYINPUT97), .A2(G197gat), .ZN(new_n381_));
  INV_X1    g180(.A(G204gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(KEYINPUT97), .A2(G197gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT21), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(G197gat), .B2(G204gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n380_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n382_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(G197gat), .A2(G204gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n385_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n388_), .A2(new_n389_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G211gat), .B(G218gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(new_n385_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n335_), .B1(new_n379_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n374_), .A2(new_n347_), .A3(new_n376_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT88), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT88), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n374_), .A2(new_n400_), .A3(new_n347_), .A4(new_n376_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n340_), .B1(new_n338_), .B2(KEYINPUT87), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G169gat), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n336_), .B(new_n340_), .C1(new_n338_), .C2(KEYINPUT87), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(new_n401_), .A3(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n408_));
  NOR2_X1   g207(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n409_));
  OAI21_X1  g208(.A(G183gat), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT85), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n360_), .A2(new_n362_), .ZN(new_n413_));
  OAI211_X1 g212(.A(KEYINPUT85), .B(G183gat), .C1(new_n408_), .C2(new_n409_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n412_), .A2(new_n359_), .A3(new_n413_), .A4(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n375_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n370_), .B1(new_n353_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n407_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n396_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n387_), .A2(new_n390_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n421_), .A2(new_n358_), .A3(KEYINPUT101), .A4(new_n378_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT19), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n397_), .A2(new_n420_), .A3(new_n422_), .A4(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n407_), .A2(new_n421_), .A3(new_n418_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT20), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n379_), .A2(new_n396_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT100), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n379_), .A2(KEYINPUT100), .A3(new_n396_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n429_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n424_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n427_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT18), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n438_), .B(new_n439_), .Z(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT27), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n379_), .A2(new_n396_), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT107), .B(KEYINPUT20), .Z(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n435_), .B1(new_n447_), .B2(new_n420_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n405_), .B1(new_n398_), .B2(KEYINPUT88), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n449_), .A2(new_n401_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n425_), .B1(new_n450_), .B2(new_n421_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n379_), .A2(KEYINPUT100), .A3(new_n396_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT100), .B1(new_n379_), .B2(new_n396_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n435_), .B(new_n451_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n448_), .B1(new_n454_), .B2(KEYINPUT108), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n454_), .A2(KEYINPUT108), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n440_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n444_), .B1(new_n457_), .B2(KEYINPUT111), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT111), .ZN(new_n459_));
  AOI211_X1 g258(.A(new_n459_), .B(new_n440_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT112), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n455_), .A2(new_n456_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n441_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n459_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT112), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n457_), .A2(KEYINPUT111), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .A4(new_n444_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n461_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT102), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n436_), .B2(new_n441_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n424_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n472_), .A2(KEYINPUT102), .A3(new_n440_), .A4(new_n427_), .ZN(new_n473_));
  AOI211_X1 g272(.A(KEYINPUT103), .B(new_n440_), .C1(new_n472_), .C2(new_n427_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT103), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n436_), .B2(new_n441_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n470_), .B(new_n473_), .C1(new_n474_), .C2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n443_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n468_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G155gat), .A2(G162gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(KEYINPUT1), .ZN(new_n481_));
  NOR2_X1   g280(.A1(G155gat), .A2(G162gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n482_), .B2(KEYINPUT1), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n481_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(new_n484_), .B2(new_n483_), .ZN(new_n486_));
  AND3_X1   g285(.A1(KEYINPUT90), .A2(G141gat), .A3(G148gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT90), .B1(G141gat), .B2(G148gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G141gat), .ZN(new_n490_));
  INV_X1    g289(.A(G148gat), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT92), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n500_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT2), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n497_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n480_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(new_n482_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n505_), .A2(KEYINPUT93), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT93), .B1(new_n505_), .B2(new_n507_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n493_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT94), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n493_), .B(new_n512_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT29), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G22gat), .B(G50gat), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n517_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n514_), .A2(new_n515_), .A3(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n524_));
  AOI211_X1 g323(.A(KEYINPUT29), .B(new_n517_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n519_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G78gat), .B(G106gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT98), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n528_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n523_), .A2(new_n526_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n511_), .A2(KEYINPUT29), .A3(new_n513_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT96), .Z(new_n536_));
  AND2_X1   g335(.A1(G228gat), .A2(G233gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n421_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n510_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n396_), .B1(new_n540_), .B2(new_n515_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n537_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n534_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n479_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G127gat), .B(G134gat), .Z(new_n549_));
  XOR2_X1   g348(.A(G113gat), .B(G120gat), .Z(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  NAND3_X1  g350(.A1(new_n511_), .A2(new_n513_), .A3(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n510_), .A2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G225gat), .A2(G233gat), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n552_), .A2(KEYINPUT4), .A3(new_n553_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT4), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n511_), .A2(new_n557_), .A3(new_n513_), .A4(new_n551_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n554_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n555_), .B1(new_n556_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G1gat), .B(G29gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(G85gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT0), .B(G57gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n555_), .B(new_n565_), .C1(new_n556_), .C2(new_n560_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(KEYINPUT109), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT109), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n561_), .A2(new_n570_), .A3(new_n566_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G71gat), .B(G99gat), .ZN(new_n574_));
  INV_X1    g373(.A(G43gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n450_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n551_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G227gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(new_n307_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT30), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT31), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n578_), .B(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n573_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n548_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT104), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n568_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n552_), .A2(KEYINPUT4), .A3(new_n553_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n559_), .A3(new_n558_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n591_), .A2(KEYINPUT104), .A3(new_n555_), .A4(new_n565_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(new_n589_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT105), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n554_), .A3(new_n558_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n552_), .A2(new_n553_), .A3(new_n559_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n566_), .A3(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n597_), .B1(new_n568_), .B2(new_n589_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n477_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT105), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n588_), .A2(new_n600_), .A3(new_n589_), .A4(new_n592_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n594_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n440_), .A2(KEYINPUT32), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT106), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n603_), .B1(new_n436_), .B2(new_n604_), .ZN(new_n605_));
  OAI211_X1 g404(.A(KEYINPUT32), .B(new_n440_), .C1(new_n436_), .C2(KEYINPUT106), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(new_n606_), .B2(new_n462_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n569_), .A2(new_n607_), .A3(new_n571_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT110), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n569_), .A2(new_n607_), .A3(KEYINPUT110), .A4(new_n571_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n602_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n547_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n461_), .A2(new_n467_), .B1(new_n443_), .B2(new_n477_), .ZN(new_n615_));
  AOI22_X1  g414(.A1(new_n545_), .A2(new_n546_), .B1(new_n571_), .B2(new_n569_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n583_), .B(KEYINPUT89), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(KEYINPUT113), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT113), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n612_), .A2(new_n613_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n619_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n621_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n586_), .B1(new_n620_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n313_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n277_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n313_), .A2(new_n276_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G229gat), .A2(G233gat), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT81), .Z(new_n630_));
  NAND3_X1  g429(.A1(new_n627_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n313_), .B(new_n276_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(G229gat), .A3(G233gat), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT82), .ZN(new_n636_));
  XOR2_X1   g435(.A(G169gat), .B(G197gat), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n634_), .A2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT83), .Z(new_n640_));
  OR2_X1    g439(.A1(new_n634_), .A2(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n625_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n334_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n572_), .A2(G1gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT113), .B1(new_n618_), .B2(new_n619_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n622_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n585_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n329_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n263_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(new_n325_), .A3(new_n642_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n573_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G1gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n648_), .A2(new_n657_), .ZN(new_n658_));
  MUX2_X1   g457(.A(new_n648_), .B(new_n658_), .S(KEYINPUT38), .Z(G1324gat));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n655_), .A2(new_n479_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(G8gat), .ZN(new_n662_));
  INV_X1    g461(.A(G8gat), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT39), .B(new_n663_), .C1(new_n655_), .C2(new_n479_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n479_), .A2(new_n663_), .ZN(new_n665_));
  OAI22_X1  g464(.A1(new_n662_), .A2(new_n664_), .B1(new_n645_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT114), .B(KEYINPUT40), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n666_), .B(new_n668_), .ZN(G1325gat));
  NAND2_X1  g468(.A1(new_n655_), .A2(new_n623_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G15gat), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT115), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT115), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n673_), .A3(G15gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(KEYINPUT41), .A3(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n646_), .A2(new_n307_), .A3(new_n623_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT41), .B1(new_n672_), .B2(new_n674_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1326gat));
  NAND3_X1  g478(.A1(new_n646_), .A2(new_n308_), .A3(new_n547_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n655_), .A2(new_n547_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT116), .B(KEYINPUT42), .Z(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(G22gat), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G22gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1327gat));
  NAND2_X1  g484(.A1(new_n291_), .A2(new_n326_), .ZN(new_n686_));
  NOR4_X1   g485(.A1(new_n625_), .A2(new_n643_), .A3(new_n263_), .A4(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G29gat), .B1(new_n687_), .B2(new_n573_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n651_), .A2(new_n689_), .A3(new_n301_), .ZN(new_n690_));
  XOR2_X1   g489(.A(KEYINPUT117), .B(KEYINPUT43), .Z(new_n691_));
  OAI21_X1  g490(.A(new_n691_), .B1(new_n625_), .B2(new_n332_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n263_), .A2(new_n325_), .A3(new_n643_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT44), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  INV_X1    g495(.A(new_n694_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n696_), .B(new_n697_), .C1(new_n690_), .C2(new_n692_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n695_), .A2(new_n698_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n573_), .A2(G29gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n688_), .B1(new_n699_), .B2(new_n700_), .ZN(G1328gat));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  INV_X1    g501(.A(G36gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n699_), .B2(new_n479_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n615_), .B(KEYINPUT118), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n687_), .A2(new_n703_), .A3(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT45), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n702_), .B1(new_n704_), .B2(new_n709_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n695_), .A2(new_n698_), .A3(new_n615_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT46), .B(new_n708_), .C1(new_n711_), .C2(new_n703_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1329gat));
  INV_X1    g512(.A(new_n695_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n694_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n583_), .A2(new_n575_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n714_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G43gat), .B1(new_n687_), .B2(new_n623_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT47), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n699_), .B2(new_n716_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1330gat));
  INV_X1    g522(.A(G50gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n687_), .A2(new_n724_), .A3(new_n547_), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT119), .B(new_n724_), .C1(new_n699_), .C2(new_n547_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT119), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n714_), .A2(new_n547_), .A3(new_n715_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(G50gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n726_), .B2(new_n729_), .ZN(G1331gat));
  NAND3_X1  g529(.A1(new_n327_), .A2(new_n333_), .A3(new_n263_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT120), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n625_), .A2(new_n642_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(KEYINPUT120), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n572_), .B1(new_n735_), .B2(KEYINPUT121), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(KEYINPUT121), .B2(new_n735_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n642_), .A2(new_n326_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n652_), .A2(new_n264_), .A3(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n572_), .A2(new_n738_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n737_), .A2(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(G1332gat));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n741_), .B2(new_n706_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT48), .Z(new_n746_));
  NAND2_X1  g545(.A1(new_n706_), .A2(new_n744_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n735_), .B2(new_n747_), .ZN(G1333gat));
  INV_X1    g547(.A(G71gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n741_), .B2(new_n623_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT49), .Z(new_n751_));
  NAND2_X1  g550(.A1(new_n623_), .A2(new_n749_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT122), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n735_), .B2(new_n753_), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n741_), .A2(new_n547_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(G78gat), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n613_), .A2(G78gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n735_), .B2(new_n758_), .ZN(G1335gat));
  NOR3_X1   g558(.A1(new_n653_), .A2(new_n325_), .A3(new_n642_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n693_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n572_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n264_), .A2(new_n686_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n733_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n573_), .A2(new_n204_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(new_n764_), .B2(new_n765_), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n761_), .B2(new_n705_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n479_), .A2(new_n205_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n764_), .B2(new_n768_), .ZN(G1337gat));
  OR2_X1    g568(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n770_));
  NAND2_X1  g569(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n771_));
  OAI21_X1  g570(.A(G99gat), .B1(new_n761_), .B2(new_n619_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n764_), .A2(new_n583_), .A3(new_n221_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n770_), .B(new_n771_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n774_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n776_), .A2(KEYINPUT123), .A3(KEYINPUT51), .A4(new_n772_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1338gat));
  OR3_X1    g577(.A1(new_n764_), .A2(G106gat), .A3(new_n613_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n693_), .A2(new_n547_), .A3(new_n760_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT124), .B(KEYINPUT52), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(G106gat), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(G106gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT53), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n779_), .B(new_n786_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1339gat));
  NAND3_X1  g587(.A1(new_n261_), .A2(new_n262_), .A3(new_n739_), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n789_), .A2(new_n301_), .A3(KEYINPUT54), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT54), .B1(new_n789_), .B2(new_n301_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n630_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n627_), .A2(new_n628_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n638_), .B1(new_n632_), .B2(new_n630_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n640_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n259_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n203_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT55), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(new_n249_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n249_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n254_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT56), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n254_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n256_), .A2(new_n806_), .A3(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n799_), .B1(new_n643_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n329_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(KEYINPUT57), .A3(new_n329_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT125), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n256_), .A2(new_n806_), .A3(new_n798_), .A4(new_n808_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n301_), .A2(new_n815_), .A3(new_n818_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n816_), .A2(new_n817_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n815_), .B1(new_n301_), .B2(new_n818_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n813_), .B(new_n814_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n793_), .B1(new_n823_), .B2(new_n326_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n548_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n825_), .A2(new_n572_), .A3(new_n583_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n824_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(G113gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n642_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT126), .B(new_n831_), .C1(new_n824_), .C2(new_n827_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n823_), .A2(new_n326_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n792_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n831_), .A2(KEYINPUT126), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(KEYINPUT126), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n826_), .A4(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n643_), .B1(new_n832_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n838_), .B2(new_n829_), .ZN(G1340gat));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n653_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n828_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n264_), .B1(new_n832_), .B2(new_n837_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n840_), .ZN(G1341gat));
  INV_X1    g643(.A(G127gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n828_), .A2(new_n845_), .A3(new_n325_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n326_), .B1(new_n832_), .B2(new_n837_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n845_), .ZN(G1342gat));
  INV_X1    g647(.A(G134gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n828_), .A2(new_n849_), .A3(new_n291_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n332_), .B1(new_n832_), .B2(new_n837_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(G1343gat));
  NOR4_X1   g651(.A1(new_n706_), .A2(new_n572_), .A3(new_n613_), .A4(new_n623_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n834_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n643_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n490_), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n264_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n491_), .ZN(G1345gat));
  NOR2_X1   g657(.A1(new_n854_), .A2(new_n326_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT61), .B(G155gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1346gat));
  OAI21_X1  g660(.A(G162gat), .B1(new_n854_), .B2(new_n332_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n329_), .A2(G162gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n854_), .B2(new_n863_), .ZN(G1347gat));
  NOR3_X1   g663(.A1(new_n547_), .A2(new_n619_), .A3(new_n573_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n814_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n810_), .B2(new_n329_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n822_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n820_), .A3(new_n819_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n325_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n706_), .B(new_n865_), .C1(new_n871_), .C2(new_n793_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G169gat), .B1(new_n872_), .B2(new_n643_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n872_), .A2(new_n643_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT62), .B(G169gat), .C1(new_n872_), .C2(new_n643_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n875_), .A2(new_n877_), .A3(new_n878_), .ZN(G1348gat));
  OAI21_X1  g678(.A(G176gat), .B1(new_n872_), .B2(new_n264_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n263_), .A2(new_n340_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n872_), .B2(new_n881_), .ZN(G1349gat));
  NOR2_X1   g681(.A1(new_n872_), .A2(new_n326_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n359_), .A3(new_n364_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n345_), .B2(new_n883_), .ZN(G1350gat));
  OAI21_X1  g684(.A(G190gat), .B1(new_n872_), .B2(new_n332_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n291_), .A2(new_n413_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n872_), .B2(new_n887_), .ZN(G1351gat));
  INV_X1    g687(.A(G197gat), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n616_), .A2(new_n619_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n834_), .A2(new_n706_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n891_), .B2(new_n643_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n824_), .A2(new_n705_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n893_), .A2(G197gat), .A3(new_n642_), .A4(new_n890_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1352gat));
  OR3_X1    g694(.A1(new_n891_), .A2(G204gat), .A3(new_n264_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G204gat), .B1(new_n891_), .B2(new_n264_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1353gat));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n899_));
  INV_X1    g698(.A(G211gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n325_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  XOR2_X1   g700(.A(new_n901_), .B(KEYINPUT127), .Z(new_n902_));
  OAI211_X1 g701(.A(new_n899_), .B(new_n900_), .C1(new_n891_), .C2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n900_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n902_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n893_), .A2(new_n890_), .A3(new_n904_), .A4(new_n905_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n903_), .A2(new_n906_), .ZN(G1354gat));
  OAI21_X1  g706(.A(G218gat), .B1(new_n891_), .B2(new_n332_), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n329_), .A2(G218gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n891_), .B2(new_n909_), .ZN(G1355gat));
endmodule


