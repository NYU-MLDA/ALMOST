//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_;
  NOR3_X1   g000(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT65), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT6), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n203_), .A2(new_n204_), .A3(new_n206_), .A4(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G85gat), .B(G92gat), .Z(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT67), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT8), .B1(new_n208_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT66), .B1(new_n213_), .B2(KEYINPUT8), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n206_), .A2(new_n207_), .ZN(new_n215_));
  AOI211_X1 g014(.A(new_n210_), .B(new_n214_), .C1(new_n215_), .C2(new_n203_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G85gat), .A3(G92gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n206_), .A2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT64), .B(G106gat), .Z(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT10), .B(G99gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n209_), .A2(KEYINPUT9), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n217_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G71gat), .B(G78gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n227_), .B1(new_n230_), .B2(KEYINPUT11), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n228_), .B(KEYINPUT68), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT11), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(KEYINPUT11), .A3(new_n227_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n226_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT12), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n225_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n217_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n235_), .A2(new_n236_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT70), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n242_), .A2(new_n245_), .A3(KEYINPUT12), .A4(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G230gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n225_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n212_), .A2(new_n216_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n246_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n240_), .A2(new_n248_), .A3(new_n249_), .A4(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n238_), .A2(new_n252_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n249_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G120gat), .B(G148gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT5), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G176gat), .B(G204gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n257_), .B(new_n261_), .Z(new_n262_));
  OR2_X1    g061(.A1(new_n262_), .A2(KEYINPUT13), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(KEYINPUT13), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G127gat), .B(G155gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT16), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G183gat), .B(G211gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT17), .ZN(new_n272_));
  INV_X1    g071(.A(G1gat), .ZN(new_n273_));
  INV_X1    g072(.A(G8gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT14), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n275_), .A2(KEYINPUT75), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(KEYINPUT75), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G15gat), .B(G22gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G8gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n276_), .A2(new_n282_), .A3(new_n277_), .A4(new_n278_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G231gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(new_n246_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n288_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n272_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n242_), .A2(new_n247_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(new_n286_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n271_), .A2(KEYINPUT17), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT76), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT78), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G190gat), .B(G218gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G134gat), .B(G162gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT36), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G29gat), .B(G36gat), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n304_), .A2(KEYINPUT72), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(KEYINPUT72), .ZN(new_n306_));
  XOR2_X1   g105(.A(G43gat), .B(G50gat), .Z(new_n307_));
  OR3_X1    g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n307_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n217_), .A2(new_n311_), .A3(new_n225_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n251_), .A2(KEYINPUT73), .A3(new_n311_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G232gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT34), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT35), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT15), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n310_), .B(new_n323_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n245_), .A2(new_n324_), .B1(new_n320_), .B2(new_n319_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n316_), .A2(new_n322_), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n322_), .B1(new_n316_), .B2(new_n325_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n302_), .A2(KEYINPUT36), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n326_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n316_), .A2(new_n325_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n321_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n316_), .A2(new_n322_), .A3(new_n325_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n328_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n303_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT37), .B1(new_n330_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n329_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n332_), .A2(new_n328_), .A3(new_n333_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n339_), .A2(new_n340_), .B1(KEYINPUT36), .B2(new_n302_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT37), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n340_), .B2(KEYINPUT74), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n338_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n299_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n267_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT79), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n351_));
  INV_X1    g150(.A(G197gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(G204gat), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT93), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(G197gat), .A3(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n353_), .A2(KEYINPUT93), .A3(G204gat), .A4(new_n354_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n357_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G211gat), .B(G218gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT21), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n357_), .A2(new_n360_), .A3(new_n361_), .A4(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n363_), .ZN(new_n369_));
  AND2_X1   g168(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n352_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT92), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n353_), .A2(new_n354_), .ZN(new_n374_));
  INV_X1    g173(.A(G204gat), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n372_), .A2(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n358_), .A2(new_n359_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(KEYINPUT92), .A3(new_n352_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n364_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n366_), .B1(new_n369_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT2), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT88), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT88), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n397_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n388_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n389_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(new_n394_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n386_), .B1(new_n385_), .B2(KEYINPUT1), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT1), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n383_), .A2(new_n408_), .A3(new_n384_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n406_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT29), .B1(new_n403_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(G228gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(G228gat), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n412_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n380_), .A2(new_n411_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n380_), .B2(new_n411_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n350_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT95), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n388_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n396_), .A2(new_n398_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n391_), .A2(new_n392_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR4_X1   g226(.A1(KEYINPUT87), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n401_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n424_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n384_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT1), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(new_n409_), .A3(new_n387_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n405_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n431_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n437_), .A2(KEYINPUT29), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G22gat), .B(G50gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT28), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n438_), .B(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n380_), .A2(new_n411_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n417_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n380_), .A2(new_n411_), .A3(new_n418_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n350_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n423_), .A2(new_n441_), .B1(new_n421_), .B2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n421_), .A2(new_n446_), .A3(new_n441_), .A4(KEYINPUT95), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G225gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G127gat), .B(G134gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G120gat), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n452_), .A2(new_n453_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n403_), .B2(new_n410_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n452_), .B(new_n453_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n431_), .A2(new_n436_), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(KEYINPUT4), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT4), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n437_), .A2(new_n461_), .A3(new_n456_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n451_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G1gat), .B(G29gat), .ZN(new_n464_));
  INV_X1    g263(.A(G85gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT0), .B(G57gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n457_), .A2(new_n459_), .B1(G225gat), .B2(G233gat), .ZN(new_n469_));
  OR3_X1    g268(.A1(new_n463_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n463_), .B2(new_n469_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n456_), .A2(KEYINPUT31), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT31), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n458_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(G99gat), .ZN(new_n479_));
  INV_X1    g278(.A(G99gat), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n474_), .A2(new_n476_), .A3(new_n477_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G227gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(G71gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n479_), .A2(new_n485_), .A3(new_n481_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G15gat), .B(G43gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT83), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT30), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(G183gat), .ZN(new_n494_));
  INV_X1    g293(.A(G190gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT23), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT23), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(G183gat), .A3(G190gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n497_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(new_n495_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(G169gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT25), .B(G183gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT26), .B(G190gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(G169gat), .ZN(new_n510_));
  INV_X1    g309(.A(G176gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G169gat), .A2(G176gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(KEYINPUT24), .A3(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n512_), .A2(KEYINPUT24), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n509_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT81), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n496_), .A2(new_n498_), .A3(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT81), .B(KEYINPUT23), .C1(new_n494_), .C2(new_n495_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI22_X1  g319(.A1(new_n503_), .A2(new_n506_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT85), .Z(new_n522_));
  INV_X1    g321(.A(new_n492_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n487_), .A2(new_n488_), .A3(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n493_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n522_), .B1(new_n493_), .B2(new_n524_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n473_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT99), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n529_));
  INV_X1    g328(.A(new_n365_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n361_), .A2(new_n360_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n531_), .B2(new_n357_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n368_), .A2(new_n363_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n372_), .A2(new_n373_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n374_), .A2(new_n375_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n378_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT21), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n532_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n516_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n500_), .A2(new_n501_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n518_), .A2(new_n519_), .A3(new_n502_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n540_), .A2(new_n542_), .B1(new_n505_), .B2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n529_), .B1(new_n539_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G226gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT19), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT96), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n380_), .A2(new_n549_), .A3(new_n521_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n380_), .B2(new_n521_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n545_), .B(new_n548_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT20), .B1(new_n380_), .B2(new_n521_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n538_), .A2(new_n368_), .A3(new_n363_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n544_), .B1(new_n554_), .B2(new_n366_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n547_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G8gat), .B(G36gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT18), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G64gat), .B(G92gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  NAND3_X1  g359(.A1(new_n552_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT27), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n545_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n547_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n553_), .A2(new_n555_), .A3(new_n547_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n560_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n560_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n543_), .A2(new_n505_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n516_), .B2(new_n541_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT20), .B(new_n548_), .C1(new_n380_), .C2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n551_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n380_), .A2(new_n549_), .A3(new_n521_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n521_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n529_), .B1(new_n539_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n380_), .A2(new_n571_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n548_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n569_), .B1(new_n575_), .B2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT27), .B1(new_n580_), .B2(new_n561_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n528_), .B1(new_n568_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT27), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n552_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n560_), .B1(new_n552_), .B2(new_n556_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n583_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n565_), .B1(new_n563_), .B2(new_n547_), .ZN(new_n587_));
  OAI211_X1 g386(.A(KEYINPUT27), .B(new_n561_), .C1(new_n587_), .C2(new_n560_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n588_), .A3(KEYINPUT99), .ZN(new_n589_));
  AOI211_X1 g388(.A(new_n450_), .B(new_n527_), .C1(new_n582_), .C2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n588_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n445_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n441_), .B1(new_n593_), .B2(KEYINPUT95), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n421_), .A2(new_n446_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n473_), .A2(new_n448_), .A3(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n591_), .B1(new_n592_), .B2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n447_), .A2(new_n472_), .A3(new_n449_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n599_), .A2(KEYINPUT98), .A3(new_n586_), .A4(new_n588_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n560_), .A2(KEYINPUT32), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n552_), .A2(new_n556_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n472_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n587_), .A2(new_n601_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n471_), .A2(KEYINPUT33), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n607_), .B(new_n468_), .C1(new_n463_), .C2(new_n469_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  AND4_X1   g408(.A1(G225gat), .A2(new_n457_), .A3(G233gat), .A4(new_n459_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n468_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n460_), .A2(new_n451_), .A3(new_n462_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT97), .B1(new_n580_), .B2(new_n561_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n580_), .A2(KEYINPUT97), .A3(new_n561_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n605_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n598_), .B(new_n600_), .C1(new_n618_), .C2(new_n450_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n525_), .A2(new_n526_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n590_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n324_), .A2(new_n284_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n310_), .A2(new_n284_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n310_), .B(new_n284_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT80), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(G113gat), .B(G141gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(G169gat), .B(G197gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n631_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n621_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n349_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n273_), .A3(new_n472_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n621_), .A2(new_n335_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n297_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n265_), .A2(new_n636_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n646_), .B2(new_n473_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n640_), .A2(new_n641_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n642_), .A2(new_n647_), .A3(new_n648_), .ZN(G1324gat));
  INV_X1    g448(.A(new_n582_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n589_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n639_), .A2(new_n274_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n646_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G8gat), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT100), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n655_), .A2(new_n659_), .A3(G8gat), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n657_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n658_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n653_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n653_), .B(new_n664_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  OAI21_X1  g467(.A(G15gat), .B1(new_n646_), .B2(new_n620_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT41), .Z(new_n670_));
  OR2_X1    g469(.A1(new_n620_), .A2(G15gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n638_), .B2(new_n671_), .ZN(G1326gat));
  INV_X1    g471(.A(new_n450_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G22gat), .B1(new_n646_), .B2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT42), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n673_), .A2(G22gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n638_), .B2(new_n676_), .ZN(G1327gat));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n265_), .A2(new_n298_), .A3(new_n636_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n598_), .A2(new_n600_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT97), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n683_), .A2(new_n617_), .A3(new_n613_), .A4(new_n609_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n603_), .A2(new_n604_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n450_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n620_), .B1(new_n681_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n527_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n673_), .B(new_n688_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n680_), .B1(new_n690_), .B2(new_n346_), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT43), .B(new_n345_), .C1(new_n687_), .C2(new_n689_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n679_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT104), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n263_), .A2(new_n264_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n635_), .A3(new_n299_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n621_), .B2(new_n345_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n690_), .A2(new_n680_), .A3(new_n346_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n695_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n694_), .B1(new_n700_), .B2(new_n704_), .ZN(new_n705_));
  AOI211_X1 g504(.A(KEYINPUT102), .B(new_n697_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n705_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT44), .B1(new_n693_), .B2(KEYINPUT102), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n700_), .A2(new_n704_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT103), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n472_), .B(new_n703_), .C1(new_n708_), .C2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G29gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n298_), .A2(new_n341_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n637_), .A2(new_n696_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(G29gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n472_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n678_), .B1(new_n713_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n717_), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT105), .B(new_n719_), .C1(new_n712_), .C2(G29gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1328gat));
  INV_X1    g520(.A(new_n652_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n695_), .B2(new_n702_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n723_), .B1(new_n708_), .B2(new_n711_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G36gat), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  INV_X1    g525(.A(G36gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n715_), .A2(new_n727_), .A3(new_n652_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT45), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n725_), .A2(KEYINPUT106), .A3(new_n726_), .A4(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n726_), .A2(KEYINPUT106), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n726_), .A2(KEYINPUT106), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n707_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n709_), .A2(KEYINPUT103), .A3(new_n710_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n727_), .B1(new_n735_), .B2(new_n723_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n729_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n731_), .B(new_n732_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n730_), .A2(new_n738_), .ZN(G1329gat));
  INV_X1    g538(.A(new_n620_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n735_), .A2(G43gat), .A3(new_n740_), .A4(new_n703_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G43gat), .B1(new_n715_), .B2(new_n740_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT47), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n741_), .A2(new_n746_), .A3(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1330gat));
  AOI21_X1  g547(.A(G50gat), .B1(new_n715_), .B2(new_n450_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n735_), .A2(new_n703_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n450_), .A2(G50gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(G1331gat));
  NOR3_X1   g551(.A1(new_n696_), .A2(new_n346_), .A3(new_n299_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n621_), .A2(new_n635_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G57gat), .B1(new_n756_), .B2(new_n472_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n298_), .A2(new_n636_), .ZN(new_n758_));
  NOR4_X1   g557(.A1(new_n267_), .A2(new_n621_), .A3(new_n335_), .A4(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n473_), .A2(KEYINPUT107), .ZN(new_n760_));
  MUX2_X1   g559(.A(KEYINPUT107), .B(new_n760_), .S(G57gat), .Z(new_n761_));
  AOI21_X1  g560(.A(new_n757_), .B1(new_n759_), .B2(new_n761_), .ZN(G1332gat));
  INV_X1    g561(.A(G64gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n759_), .B2(new_n652_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT48), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n756_), .A2(new_n763_), .A3(new_n652_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1333gat));
  AOI21_X1  g566(.A(new_n484_), .B1(new_n759_), .B2(new_n740_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT49), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n756_), .A2(new_n484_), .A3(new_n740_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1334gat));
  NAND2_X1  g570(.A1(new_n759_), .A2(new_n450_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G78gat), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT50), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n673_), .A2(G78gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n755_), .B2(new_n775_), .ZN(G1335gat));
  XNOR2_X1  g575(.A(new_n265_), .B(KEYINPUT71), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(new_n714_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(new_n754_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n465_), .A3(new_n472_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n265_), .A2(new_n299_), .A3(new_n636_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n691_), .A2(new_n692_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT108), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n781_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT109), .B(new_n781_), .C1(new_n783_), .C2(new_n785_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n473_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n780_), .B1(new_n790_), .B2(new_n465_), .ZN(G1336gat));
  INV_X1    g590(.A(G92gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n779_), .A2(new_n792_), .A3(new_n652_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n788_), .A2(new_n789_), .A3(new_n722_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n792_), .ZN(G1337gat));
  INV_X1    g594(.A(new_n222_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n779_), .A2(new_n740_), .A3(new_n796_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n788_), .A2(new_n789_), .A3(new_n620_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n480_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n797_), .C1(new_n798_), .C2(new_n480_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1338gat));
  NOR2_X1   g602(.A1(new_n673_), .A2(new_n221_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n778_), .A2(new_n754_), .A3(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT110), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n781_), .A2(new_n673_), .ZN(new_n807_));
  OAI21_X1  g606(.A(G106gat), .B1(new_n782_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n809_), .A2(KEYINPUT52), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(KEYINPUT52), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n806_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT53), .ZN(G1339gat));
  OR2_X1    g612(.A1(new_n257_), .A2(new_n261_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n625_), .A2(new_n628_), .A3(new_n634_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n634_), .B1(new_n626_), .B2(new_n624_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT113), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT114), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n622_), .A2(new_n623_), .A3(new_n627_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n818_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n814_), .B(new_n815_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n253_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n240_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n255_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n253_), .A2(new_n824_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n826_), .A2(KEYINPUT112), .A3(new_n255_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n825_), .A2(new_n829_), .A3(new_n830_), .A4(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n261_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n261_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(KEYINPUT115), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n261_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n836_), .A2(KEYINPUT115), .A3(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n823_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT58), .B(new_n823_), .C1(new_n835_), .C2(new_n838_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n841_), .A2(new_n346_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n635_), .A2(new_n814_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n836_), .A2(new_n837_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n833_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n815_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n262_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n341_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT57), .B(new_n341_), .C1(new_n846_), .C2(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n644_), .B1(new_n843_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n696_), .A2(new_n636_), .A3(new_n345_), .A4(new_n298_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(KEYINPUT54), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n758_), .A2(new_n265_), .A3(new_n346_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(KEYINPUT111), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n856_), .A2(KEYINPUT54), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n854_), .A2(new_n862_), .ZN(new_n863_));
  NOR4_X1   g662(.A1(new_n652_), .A2(new_n450_), .A3(new_n473_), .A4(new_n620_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT116), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G113gat), .B1(new_n867_), .B2(new_n635_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n299_), .B1(new_n843_), .B2(new_n853_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n862_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n865_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(KEYINPUT59), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n866_), .A2(KEYINPUT59), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n635_), .A2(G113gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT117), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n868_), .B1(new_n873_), .B2(new_n875_), .ZN(G1340gat));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n777_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G120gat), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n879_));
  AOI21_X1  g678(.A(G120gat), .B1(new_n265_), .B2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n879_), .B2(G120gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT118), .B1(new_n867_), .B2(new_n881_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n867_), .A2(KEYINPUT118), .A3(new_n881_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n878_), .B1(new_n882_), .B2(new_n883_), .ZN(G1341gat));
  INV_X1    g683(.A(G127gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n866_), .B2(new_n299_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n887_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n644_), .A2(new_n885_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n888_), .A2(new_n889_), .B1(new_n873_), .B2(new_n890_), .ZN(G1342gat));
  INV_X1    g690(.A(G134gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n866_), .B2(new_n341_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n894_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n345_), .A2(new_n892_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT121), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n895_), .A2(new_n896_), .B1(new_n873_), .B2(new_n898_), .ZN(G1343gat));
  NOR3_X1   g698(.A1(new_n652_), .A2(new_n673_), .A3(new_n473_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n863_), .A2(new_n620_), .A3(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n636_), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n267_), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g704(.A1(new_n901_), .A2(new_n299_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT61), .B(G155gat), .Z(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1346gat));
  INV_X1    g707(.A(G162gat), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n901_), .A2(new_n909_), .A3(new_n345_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n901_), .B2(new_n341_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n912_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n910_), .B1(new_n913_), .B2(new_n914_), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n722_), .A2(new_n527_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n450_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(new_n869_), .B2(new_n862_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n510_), .B1(new_n920_), .B2(new_n635_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT124), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n851_), .A2(new_n852_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n841_), .A2(new_n346_), .A3(new_n842_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n298_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n857_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n635_), .B(new_n918_), .C1(new_n926_), .C2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(G169gat), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n929_), .A2(new_n930_), .A3(KEYINPUT62), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n928_), .A2(new_n922_), .A3(G169gat), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n921_), .A2(KEYINPUT123), .A3(new_n922_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n923_), .A2(new_n931_), .A3(new_n934_), .A4(new_n935_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT22), .B(G169gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n920_), .A2(new_n635_), .A3(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1348gat));
  AOI21_X1  g738(.A(G176gat), .B1(new_n920_), .B2(new_n265_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n450_), .B1(new_n854_), .B2(new_n862_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n267_), .A2(new_n511_), .A3(new_n917_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(G1349gat));
  NAND3_X1  g742(.A1(new_n941_), .A2(new_n298_), .A3(new_n916_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n644_), .A2(new_n507_), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n944_), .A2(new_n494_), .B1(new_n920_), .B2(new_n945_), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n920_), .A2(new_n508_), .A3(new_n335_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n920_), .A2(new_n346_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n947_), .B1(new_n949_), .B2(new_n495_), .ZN(G1351gat));
  NOR2_X1   g749(.A1(new_n722_), .A2(new_n597_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n297_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n620_), .B(new_n951_), .C1(new_n952_), .C2(new_n927_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n953_), .A2(new_n636_), .ZN(new_n954_));
  XOR2_X1   g753(.A(KEYINPUT125), .B(G197gat), .Z(new_n955_));
  XNOR2_X1  g754(.A(new_n954_), .B(new_n955_), .ZN(G1352gat));
  OAI21_X1  g755(.A(new_n375_), .B1(new_n953_), .B2(new_n267_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n740_), .B1(new_n854_), .B2(new_n862_), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n958_), .A2(new_n377_), .A3(new_n777_), .A4(new_n951_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n959_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(KEYINPUT126), .ZN(G1353gat));
  NAND3_X1  g760(.A1(new_n958_), .A2(new_n297_), .A3(new_n951_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n963_));
  AND2_X1   g762(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n964_));
  NOR3_X1   g763(.A1(new_n962_), .A2(new_n963_), .A3(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n965_), .B1(new_n962_), .B2(new_n963_), .ZN(G1354gat));
  OAI21_X1  g765(.A(G218gat), .B1(new_n953_), .B2(new_n345_), .ZN(new_n967_));
  OR2_X1    g766(.A1(new_n341_), .A2(G218gat), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n967_), .B1(new_n953_), .B2(new_n968_), .ZN(G1355gat));
endmodule


