//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203_));
  XOR2_X1   g002(.A(G85gat), .B(G92gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT9), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT10), .B(G99gat), .Z(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(G85gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n205_), .A2(new_n208_), .A3(new_n213_), .A4(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G57gat), .B(G64gat), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n218_), .A2(KEYINPUT11), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(KEYINPUT11), .ZN(new_n220_));
  XOR2_X1   g019(.A(G71gat), .B(G78gat), .Z(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n220_), .A2(new_n221_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  INV_X1    g024(.A(new_n213_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n207_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n225_), .B(new_n204_), .C1(new_n226_), .C2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n231_), .B(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n213_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n225_), .B1(new_n237_), .B2(new_n204_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n232_), .B1(new_n238_), .B2(KEYINPUT67), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240_));
  AOI211_X1 g039(.A(new_n240_), .B(new_n225_), .C1(new_n237_), .C2(new_n204_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n217_), .B(new_n224_), .C1(new_n239_), .C2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n238_), .A2(KEYINPUT67), .ZN(new_n244_));
  INV_X1    g043(.A(new_n241_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n232_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n224_), .B1(new_n246_), .B2(new_n217_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n247_), .B2(KEYINPUT12), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G230gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n217_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n224_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT12), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n250_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AOI211_X1 g054(.A(KEYINPUT68), .B(KEYINPUT12), .C1(new_n251_), .C2(new_n252_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n248_), .B(new_n249_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(G230gat), .B(G233gat), .C1(new_n247_), .C2(new_n243_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G120gat), .B(G148gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(G176gat), .B(G204gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n257_), .A2(new_n258_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n264_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n203_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n257_), .A2(new_n258_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n263_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n257_), .A2(new_n258_), .A3(new_n264_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(KEYINPUT70), .A3(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n271_), .A3(KEYINPUT13), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT13), .B1(new_n267_), .B2(new_n271_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT71), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n267_), .A2(new_n271_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT13), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n276_), .B1(new_n279_), .B2(new_n272_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n202_), .B1(new_n275_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G15gat), .B(G22gat), .ZN(new_n282_));
  INV_X1    g081(.A(G1gat), .ZN(new_n283_));
  INV_X1    g082(.A(G8gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT14), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G1gat), .B(G8gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G231gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(new_n252_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G127gat), .B(G155gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT16), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G183gat), .B(G211gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT17), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n298_), .B(KEYINPUT78), .Z(new_n299_));
  AND2_X1   g098(.A1(new_n295_), .A2(new_n296_), .ZN(new_n300_));
  OR3_X1    g099(.A1(new_n291_), .A2(new_n297_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G29gat), .B(G36gat), .Z(new_n304_));
  XOR2_X1   g103(.A(G43gat), .B(G50gat), .Z(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT15), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n251_), .A2(new_n308_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n306_), .B(new_n217_), .C1(new_n239_), .C2(new_n241_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT35), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(new_n314_), .A3(new_n310_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G232gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n313_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(G190gat), .B(G218gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT74), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G134gat), .B(G162gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT36), .ZN(new_n325_));
  INV_X1    g124(.A(new_n318_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n311_), .A2(new_n312_), .A3(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n319_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n319_), .A2(new_n327_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n329_), .A2(KEYINPUT77), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n323_), .B(KEYINPUT36), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT75), .Z(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n329_), .B2(KEYINPUT77), .ZN(new_n333_));
  AOI211_X1 g132(.A(KEYINPUT37), .B(new_n328_), .C1(new_n330_), .C2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT37), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n319_), .B2(new_n327_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT76), .B1(new_n328_), .B2(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n336_), .A2(KEYINPUT76), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n335_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n303_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT79), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n338_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT37), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n328_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n335_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n303_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n341_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT71), .B1(new_n273_), .B2(new_n274_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n279_), .A2(new_n276_), .A3(new_n272_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(KEYINPUT72), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n281_), .A2(new_n349_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT100), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT25), .B(G183gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT26), .B(G190gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n356_), .A2(new_n357_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G183gat), .A2(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT23), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(G183gat), .A3(G190gat), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(G169gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n365_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n371_), .B(new_n372_), .C1(G183gat), .C2(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G71gat), .B(G99gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(G15gat), .B(G43gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n375_), .B(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G127gat), .B(G134gat), .Z(new_n380_));
  XOR2_X1   g179(.A(G113gat), .B(G120gat), .Z(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n379_), .B(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n385_), .B(KEYINPUT81), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT30), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT31), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n384_), .B(new_n388_), .Z(new_n389_));
  XOR2_X1   g188(.A(new_n389_), .B(KEYINPUT82), .Z(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT27), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT18), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT19), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G197gat), .ZN(new_n400_));
  INV_X1    g199(.A(G204gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G197gat), .A2(G204gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(KEYINPUT21), .A3(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G211gat), .B(G218gat), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G197gat), .A2(G204gat), .ZN(new_n407_));
  AND2_X1   g206(.A1(G197gat), .A2(G204gat), .ZN(new_n408_));
  AND2_X1   g207(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n409_));
  NOR2_X1   g208(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n410_));
  OAI22_X1  g209(.A1(new_n407_), .A2(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n402_), .A2(new_n403_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT86), .B(KEYINPUT21), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT87), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n406_), .A2(new_n413_), .A3(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT88), .B1(new_n404_), .B2(new_n405_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n406_), .A2(new_n418_), .A3(new_n413_), .A4(new_n416_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n360_), .B(KEYINPUT91), .ZN(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT22), .B(G169gat), .Z(new_n424_));
  OAI211_X1 g223(.A(new_n373_), .B(new_n423_), .C1(G176gat), .C2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n368_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n428_));
  INV_X1    g227(.A(new_n375_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(new_n422_), .B2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n427_), .B1(new_n430_), .B2(KEYINPUT90), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT90), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n375_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n432_), .B1(new_n433_), .B2(new_n428_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n399_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT87), .B1(new_n414_), .B2(new_n415_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n404_), .A2(new_n405_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n418_), .B1(new_n438_), .B2(new_n416_), .ZN(new_n439_));
  AND4_X1   g238(.A1(new_n418_), .A2(new_n406_), .A3(new_n413_), .A4(new_n416_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n426_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n420_), .A2(new_n375_), .A3(new_n421_), .ZN(new_n442_));
  AND4_X1   g241(.A1(KEYINPUT20), .A2(new_n441_), .A3(new_n399_), .A4(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n396_), .B1(new_n435_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n429_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n422_), .A2(new_n426_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n434_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AOI211_X1 g247(.A(new_n396_), .B(new_n443_), .C1(new_n448_), .C2(new_n398_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n444_), .B1(new_n449_), .B2(KEYINPUT92), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n443_), .B1(new_n448_), .B2(new_n398_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n396_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(KEYINPUT92), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n392_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n448_), .A2(new_n398_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n443_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n452_), .A3(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n426_), .B(KEYINPUT98), .ZN(new_n459_));
  INV_X1    g258(.A(new_n422_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT20), .B(new_n442_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n398_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n431_), .A2(new_n399_), .A3(new_n434_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(KEYINPUT27), .B(new_n458_), .C1(new_n464_), .C2(new_n452_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n455_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G155gat), .ZN(new_n468_));
  INV_X1    g267(.A(G162gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n469_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT2), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n472_), .A2(new_n473_), .B1(G141gat), .B2(G148gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(KEYINPUT84), .A2(KEYINPUT2), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n481_));
  INV_X1    g280(.A(G141gat), .ZN(new_n482_));
  INV_X1    g281(.A(G148gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(KEYINPUT85), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n485_));
  OAI22_X1  g284(.A1(KEYINPUT83), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n471_), .B1(new_n480_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT1), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n471_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n482_), .A2(new_n483_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G141gat), .A2(G148gat), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n470_), .B1(new_n488_), .B2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n470_), .A2(new_n489_), .A3(new_n491_), .A4(new_n492_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT29), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n460_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G228gat), .A2(G233gat), .ZN(new_n501_));
  INV_X1    g300(.A(G78gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(new_n207_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n500_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(new_n499_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT28), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G22gat), .B(G50gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n507_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n505_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n511_), .B2(new_n510_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n505_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n383_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n474_), .A2(new_n475_), .B1(new_n478_), .B2(new_n477_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n517_), .A2(new_n485_), .A3(new_n484_), .A4(new_n486_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n493_), .B1(new_n518_), .B2(new_n471_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n382_), .B(new_n496_), .C1(new_n519_), .C2(new_n470_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n516_), .A2(new_n520_), .A3(KEYINPUT4), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G225gat), .A2(G233gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT4), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n524_), .B(new_n383_), .C1(new_n495_), .C2(new_n497_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n516_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G1gat), .B(G29gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G57gat), .B(G85gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n467_), .A2(new_n515_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n515_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n452_), .A2(KEYINPUT32), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n464_), .A2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n451_), .A2(new_n542_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n543_), .A2(new_n537_), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n516_), .A2(new_n520_), .A3(new_n523_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n533_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT95), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n546_), .A2(new_n549_), .A3(new_n533_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n521_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n552_), .A2(KEYINPUT96), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(KEYINPUT96), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT33), .B1(new_n528_), .B2(new_n533_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n526_), .A2(new_n557_), .A3(new_n535_), .A4(new_n527_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n554_), .A2(new_n555_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT92), .B1(new_n451_), .B2(new_n452_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n451_), .A2(new_n452_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n560_), .B1(new_n563_), .B2(new_n453_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n458_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n566_), .A2(new_n560_), .A3(new_n453_), .A4(new_n444_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n559_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n545_), .B1(new_n569_), .B2(KEYINPUT97), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n556_), .A2(new_n558_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n521_), .A2(new_n525_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n573_), .A2(new_n522_), .B1(new_n547_), .B2(KEYINPUT95), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n574_), .B2(new_n550_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n571_), .B1(new_n575_), .B2(new_n553_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT93), .B1(new_n450_), .B2(new_n454_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(new_n567_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n541_), .B1(new_n570_), .B2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n540_), .B1(new_n581_), .B2(KEYINPUT99), .ZN(new_n582_));
  INV_X1    g381(.A(new_n545_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n584_));
  AOI211_X1 g383(.A(KEYINPUT97), .B(new_n576_), .C1(new_n577_), .C2(new_n567_), .ZN(new_n585_));
  OAI211_X1 g384(.A(KEYINPUT99), .B(new_n515_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n391_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n515_), .A2(new_n466_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n589_), .A2(new_n538_), .A3(new_n389_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n306_), .B(new_n288_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT80), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(G229gat), .A3(G233gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n307_), .A2(new_n288_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n306_), .A2(new_n288_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G113gat), .B(G141gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G169gat), .B(G197gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  XNOR2_X1  g402(.A(new_n600_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n355_), .B1(new_n592_), .B2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n515_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n539_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n390_), .B1(new_n609_), .B2(new_n586_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n355_), .B(new_n605_), .C1(new_n610_), .C2(new_n590_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n354_), .B1(new_n606_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n607_), .A2(new_n608_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n586_), .A3(new_n540_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n590_), .B1(new_n618_), .B2(new_n391_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT100), .B1(new_n619_), .B2(new_n604_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n611_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(KEYINPUT101), .A3(new_n354_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n615_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT101), .B1(new_n621_), .B2(new_n354_), .ZN(new_n624_));
  AOI211_X1 g423(.A(new_n614_), .B(new_n353_), .C1(new_n620_), .C2(new_n611_), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT102), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n537_), .A2(G1gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n623_), .A2(new_n626_), .A3(KEYINPUT103), .A4(new_n627_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(KEYINPUT38), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT104), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n630_), .A2(new_n634_), .A3(KEYINPUT38), .A4(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT38), .B1(new_n630_), .B2(new_n631_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n275_), .A2(new_n280_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n605_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT105), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(new_n303_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n619_), .A2(new_n344_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n283_), .B1(new_n644_), .B2(new_n538_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n637_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n636_), .A2(new_n646_), .ZN(G1324gat));
  NOR2_X1   g446(.A1(new_n466_), .A2(G8gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n623_), .A2(new_n626_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n623_), .A2(new_n626_), .A3(KEYINPUT106), .A4(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G8gat), .B1(new_n643_), .B2(new_n466_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT39), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(G8gat), .C1(new_n643_), .C2(new_n466_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n653_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n653_), .A2(new_n658_), .A3(KEYINPUT40), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n643_), .B2(new_n391_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT41), .Z(new_n665_));
  NOR2_X1   g464(.A1(new_n624_), .A2(new_n625_), .ZN(new_n666_));
  INV_X1    g465(.A(G15gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n390_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(G1326gat));
  OAI21_X1  g468(.A(G22gat), .B1(new_n643_), .B2(new_n515_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT42), .ZN(new_n671_));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n666_), .A2(new_n672_), .A3(new_n541_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(G1327gat));
  INV_X1    g473(.A(new_n344_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n303_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n621_), .A2(new_n638_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G29gat), .B1(new_n678_), .B2(new_n538_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n346_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT43), .B1(new_n592_), .B2(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(new_n303_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n592_), .A2(KEYINPUT43), .A3(new_n680_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n640_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n685_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n538_), .A2(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n679_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  NOR3_X1   g489(.A1(new_n677_), .A2(G36gat), .A3(new_n466_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT45), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n686_), .A2(new_n467_), .A3(new_n687_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G36gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(G1329gat));
  INV_X1    g496(.A(G43gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n389_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n686_), .A2(new_n687_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT107), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n686_), .A2(new_n702_), .A3(new_n687_), .A4(new_n699_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n698_), .B1(new_n677_), .B2(new_n391_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n701_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT47), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n701_), .A2(new_n707_), .A3(new_n703_), .A4(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1330gat));
  AOI21_X1  g508(.A(G50gat), .B1(new_n678_), .B2(new_n541_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n541_), .A2(G50gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n688_), .B2(new_n711_), .ZN(G1331gat));
  NOR2_X1   g511(.A1(new_n619_), .A2(new_n605_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n638_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n349_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(G57gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n538_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n281_), .A2(new_n352_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n642_), .A2(new_n604_), .A3(new_n303_), .A4(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G57gat), .B1(new_n719_), .B2(new_n537_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(G1332gat));
  OAI21_X1  g520(.A(G64gat), .B1(new_n719_), .B2(new_n466_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT48), .ZN(new_n723_));
  INV_X1    g522(.A(G64gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n715_), .A2(new_n724_), .A3(new_n467_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n719_), .B2(new_n391_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT49), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n391_), .A2(G71gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT108), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n715_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n731_), .ZN(G1334gat));
  OAI21_X1  g531(.A(G78gat), .B1(new_n719_), .B2(new_n515_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT50), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n715_), .A2(new_n502_), .A3(new_n541_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1335gat));
  NOR2_X1   g535(.A1(new_n638_), .A2(new_n605_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n682_), .A2(new_n683_), .A3(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n537_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n713_), .A2(new_n718_), .A3(new_n676_), .ZN(new_n740_));
  INV_X1    g539(.A(G85gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n538_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n740_), .B2(new_n467_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n738_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n467_), .A2(new_n214_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT109), .Z(new_n747_));
  AOI21_X1  g546(.A(new_n744_), .B1(new_n745_), .B2(new_n747_), .ZN(G1337gat));
  AOI21_X1  g547(.A(new_n228_), .B1(new_n745_), .B2(new_n390_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n389_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n206_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n740_), .B2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n752_), .B(new_n753_), .Z(G1338gat));
  NAND3_X1  g553(.A1(new_n740_), .A2(new_n207_), .A3(new_n541_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n745_), .A2(new_n541_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(G106gat), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n757_), .B1(new_n756_), .B2(G106gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT53), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n755_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1339gat));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT59), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n346_), .A2(new_n604_), .A3(new_n303_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n273_), .A2(new_n274_), .ZN(new_n769_));
  OR3_X1    g568(.A1(new_n768_), .A2(new_n769_), .A3(KEYINPUT54), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT54), .B1(new_n768_), .B2(new_n769_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n248_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n249_), .B1(new_n774_), .B2(KEYINPUT112), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n248_), .B(new_n776_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n775_), .A2(new_n777_), .B1(new_n778_), .B2(new_n257_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n242_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n255_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n253_), .A2(new_n250_), .A3(new_n254_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n783_), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n249_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n257_), .B2(new_n778_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n779_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n263_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT56), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n788_), .A2(new_n791_), .A3(new_n263_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n790_), .A2(new_n605_), .A3(new_n270_), .A4(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n603_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n600_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n594_), .A2(new_n597_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n794_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n797_), .A2(KEYINPUT114), .ZN(new_n798_));
  AND4_X1   g597(.A1(G229gat), .A2(new_n596_), .A3(G233gat), .A4(new_n598_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n797_), .B2(KEYINPUT114), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n795_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n267_), .A2(new_n271_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n793_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n675_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n344_), .B1(new_n793_), .B2(new_n802_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT57), .B1(new_n808_), .B2(KEYINPUT115), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n265_), .B1(new_n789_), .B2(KEYINPUT56), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n801_), .A3(new_n792_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n810_), .A2(KEYINPUT58), .A3(new_n801_), .A4(new_n792_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n680_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n807_), .A2(new_n809_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n773_), .B1(new_n816_), .B2(new_n302_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n767_), .B1(new_n817_), .B2(KEYINPUT116), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n589_), .A2(new_n389_), .A3(new_n537_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n816_), .A2(new_n302_), .ZN(new_n823_));
  AOI221_X4 g622(.A(new_n820_), .B1(KEYINPUT116), .B2(new_n767_), .C1(new_n823_), .C2(new_n772_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n605_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G113gat), .ZN(new_n826_));
  INV_X1    g625(.A(new_n817_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n819_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n828_), .A2(G113gat), .A3(new_n604_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n766_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n831_));
  AOI211_X1 g630(.A(KEYINPUT117), .B(new_n829_), .C1(new_n825_), .C2(G113gat), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1340gat));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n638_), .B2(KEYINPUT60), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT118), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n821_), .B(new_n836_), .C1(KEYINPUT60), .C2(new_n834_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(KEYINPUT119), .Z(new_n838_));
  OR2_X1    g637(.A1(new_n822_), .A2(new_n824_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n839_), .A2(new_n718_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n840_), .B2(new_n834_), .ZN(G1341gat));
  INV_X1    g640(.A(G127gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n821_), .A2(new_n842_), .A3(new_n303_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n839_), .A2(new_n303_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(G1342gat));
  AOI21_X1  g644(.A(G134gat), .B1(new_n821_), .B2(new_n344_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n680_), .A2(G134gat), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT120), .Z(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n839_), .B2(new_n848_), .ZN(G1343gat));
  NOR3_X1   g648(.A1(new_n817_), .A2(new_n390_), .A3(new_n515_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n467_), .A2(new_n537_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n604_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n482_), .ZN(G1344gat));
  INV_X1    g653(.A(new_n718_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n852_), .A2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(new_n483_), .ZN(G1345gat));
  OR3_X1    g656(.A1(new_n852_), .A2(KEYINPUT121), .A3(new_n302_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT121), .B1(new_n852_), .B2(new_n302_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1346gat));
  INV_X1    g662(.A(new_n852_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G162gat), .B1(new_n864_), .B2(new_n344_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n680_), .A2(G162gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT122), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n864_), .B2(new_n867_), .ZN(G1347gat));
  NOR2_X1   g667(.A1(new_n466_), .A2(new_n538_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n869_), .A2(new_n390_), .A3(new_n515_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n827_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n605_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n424_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n873_), .A2(G169gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(KEYINPUT62), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(KEYINPUT62), .B2(new_n875_), .ZN(G1348gat));
  OR3_X1    g676(.A1(new_n871_), .A2(G176gat), .A3(new_n638_), .ZN(new_n878_));
  OAI21_X1  g677(.A(G176gat), .B1(new_n871_), .B2(new_n855_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1349gat));
  NOR2_X1   g679(.A1(new_n871_), .A2(new_n302_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n356_), .B1(new_n882_), .B2(G183gat), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  OR2_X1    g683(.A1(KEYINPUT123), .A2(G183gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n881_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n871_), .B2(new_n346_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n344_), .A2(new_n357_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n871_), .B2(new_n890_), .ZN(G1351gat));
  NAND2_X1  g690(.A1(new_n850_), .A2(new_n869_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n604_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n400_), .ZN(G1352gat));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n855_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n401_), .ZN(G1353gat));
  NOR3_X1   g695(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n897_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n892_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n303_), .A2(new_n902_), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT125), .Z(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(new_n905_));
  MUX2_X1   g704(.A(new_n897_), .B(new_n900_), .S(new_n905_), .Z(G1354gat));
  INV_X1    g705(.A(G218gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n901_), .A2(new_n907_), .A3(new_n344_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n892_), .A2(new_n346_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n907_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n908_), .B(KEYINPUT127), .C1(new_n909_), .C2(new_n907_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1355gat));
endmodule


