//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT35), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT10), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n219_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT65), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n211_), .B(new_n217_), .C1(new_n223_), .C2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n219_), .A2(new_n221_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(new_n213_), .A3(new_n215_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AOI211_X1 g030(.A(KEYINPUT8), .B(new_n227_), .C1(new_n231_), .C2(new_n211_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n211_), .A2(new_n230_), .A3(new_n229_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n227_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n226_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT66), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n226_), .B(new_n239_), .C1(new_n232_), .C2(new_n236_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n206_), .B1(new_n241_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT73), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(KEYINPUT73), .B(new_n206_), .C1(new_n241_), .C2(new_n247_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n246_), .B(KEYINPUT15), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n237_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT72), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n251_), .A3(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n204_), .A2(new_n205_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n248_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n258_), .B(new_n253_), .C1(new_n205_), .C2(new_n204_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G134gat), .B(G162gat), .Z(new_n261_));
  XNOR2_X1  g060(.A(G190gat), .B(G218gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT36), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n263_), .A2(new_n264_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n260_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n257_), .A2(new_n264_), .A3(new_n263_), .A4(new_n259_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT74), .B(KEYINPUT37), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G15gat), .B(G22gat), .ZN(new_n276_));
  INV_X1    g075(.A(G1gat), .ZN(new_n277_));
  INV_X1    g076(.A(G8gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT14), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G8gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT75), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G231gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G71gat), .B(G78gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(G57gat), .B(G64gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n286_), .B1(KEYINPUT11), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n287_), .B2(KEYINPUT11), .ZN(new_n290_));
  INV_X1    g089(.A(G64gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G57gat), .ZN(new_n292_));
  INV_X1    g091(.A(G57gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G64gat), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n292_), .A2(new_n294_), .A3(new_n289_), .A4(KEYINPUT11), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n288_), .B1(new_n290_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(new_n294_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT11), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT67), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n299_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(new_n286_), .A4(new_n295_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n285_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n285_), .A2(new_n303_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G127gat), .B(G155gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(G183gat), .B(G211gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT17), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n304_), .A2(new_n305_), .A3(KEYINPUT77), .A4(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n304_), .A2(new_n305_), .A3(new_n311_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n310_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT17), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n312_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n275_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT78), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  INV_X1    g123(.A(G176gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OR3_X1    g125(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT82), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n329_), .B1(new_n330_), .B2(G183gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(G190gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT25), .B(G183gat), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n331_), .B(new_n332_), .C1(new_n333_), .C2(new_n329_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT23), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n328_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n335_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n339_), .B2(new_n335_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G169gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT84), .ZN(new_n347_));
  XOR2_X1   g146(.A(G71gat), .B(G99gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n345_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G15gat), .B(G43gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT83), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT30), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n353_), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT85), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G127gat), .B(G134gat), .Z(new_n357_));
  XOR2_X1   g156(.A(G113gat), .B(G120gat), .Z(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  XOR2_X1   g158(.A(new_n359_), .B(KEYINPUT31), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n354_), .A2(KEYINPUT85), .A3(new_n355_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G1gat), .B(G29gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G85gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G57gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G141gat), .ZN(new_n371_));
  INV_X1    g170(.A(G148gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G141gat), .A2(G148gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT2), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G155gat), .ZN(new_n379_));
  INV_X1    g178(.A(G162gat), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n378_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT1), .B1(new_n379_), .B2(new_n380_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT1), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(G155gat), .A3(G162gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n388_), .A3(new_n384_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n376_), .A3(new_n373_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n390_), .A2(new_n391_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n385_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n359_), .ZN(new_n396_));
  OR3_X1    g195(.A1(new_n394_), .A2(KEYINPUT100), .A3(new_n359_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n359_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n385_), .B(new_n398_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT100), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(KEYINPUT99), .A3(new_n359_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT99), .B1(new_n394_), .B2(new_n359_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n397_), .B(new_n400_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n370_), .B(new_n396_), .C1(new_n404_), .C2(new_n395_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n397_), .A2(new_n400_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n401_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n369_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n368_), .B1(new_n405_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n405_), .A2(new_n368_), .A3(new_n409_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n364_), .A2(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n394_), .A2(KEYINPUT29), .ZN(new_n415_));
  XOR2_X1   g214(.A(G22gat), .B(G50gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT28), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n415_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n419_), .B(KEYINPUT92), .Z(new_n420_));
  INV_X1    g219(.A(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT87), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(G228gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(G228gat), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(KEYINPUT91), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT88), .B(G197gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(G204gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(G197gat), .B2(G204gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(G211gat), .B(G218gat), .Z(new_n431_));
  AND2_X1   g230(.A1(new_n431_), .A2(KEYINPUT90), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT21), .B1(new_n431_), .B2(KEYINPUT90), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT21), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n428_), .A2(G204gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n436_), .B1(G197gat), .B2(G204gat), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n431_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n435_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n437_), .A2(new_n440_), .A3(new_n435_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n434_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n394_), .A2(KEYINPUT29), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n427_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n434_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n443_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n447_), .B1(new_n448_), .B2(new_n441_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n394_), .A2(KEYINPUT29), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n425_), .B(KEYINPUT91), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n420_), .B1(new_n446_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n418_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT94), .ZN(new_n456_));
  INV_X1    g255(.A(new_n452_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n426_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n420_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(new_n453_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT94), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n462_), .B(new_n418_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n456_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n461_), .B1(new_n456_), .B2(new_n463_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G8gat), .B(G36gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT18), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G64gat), .B(G92gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n338_), .A2(KEYINPUT96), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n336_), .A2(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n473_), .A2(new_n343_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n341_), .A2(KEYINPUT96), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n333_), .A2(new_n332_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n476_), .A2(new_n336_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n474_), .A2(new_n475_), .B1(new_n328_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n444_), .A2(KEYINPUT98), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n449_), .B2(new_n345_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G226gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT19), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n447_), .B(new_n478_), .C1(new_n448_), .C2(new_n441_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT98), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n479_), .A2(new_n481_), .A3(new_n484_), .A4(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n483_), .B(KEYINPUT95), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n478_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n480_), .B1(new_n449_), .B2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n337_), .A2(new_n344_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n447_), .B(new_n493_), .C1(new_n448_), .C2(new_n441_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n490_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n488_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n494_), .B(KEYINPUT20), .C1(new_n444_), .C2(new_n478_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n489_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(KEYINPUT97), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n471_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(new_n496_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(KEYINPUT97), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n470_), .A4(new_n488_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT27), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n481_), .A2(new_n485_), .ZN(new_n507_));
  OAI22_X1  g306(.A1(new_n507_), .A2(new_n484_), .B1(new_n489_), .B2(new_n498_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n508_), .B2(new_n471_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n505_), .A2(new_n506_), .B1(new_n504_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n414_), .A2(new_n466_), .A3(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(KEYINPUT32), .A3(new_n470_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n470_), .A2(KEYINPUT32), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT102), .Z(new_n514_));
  NAND4_X1  g313(.A1(new_n502_), .A2(new_n503_), .A3(new_n488_), .A4(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n412_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n512_), .B(new_n515_), .C1(new_n516_), .C2(new_n410_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n369_), .B(new_n396_), .C1(new_n404_), .C2(new_n395_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT101), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n406_), .A2(KEYINPUT4), .A3(new_n408_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT101), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n369_), .A4(new_n396_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n404_), .A2(new_n369_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(new_n368_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n519_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT33), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n412_), .A2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n405_), .A2(KEYINPUT33), .A3(new_n368_), .A4(new_n409_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n517_), .B1(new_n526_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n461_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n459_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT93), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n462_), .B1(new_n534_), .B2(new_n418_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n463_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n532_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n456_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n413_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n531_), .A2(new_n466_), .B1(new_n539_), .B2(new_n510_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n364_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n511_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n303_), .A2(KEYINPUT12), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n211_), .A2(new_n217_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT65), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n224_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT9), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT64), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT64), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT9), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n218_), .B1(new_n551_), .B2(new_n221_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n544_), .B1(new_n546_), .B2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n208_), .A2(new_n210_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n229_), .A2(new_n230_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n235_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT8), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n234_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n553_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT68), .B1(new_n543_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT12), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT68), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n237_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n303_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n238_), .A2(new_n566_), .A3(new_n240_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n565_), .B(new_n567_), .C1(KEYINPUT12), .C2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT69), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n563_), .B1(new_n237_), .B2(new_n562_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n237_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n567_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT12), .B1(new_n241_), .B2(new_n303_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT69), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n576_), .A2(new_n578_), .A3(new_n579_), .A4(new_n570_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n567_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n571_), .B1(new_n581_), .B2(new_n568_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n572_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G120gat), .B(G148gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n572_), .A2(new_n580_), .A3(new_n582_), .A4(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(KEYINPUT71), .B2(KEYINPUT13), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n282_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n246_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n247_), .A2(new_n282_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT79), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(G229gat), .A3(G233gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n252_), .A2(new_n282_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n598_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(G113gat), .B(G141gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT80), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G169gat), .B(G197gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n602_), .A2(new_n605_), .A3(new_n610_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(KEYINPUT81), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT81), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n596_), .B1(new_n614_), .B2(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n542_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n321_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n413_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n620_), .A2(G1gat), .A3(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n622_), .A2(KEYINPUT38), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(KEYINPUT38), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n414_), .A2(new_n466_), .A3(new_n510_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n531_), .A2(new_n466_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n539_), .A2(new_n510_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n625_), .B1(new_n628_), .B2(new_n364_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n615_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n596_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n319_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n269_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n629_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n635_), .B2(new_n621_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n623_), .A2(new_n624_), .A3(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(new_n510_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n634_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT103), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n634_), .A2(new_n641_), .A3(new_n638_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(G8gat), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(KEYINPUT104), .A3(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n640_), .A2(G8gat), .A3(new_n642_), .A4(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n321_), .A2(new_n619_), .A3(new_n278_), .A4(new_n638_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n645_), .A2(KEYINPUT40), .A3(new_n647_), .A4(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n635_), .B2(new_n364_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT41), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n620_), .A2(G15gat), .A3(new_n364_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1326gat));
  OAI21_X1  g456(.A(G22gat), .B1(new_n635_), .B2(new_n466_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT42), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n466_), .A2(G22gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n620_), .B2(new_n660_), .ZN(G1327gat));
  INV_X1    g460(.A(new_n319_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n631_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n664_), .B1(new_n629_), .B2(new_n275_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n541_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n274_), .B1(new_n668_), .B2(new_n625_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n664_), .A3(KEYINPUT43), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n663_), .B1(new_n667_), .B2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n663_), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT105), .B(new_n666_), .C1(new_n542_), .C2(new_n274_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT43), .B1(new_n669_), .B2(new_n664_), .ZN(new_n676_));
  OAI211_X1 g475(.A(KEYINPUT44), .B(new_n674_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n673_), .A2(new_n413_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G29gat), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n269_), .A2(new_n319_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n542_), .A2(new_n618_), .A3(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n621_), .A2(G29gat), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT107), .Z(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n681_), .B2(new_n683_), .ZN(G1328gat));
  OAI211_X1 g483(.A(new_n638_), .B(new_n677_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n510_), .A2(G36gat), .ZN(new_n687_));
  OR3_X1    g486(.A1(new_n681_), .A2(KEYINPUT108), .A3(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT108), .B1(new_n681_), .B2(new_n687_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(KEYINPUT45), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT45), .B1(new_n688_), .B2(new_n689_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n686_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n686_), .A2(KEYINPUT46), .A3(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1329gat));
  AND2_X1   g496(.A1(new_n541_), .A2(G43gat), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n677_), .B(new_n698_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT109), .B(G43gat), .Z(new_n700_));
  OAI21_X1  g499(.A(new_n700_), .B1(new_n681_), .B2(new_n364_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(G1330gat));
  INV_X1    g503(.A(new_n466_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n673_), .A2(G50gat), .A3(new_n705_), .A4(new_n677_), .ZN(new_n706_));
  INV_X1    g505(.A(G50gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n707_), .B1(new_n681_), .B2(new_n466_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1331gat));
  INV_X1    g508(.A(new_n596_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n319_), .A2(new_n617_), .A3(new_n614_), .ZN(new_n711_));
  OR4_X1    g510(.A1(new_n633_), .A2(new_n629_), .A3(new_n710_), .A4(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G57gat), .B1(new_n712_), .B2(new_n621_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n321_), .A2(new_n596_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n629_), .A2(new_n615_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n413_), .A2(new_n293_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(G1332gat));
  OAI21_X1  g517(.A(G64gat), .B1(new_n712_), .B2(new_n510_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n638_), .A2(new_n291_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n716_), .B2(new_n722_), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n712_), .B2(new_n364_), .ZN(new_n724_));
  XOR2_X1   g523(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n364_), .A2(G71gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n716_), .B2(new_n727_), .ZN(G1334gat));
  OAI21_X1  g527(.A(G78gat), .B1(new_n712_), .B2(new_n466_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT50), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n466_), .A2(G78gat), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT113), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n716_), .B2(new_n732_), .ZN(G1335gat));
  NAND3_X1  g532(.A1(new_n715_), .A2(new_n596_), .A3(new_n680_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(G85gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n413_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n667_), .A2(new_n670_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n710_), .A2(new_n319_), .A3(new_n615_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n413_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n737_), .B1(new_n743_), .B2(new_n736_), .ZN(G1336gat));
  INV_X1    g543(.A(G92gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n735_), .A2(new_n745_), .A3(new_n638_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n741_), .A2(new_n638_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n748_), .B2(new_n745_), .ZN(G1337gat));
  OAI21_X1  g548(.A(G99gat), .B1(new_n740_), .B2(new_n364_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n735_), .A2(new_n214_), .A3(new_n216_), .A4(new_n541_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n735_), .A2(new_n215_), .A3(new_n705_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n705_), .B(new_n739_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(G106gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G106gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n754_), .B(new_n760_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1339gat));
  NAND2_X1  g563(.A1(new_n617_), .A2(new_n614_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n601_), .A2(new_n604_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n604_), .B1(new_n597_), .B2(new_n246_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n610_), .B1(new_n603_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n613_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n591_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n572_), .A2(new_n580_), .A3(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n576_), .A2(new_n578_), .A3(KEYINPUT55), .A4(new_n570_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n776_), .B(new_n571_), .C1(new_n575_), .C2(new_n577_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n588_), .B1(new_n774_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n572_), .A2(new_n580_), .A3(new_n773_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n571_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT116), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n777_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n784_), .A2(new_n787_), .A3(new_n775_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(KEYINPUT56), .A3(new_n588_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n772_), .B1(new_n783_), .B2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n766_), .B(new_n274_), .C1(new_n790_), .C2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(KEYINPUT58), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n772_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n788_), .A2(KEYINPUT56), .A3(new_n588_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n588_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n791_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n766_), .B1(new_n800_), .B2(new_n274_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n795_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n615_), .A2(new_n591_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n783_), .B2(new_n789_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n592_), .A2(new_n771_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n269_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT57), .B(new_n269_), .C1(new_n804_), .C2(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n662_), .B1(new_n802_), .B2(new_n811_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n711_), .A2(KEYINPUT115), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n711_), .A2(KEYINPUT115), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n710_), .A2(new_n275_), .A3(new_n813_), .A4(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT54), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n812_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n705_), .A2(new_n638_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n621_), .A2(new_n364_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n817_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n815_), .B(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n795_), .B2(new_n801_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n274_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT118), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(KEYINPUT119), .A3(new_n794_), .A4(new_n793_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n591_), .B(new_n615_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n805_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT57), .B1(new_n832_), .B2(new_n269_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n810_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n827_), .A2(new_n830_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n825_), .B1(new_n836_), .B2(new_n662_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n820_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n765_), .B(new_n823_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G113gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n836_), .A2(new_n662_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n816_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n821_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n630_), .A2(G113gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(G1340gat));
  OAI21_X1  g645(.A(new_n823_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n847_));
  OAI21_X1  g646(.A(G120gat), .B1(new_n847_), .B2(new_n710_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n849_));
  AOI21_X1  g648(.A(G120gat), .B1(new_n596_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT121), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n849_), .B2(G120gat), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n838_), .B(new_n851_), .C1(new_n850_), .C2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n848_), .A2(new_n854_), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n847_), .B2(new_n662_), .ZN(new_n856_));
  OR3_X1    g655(.A1(new_n844_), .A2(G127gat), .A3(new_n662_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1342gat));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n859_), .B(new_n860_), .C1(new_n844_), .C2(new_n269_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n837_), .A2(new_n269_), .A3(new_n820_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT122), .B1(new_n862_), .B2(G134gat), .ZN(new_n863_));
  INV_X1    g662(.A(new_n823_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n844_), .B2(KEYINPUT59), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n275_), .A2(new_n860_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n861_), .A2(new_n863_), .B1(new_n865_), .B2(new_n866_), .ZN(G1343gat));
  NAND3_X1  g666(.A1(new_n705_), .A2(new_n413_), .A3(new_n364_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n638_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n842_), .B2(new_n816_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n615_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n596_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n871_), .B2(new_n319_), .ZN(new_n877_));
  NOR4_X1   g676(.A1(new_n837_), .A2(KEYINPUT123), .A3(new_n662_), .A4(new_n870_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n877_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n829_), .A2(new_n794_), .A3(new_n793_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n811_), .B1(new_n882_), .B2(new_n826_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n319_), .B1(new_n883_), .B2(new_n830_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n319_), .B(new_n869_), .C1(new_n884_), .C2(new_n825_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT123), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n871_), .A2(new_n876_), .A3(new_n319_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n879_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n881_), .A2(new_n888_), .ZN(G1346gat));
  INV_X1    g688(.A(new_n871_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G162gat), .B1(new_n890_), .B2(new_n275_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n871_), .A2(new_n380_), .A3(new_n633_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1347gat));
  NAND2_X1  g692(.A1(new_n638_), .A2(new_n414_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT124), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n705_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n817_), .A2(new_n615_), .A3(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT62), .B1(new_n897_), .B2(KEYINPUT22), .ZN(new_n898_));
  OAI21_X1  g697(.A(G169gat), .B1(new_n897_), .B2(KEYINPUT62), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n324_), .B2(new_n898_), .ZN(G1348gat));
  AND2_X1   g700(.A1(new_n817_), .A2(new_n896_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G176gat), .B1(new_n902_), .B2(new_n596_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n837_), .A2(new_n705_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n895_), .A2(new_n325_), .A3(new_n710_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  NOR2_X1   g705(.A1(new_n895_), .A2(new_n662_), .ZN(new_n907_));
  AOI21_X1  g706(.A(G183gat), .B1(new_n904_), .B2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n662_), .A2(new_n333_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n902_), .B2(new_n909_), .ZN(G1350gat));
  NAND2_X1  g709(.A1(new_n902_), .A2(new_n274_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(G190gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n902_), .A2(new_n633_), .A3(new_n332_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1351gat));
  AND3_X1   g713(.A1(new_n638_), .A2(new_n539_), .A3(new_n364_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n843_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n630_), .ZN(new_n917_));
  INV_X1    g716(.A(G197gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1352gat));
  NOR2_X1   g718(.A1(new_n916_), .A2(new_n710_), .ZN(new_n920_));
  INV_X1    g719(.A(G204gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1353gat));
  INV_X1    g721(.A(new_n916_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n662_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n924_));
  OR3_X1    g723(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  OAI21_X1  g725(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n923_), .A2(new_n924_), .B1(new_n927_), .B2(new_n925_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1354gat));
  INV_X1    g728(.A(G218gat), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n916_), .A2(new_n930_), .A3(new_n275_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n843_), .A2(new_n633_), .A3(new_n915_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933_));
  AOI21_X1  g732(.A(G218gat), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT126), .B1(new_n916_), .B2(new_n269_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n931_), .B1(new_n934_), .B2(new_n935_), .ZN(G1355gat));
endmodule


