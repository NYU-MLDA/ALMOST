//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT71), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G230gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT64), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT7), .Z(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n209_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT68), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n217_), .B(new_n209_), .C1(new_n211_), .C2(new_n214_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(KEYINPUT8), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n212_), .B(KEYINPUT6), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT67), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n220_), .B(new_n209_), .C1(new_n222_), .C2(new_n211_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n214_), .B(KEYINPUT67), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT10), .B(G99gat), .Z(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n206_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT66), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(G85gat), .B2(G92gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n229_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n224_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G57gat), .B(G64gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n240_), .A2(KEYINPUT69), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(KEYINPUT69), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n241_), .A2(new_n242_), .A3(KEYINPUT11), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT11), .B1(new_n241_), .B2(new_n242_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G71gat), .B(G78gat), .Z(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n239_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n237_), .B1(new_n219_), .B2(new_n223_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n248_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n205_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G120gat), .B(G148gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT5), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G176gat), .B(G204gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT12), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(new_n251_), .B2(new_n248_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n224_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n219_), .A2(KEYINPUT70), .A3(new_n223_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n237_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n248_), .A2(new_n260_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n261_), .B(new_n252_), .C1(new_n265_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n205_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n254_), .B(new_n259_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n264_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT70), .B1(new_n219_), .B2(new_n223_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n238_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n266_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n275_), .A2(new_n205_), .A3(new_n252_), .A4(new_n261_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n259_), .B1(new_n276_), .B2(new_n254_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n203_), .B1(new_n271_), .B2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n265_), .A2(new_n267_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n261_), .A2(new_n252_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n269_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n258_), .B1(new_n281_), .B2(new_n253_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(KEYINPUT71), .A3(new_n270_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT13), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n278_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n278_), .A2(new_n283_), .A3(KEYINPUT72), .A4(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n278_), .A2(new_n283_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(KEYINPUT13), .ZN(new_n292_));
  AOI211_X1 g091(.A(KEYINPUT73), .B(new_n284_), .C1(new_n278_), .C2(new_n283_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n289_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G229gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296_));
  INV_X1    g095(.A(G8gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  XOR2_X1   g100(.A(G29gat), .B(G36gat), .Z(new_n302_));
  XOR2_X1   g101(.A(G43gat), .B(G50gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n302_), .B(new_n303_), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n299_), .B(new_n300_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n295_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT81), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT76), .B(KEYINPUT15), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n304_), .B(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n312_), .A2(new_n301_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n305_), .A3(new_n295_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G113gat), .B(G141gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G169gat), .B(G197gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n314_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(KEYINPUT82), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n319_), .A2(new_n323_), .A3(new_n320_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G231gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n307_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(new_n248_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G127gat), .B(G155gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G183gat), .B(G211gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT17), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n329_), .A2(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n334_), .A2(KEYINPUT17), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n329_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n326_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n338_), .A2(new_n326_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n294_), .A2(new_n325_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT104), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT23), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(G183gat), .A3(G190gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G183gat), .ZN(new_n352_));
  INV_X1    g151(.A(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n348_), .A2(KEYINPUT87), .A3(G183gat), .A4(G190gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(KEYINPUT86), .A2(G176gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(KEYINPUT86), .A2(G176gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G169gat), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n357_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT24), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n347_), .A2(new_n349_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(KEYINPUT84), .A2(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT26), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT26), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n352_), .A2(KEYINPUT25), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(G183gat), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .A4(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT85), .B1(new_n375_), .B2(new_n357_), .ZN(new_n376_));
  INV_X1    g175(.A(G169gat), .ZN(new_n377_));
  INV_X1    g176(.A(G176gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT85), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT24), .A4(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n366_), .A2(new_n374_), .A3(new_n376_), .A4(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n363_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(G71gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G99gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n384_), .B(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G127gat), .B(G134gat), .Z(new_n390_));
  XOR2_X1   g189(.A(G113gat), .B(G120gat), .Z(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  XNOR2_X1  g191(.A(new_n389_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G15gat), .B(G43gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT88), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT30), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT31), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n397_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G22gat), .B(G50gat), .Z(new_n402_));
  NAND2_X1  g201(.A1(G141gat), .A2(G148gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT2), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G141gat), .A2(G148gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT3), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n404_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(G155gat), .A2(G162gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(G155gat), .A2(G162gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT1), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n412_), .B1(new_n411_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT89), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n411_), .B2(new_n415_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n406_), .A2(new_n403_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n414_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT28), .B1(new_n424_), .B2(KEYINPUT29), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT90), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n410_), .A2(new_n413_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT28), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n425_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n426_), .B1(new_n425_), .B2(new_n430_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n402_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n402_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n431_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(G197gat), .A2(G204gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G197gat), .A2(G204gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT21), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(KEYINPUT21), .A3(new_n440_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G211gat), .B(G218gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n444_), .A2(new_n445_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G228gat), .ZN(new_n449_));
  INV_X1    g248(.A(G233gat), .ZN(new_n450_));
  OAI221_X1 g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .C1(new_n427_), .C2(new_n429_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n448_), .B1(new_n427_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n449_), .A2(new_n450_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT92), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT92), .B1(new_n454_), .B2(new_n455_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n451_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G78gat), .B(G106gat), .Z(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n460_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n454_), .A2(new_n455_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT92), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n456_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n462_), .B1(new_n466_), .B2(new_n451_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n438_), .B1(new_n461_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n459_), .A2(new_n460_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n462_), .A3(new_n451_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n434_), .A4(new_n437_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G1gat), .B(G29gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G85gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT0), .B(G57gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  NAND2_X1  g275(.A1(new_n424_), .A2(new_n392_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n390_), .B(new_n391_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n427_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G225gat), .A2(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n477_), .A2(KEYINPUT4), .A3(new_n479_), .ZN(new_n485_));
  OR3_X1    g284(.A1(new_n427_), .A2(KEYINPUT4), .A3(new_n478_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n482_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n476_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n489_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n485_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT99), .Z(new_n493_));
  INV_X1    g292(.A(new_n476_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n494_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n490_), .B(new_n491_), .C1(new_n493_), .C2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G8gat), .B(G36gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G64gat), .B(G92gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n502_));
  AND2_X1   g301(.A1(G226gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n351_), .A2(new_n355_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n353_), .A2(KEYINPUT26), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n369_), .A2(G190gat), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n371_), .A2(new_n373_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n375_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n512_), .B2(new_n381_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .A4(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n510_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n351_), .A2(new_n355_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT95), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT96), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n347_), .A2(new_n349_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n354_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n362_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(new_n362_), .B2(new_n520_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n514_), .B(new_n517_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n448_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT97), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(KEYINPUT97), .A3(new_n448_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n363_), .A2(new_n446_), .A3(new_n383_), .A4(new_n447_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT20), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT94), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n505_), .B1(new_n528_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n522_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n362_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n448_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(new_n517_), .A4(new_n514_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n505_), .A2(KEYINPUT20), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n448_), .B2(new_n384_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n501_), .B1(new_n535_), .B2(new_n543_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n523_), .A2(KEYINPUT97), .A3(new_n448_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT97), .B1(new_n523_), .B2(new_n448_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n534_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n504_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n501_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n543_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n544_), .A2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n496_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n362_), .A2(new_n520_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n515_), .A2(new_n516_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT20), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT100), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n384_), .A2(new_n448_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(KEYINPUT100), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n504_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(new_n547_), .B2(new_n504_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(KEYINPUT32), .A3(new_n549_), .ZN(new_n564_));
  OR3_X1    g363(.A1(new_n484_), .A2(new_n487_), .A3(new_n476_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n488_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n543_), .B1(new_n547_), .B2(new_n504_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n549_), .A2(KEYINPUT32), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n472_), .B1(new_n553_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT27), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n563_), .A2(new_n501_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n567_), .B2(new_n549_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n552_), .A2(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n566_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n472_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n401_), .B1(new_n572_), .B2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n400_), .A2(new_n566_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT101), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n576_), .B2(new_n472_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n549_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n584_));
  AOI211_X1 g383(.A(new_n501_), .B(new_n543_), .C1(new_n547_), .C2(new_n504_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n573_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n574_), .A2(new_n551_), .A3(KEYINPUT27), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n586_), .A2(new_n472_), .A3(new_n587_), .A4(new_n582_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n581_), .B1(new_n583_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT102), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n472_), .A3(new_n587_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT101), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n588_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT102), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(new_n581_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n580_), .B1(new_n591_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT35), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n251_), .A2(new_n304_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n265_), .B2(new_n312_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n601_), .A2(new_n598_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  OAI221_X1 g404(.A(new_n602_), .B1(new_n598_), .B2(new_n601_), .C1(new_n265_), .C2(new_n312_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT36), .ZN(new_n608_));
  XOR2_X1   g407(.A(G190gat), .B(G218gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT77), .ZN(new_n610_));
  XOR2_X1   g409(.A(G134gat), .B(G162gat), .Z(new_n611_));
  XOR2_X1   g410(.A(new_n610_), .B(new_n611_), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(KEYINPUT78), .ZN(new_n614_));
  INV_X1    g413(.A(new_n612_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT36), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n616_), .B1(new_n619_), .B2(new_n615_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n614_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n597_), .A2(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n294_), .A2(KEYINPUT104), .A3(new_n325_), .A4(new_n342_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n345_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n202_), .B1(new_n627_), .B2(new_n566_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT105), .Z(new_n629_));
  NOR3_X1   g428(.A1(new_n271_), .A2(new_n277_), .A3(new_n203_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT71), .B1(new_n282_), .B2(new_n270_), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT13), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT73), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n291_), .A2(new_n290_), .A3(KEYINPUT13), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n633_), .A2(new_n634_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT74), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n572_), .A2(new_n579_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n400_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n595_), .B1(new_n594_), .B2(new_n581_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n581_), .ZN(new_n640_));
  AOI211_X1 g439(.A(KEYINPUT102), .B(new_n640_), .C1(new_n593_), .C2(new_n588_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n638_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n325_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT83), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n322_), .A2(KEYINPUT83), .A3(new_n324_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n642_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n614_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n620_), .A2(new_n621_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n648_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n617_), .A2(KEYINPUT37), .A3(new_n622_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AND4_X1   g453(.A1(new_n342_), .A2(new_n636_), .A3(new_n647_), .A4(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n657_));
  AOI21_X1  g456(.A(G1gat), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n566_), .A3(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n656_), .A2(new_n657_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n629_), .A2(new_n661_), .ZN(G1324gat));
  NAND2_X1  g461(.A1(new_n586_), .A2(new_n587_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n345_), .A2(new_n663_), .A3(new_n625_), .A4(new_n626_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n664_), .A2(KEYINPUT106), .A3(G8gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT106), .B1(new_n664_), .B2(G8gat), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n667_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n655_), .A2(new_n297_), .A3(new_n663_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n668_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1325gat));
  INV_X1    g474(.A(G15gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n627_), .B2(new_n401_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT41), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n655_), .A2(new_n676_), .A3(new_n401_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1326gat));
  INV_X1    g479(.A(G22gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n627_), .B2(new_n578_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT42), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n655_), .A2(new_n681_), .A3(new_n578_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1327gat));
  INV_X1    g484(.A(G29gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n294_), .A2(new_n325_), .A3(new_n341_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n597_), .B2(new_n654_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n642_), .A2(new_n689_), .A3(new_n653_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n687_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT108), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n635_), .A2(new_n643_), .A3(new_n342_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n642_), .A2(new_n689_), .A3(new_n653_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n689_), .B1(new_n642_), .B2(new_n653_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698_));
  INV_X1    g497(.A(new_n692_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n693_), .A2(new_n700_), .B1(KEYINPUT44), .B2(new_n691_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n686_), .B1(new_n701_), .B2(new_n566_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n623_), .A2(new_n342_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n635_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n647_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n566_), .A2(new_n686_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT109), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OR3_X1    g509(.A1(new_n702_), .A2(KEYINPUT110), .A3(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT110), .B1(new_n702_), .B2(new_n710_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n706_), .A2(new_n714_), .A3(new_n663_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT45), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n576_), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n691_), .A2(KEYINPUT108), .A3(new_n692_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n698_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT111), .B(new_n717_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G36gat), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n693_), .A2(new_n700_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT111), .B1(new_n722_), .B2(new_n717_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n716_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(KEYINPUT46), .B(new_n716_), .C1(new_n721_), .C2(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1329gat));
  NAND2_X1  g527(.A1(new_n691_), .A2(KEYINPUT44), .ZN(new_n729_));
  INV_X1    g528(.A(G43gat), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n400_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n729_), .B(new_n731_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT112), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n701_), .A2(new_n734_), .A3(new_n731_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n706_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n730_), .B1(new_n736_), .B2(new_n400_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n733_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT47), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n733_), .A2(new_n735_), .A3(new_n740_), .A4(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1330gat));
  AOI21_X1  g541(.A(G50gat), .B1(new_n706_), .B2(new_n578_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n578_), .A2(G50gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n701_), .B2(new_n744_), .ZN(G1331gat));
  NAND2_X1  g544(.A1(new_n642_), .A2(new_n643_), .ZN(new_n746_));
  NOR4_X1   g545(.A1(new_n746_), .A2(new_n294_), .A3(new_n341_), .A4(new_n653_), .ZN(new_n747_));
  INV_X1    g546(.A(G57gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n566_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n636_), .A2(new_n341_), .A3(new_n646_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n625_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(new_n566_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n752_), .B2(new_n748_), .ZN(G1332gat));
  INV_X1    g552(.A(G64gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n747_), .A2(new_n754_), .A3(new_n663_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n751_), .A2(new_n663_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(G64gat), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(KEYINPUT48), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(KEYINPUT48), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1333gat));
  NAND3_X1  g559(.A1(new_n747_), .A2(new_n386_), .A3(new_n401_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n751_), .A2(new_n401_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G71gat), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n763_), .A2(KEYINPUT49), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(KEYINPUT49), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(G1334gat));
  INV_X1    g565(.A(G78gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n747_), .A2(new_n767_), .A3(new_n578_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n751_), .A2(new_n578_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G78gat), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(KEYINPUT50), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(KEYINPUT50), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(G1335gat));
  NAND2_X1  g572(.A1(new_n688_), .A2(new_n690_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n294_), .A2(new_n325_), .A3(new_n342_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n577_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n636_), .A2(new_n704_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n746_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(KEYINPUT113), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT113), .B1(new_n778_), .B2(new_n779_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n577_), .A2(G85gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n777_), .B1(new_n782_), .B2(new_n783_), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n776_), .B2(new_n576_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n576_), .A2(G92gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n782_), .B2(new_n786_), .ZN(G1337gat));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n226_), .B(new_n401_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G99gat), .B1(new_n776_), .B2(new_n400_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n788_), .B(KEYINPUT51), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT114), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(KEYINPUT51), .ZN(new_n794_));
  AND4_X1   g593(.A1(new_n793_), .A2(new_n789_), .A3(new_n790_), .A4(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n791_), .A2(new_n795_), .ZN(G1338gat));
  NOR2_X1   g595(.A1(new_n472_), .A2(G106gat), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n774_), .A2(new_n578_), .A3(new_n775_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G106gat), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(KEYINPUT52), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(KEYINPUT52), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n782_), .A2(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g603(.A1(new_n594_), .A2(new_n566_), .A3(new_n401_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n806_));
  INV_X1    g605(.A(new_n268_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT55), .A3(new_n205_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n276_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n268_), .A2(new_n269_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n258_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n258_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n305_), .A2(new_n308_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n317_), .B1(new_n818_), .B2(new_n295_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n819_), .A2(KEYINPUT118), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(KEYINPUT118), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n313_), .A2(G229gat), .A3(G233gat), .A4(new_n305_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n318_), .ZN(new_n824_));
  XOR2_X1   g623(.A(new_n824_), .B(KEYINPUT119), .Z(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n270_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n817_), .A2(KEYINPUT58), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n653_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT58), .B1(new_n817_), .B2(new_n827_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n806_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n830_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n832_), .A2(KEYINPUT121), .A3(new_n653_), .A4(new_n828_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n325_), .A2(new_n270_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n291_), .A2(new_n825_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n623_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n837_), .A2(new_n838_), .A3(KEYINPUT57), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT57), .B1(new_n837_), .B2(new_n838_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n831_), .B(new_n833_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n341_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n843_));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n341_), .B(new_n845_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n294_), .A2(new_n654_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n844_), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT117), .Z(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n294_), .A2(new_n654_), .A3(new_n849_), .A4(new_n846_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n805_), .B1(new_n842_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G113gat), .B1(new_n854_), .B2(new_n325_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n855_), .A2(KEYINPUT122), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(KEYINPUT122), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n841_), .A2(new_n341_), .B1(new_n852_), .B2(new_n851_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT59), .B1(new_n858_), .B2(new_n805_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n805_), .A2(KEYINPUT59), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n837_), .A2(new_n838_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n837_), .A2(new_n838_), .A3(KEYINPUT57), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n832_), .A2(new_n653_), .A3(new_n828_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n342_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n853_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n860_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n859_), .A2(new_n869_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n646_), .A2(G113gat), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n856_), .A2(new_n857_), .B1(new_n870_), .B2(new_n871_), .ZN(G1340gat));
  XNOR2_X1  g671(.A(new_n294_), .B(KEYINPUT74), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n859_), .A2(new_n873_), .A3(new_n869_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n859_), .A2(new_n876_), .A3(new_n873_), .A4(new_n869_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(G120gat), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(G120gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n294_), .B2(KEYINPUT60), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n854_), .B(new_n880_), .C1(KEYINPUT60), .C2(new_n879_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(G1341gat));
  NAND2_X1  g681(.A1(new_n870_), .A2(new_n342_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G127gat), .ZN(new_n884_));
  INV_X1    g683(.A(new_n854_), .ZN(new_n885_));
  OR3_X1    g684(.A1(new_n885_), .A2(G127gat), .A3(new_n341_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1342gat));
  NAND2_X1  g686(.A1(new_n870_), .A2(new_n653_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G134gat), .ZN(new_n889_));
  OR3_X1    g688(.A1(new_n885_), .A2(G134gat), .A3(new_n623_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1343gat));
  NOR3_X1   g690(.A1(new_n663_), .A2(new_n577_), .A3(new_n472_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n858_), .A2(new_n401_), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n325_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n873_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g697(.A1(new_n842_), .A2(new_n853_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n899_), .A2(new_n342_), .A3(new_n400_), .A4(new_n892_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT124), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n858_), .A2(new_n401_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(new_n342_), .A4(new_n892_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n901_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1346gat));
  INV_X1    g707(.A(G162gat), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n902_), .A2(new_n909_), .A3(new_n624_), .A4(new_n892_), .ZN(new_n910_));
  NOR4_X1   g709(.A1(new_n858_), .A2(new_n401_), .A3(new_n654_), .A4(new_n893_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n909_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT125), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n910_), .B(new_n914_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1347gat));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n640_), .A2(new_n576_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n578_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n643_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n917_), .B1(new_n922_), .B2(new_n377_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n361_), .ZN(new_n924_));
  OAI211_X1 g723(.A(KEYINPUT62), .B(G169gat), .C1(new_n921_), .C2(new_n643_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(G1348gat));
  INV_X1    g725(.A(new_n921_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n635_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n858_), .A2(new_n578_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n636_), .A2(new_n378_), .A3(new_n919_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n928_), .A2(new_n360_), .B1(new_n929_), .B2(new_n930_), .ZN(G1349gat));
  AOI211_X1 g730(.A(new_n341_), .B(new_n921_), .C1(new_n371_), .C2(new_n373_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n929_), .A2(new_n342_), .A3(new_n918_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n352_), .B2(new_n933_), .ZN(G1350gat));
  AND3_X1   g733(.A1(new_n624_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n927_), .A2(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(G190gat), .B1(new_n921_), .B2(new_n654_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n936_), .A2(KEYINPUT126), .A3(new_n937_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1351gat));
  NOR3_X1   g741(.A1(new_n576_), .A2(new_n566_), .A3(new_n472_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n902_), .A2(new_n325_), .A3(new_n943_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g744(.A1(new_n902_), .A2(new_n943_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n636_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n947_), .B(new_n948_), .ZN(G1353gat));
  INV_X1    g748(.A(new_n946_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  AND2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n950_), .B(new_n342_), .C1(new_n951_), .C2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n946_), .A2(new_n341_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n954_), .B2(new_n951_), .ZN(G1354gat));
  OR3_X1    g754(.A1(new_n946_), .A2(G218gat), .A3(new_n623_), .ZN(new_n956_));
  OAI21_X1  g755(.A(G218gat), .B1(new_n946_), .B2(new_n654_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1355gat));
endmodule


