//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT74), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208_));
  INV_X1    g007(.A(G1gat), .ZN(new_n209_));
  INV_X1    g008(.A(G8gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G1gat), .B(G8gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G29gat), .B(G36gat), .Z(new_n215_));
  INV_X1    g014(.A(G43gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G29gat), .B(G36gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G43gat), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n217_), .A2(G50gat), .A3(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(G50gat), .B1(new_n217_), .B2(new_n219_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT15), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G50gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n219_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n218_), .A2(G43gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n217_), .A2(G50gat), .A3(new_n219_), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT15), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n214_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n214_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(new_n228_), .A3(new_n227_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n230_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n227_), .A2(new_n228_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n214_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n231_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n207_), .B1(new_n234_), .B2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n231_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT74), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n206_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n206_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n235_), .A2(new_n214_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n222_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n227_), .A2(KEYINPUT15), .A3(new_n228_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n246_), .B1(new_n249_), .B2(new_n214_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n241_), .B1(new_n250_), .B2(new_n231_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n244_), .B(new_n245_), .C1(new_n251_), .C2(new_n207_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n243_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G230gat), .A2(G233gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT10), .B(G99gat), .Z(new_n256_));
  INV_X1    g055(.A(G106gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G85gat), .B(G92gat), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT9), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT9), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(G85gat), .A3(G92gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G99gat), .A2(G106gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT6), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n258_), .A2(new_n260_), .A3(new_n262_), .A4(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n266_));
  OR3_X1    g065(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT8), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n259_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n268_), .B2(new_n259_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n265_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT64), .B(G71gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G78gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(G57gat), .B(G64gat), .Z(new_n275_));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n276_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n274_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(G78gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n273_), .B(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n275_), .A2(new_n276_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n255_), .B1(new_n272_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT12), .B1(new_n272_), .B2(new_n284_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n272_), .A2(new_n284_), .A3(KEYINPUT12), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n279_), .A2(new_n283_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n291_), .B(new_n265_), .C1(new_n271_), .C2(new_n270_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(KEYINPUT66), .A3(new_n255_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n287_), .A2(new_n289_), .A3(new_n290_), .A4(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n272_), .A2(new_n284_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n292_), .A3(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n272_), .A2(new_n284_), .A3(KEYINPUT65), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n297_), .A2(G230gat), .A3(G233gat), .A4(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G120gat), .B(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(G204gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT5), .ZN(new_n303_));
  INV_X1    g102(.A(G176gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n294_), .A2(new_n299_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n305_), .B1(new_n294_), .B2(new_n299_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT13), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(KEYINPUT67), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(KEYINPUT67), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n310_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n309_), .B1(KEYINPUT67), .B2(new_n311_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G127gat), .B(G134gat), .Z(new_n317_));
  OR2_X1    g116(.A1(G113gat), .A2(G120gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G113gat), .A2(G120gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT78), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT78), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n322_), .A3(new_n319_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n317_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT79), .ZN(new_n325_));
  INV_X1    g124(.A(new_n324_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n321_), .A2(new_n323_), .A3(new_n317_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n325_), .B1(new_n328_), .B2(KEYINPUT79), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT80), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G155gat), .A3(G162gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT81), .B1(new_n334_), .B2(KEYINPUT1), .ZN(new_n335_));
  OR2_X1    g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(KEYINPUT1), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n331_), .A2(new_n333_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .A4(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n334_), .A2(KEYINPUT83), .A3(new_n336_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT83), .B1(new_n334_), .B2(new_n336_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n342_), .B1(KEYINPUT82), .B2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT82), .B(KEYINPUT3), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(new_n342_), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n344_), .B(KEYINPUT2), .Z(new_n352_));
  OAI22_X1  g151(.A1(new_n346_), .A2(new_n347_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n345_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n329_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n327_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT99), .B1(new_n357_), .B2(new_n324_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT99), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n326_), .A2(new_n359_), .A3(new_n327_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n358_), .A2(new_n360_), .A3(new_n345_), .A4(new_n353_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n355_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT100), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT100), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n355_), .A2(new_n364_), .A3(new_n356_), .A4(new_n361_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n356_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n355_), .B2(new_n361_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT4), .B1(new_n329_), .B2(new_n354_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n367_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT0), .B(G57gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G85gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(G1gat), .B(G29gat), .Z(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n371_), .A2(new_n378_), .A3(new_n363_), .A4(new_n365_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT19), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n205_), .A2(G204gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT85), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(G197gat), .B2(new_n301_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n205_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n384_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G211gat), .B(G218gat), .Z(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT21), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT88), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n388_), .A2(KEYINPUT88), .A3(KEYINPUT21), .A4(new_n389_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT21), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n395_), .B(new_n384_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n301_), .A2(G197gat), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n395_), .B1(new_n399_), .B2(new_n384_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(new_n389_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT85), .B1(new_n205_), .B2(G204gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n385_), .A2(new_n301_), .A3(G197gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n404_), .A2(KEYINPUT86), .A3(new_n395_), .A4(new_n384_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n398_), .A2(new_n401_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT87), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT87), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n398_), .A2(new_n405_), .A3(new_n408_), .A4(new_n401_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n394_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G183gat), .A2(G190gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT23), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(G183gat), .B2(G190gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n203_), .A2(new_n304_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT22), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(KEYINPUT75), .B2(G169gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(KEYINPUT75), .A2(G169gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n304_), .B1(new_n418_), .B2(KEYINPUT22), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n413_), .B(new_n415_), .C1(new_n417_), .C2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G169gat), .A2(G176gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n415_), .A2(KEYINPUT24), .A3(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n422_), .A2(KEYINPUT24), .ZN(new_n424_));
  OR2_X1    g223(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G190gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n423_), .A2(new_n424_), .A3(new_n429_), .A4(new_n412_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n420_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT20), .B(new_n383_), .C1(new_n410_), .C2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n416_), .A2(G169gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n203_), .A2(KEYINPUT22), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n304_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT95), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n414_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n414_), .A2(new_n438_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT96), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT96), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT22), .B(G169gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT95), .B1(new_n444_), .B2(new_n304_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n443_), .B(new_n440_), .C1(new_n445_), .C2(new_n414_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(new_n446_), .A3(new_n413_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n424_), .A2(new_n412_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT94), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n427_), .A2(KEYINPUT93), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT93), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n428_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n424_), .A2(KEYINPUT94), .A3(new_n412_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n450_), .A2(new_n454_), .A3(new_n423_), .A4(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n447_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT97), .B1(new_n410_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n410_), .A2(new_n457_), .A3(KEYINPUT97), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n434_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n407_), .A2(new_n409_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n394_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n447_), .A2(new_n456_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n410_), .B2(new_n432_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n382_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n461_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT18), .B(G64gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(G92gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G8gat), .B(G36gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(new_n474_), .Z(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT98), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n461_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT27), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n471_), .A2(KEYINPUT98), .A3(new_n476_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT101), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n464_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n410_), .A2(KEYINPUT89), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n465_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n484_), .B1(new_n488_), .B2(new_n467_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n464_), .A2(new_n431_), .ZN(new_n490_));
  AOI211_X1 g289(.A(new_n485_), .B(new_n394_), .C1(new_n407_), .C2(new_n409_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT89), .B1(new_n462_), .B2(new_n463_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n457_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n489_), .A2(new_n490_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n382_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n469_), .A2(new_n382_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n475_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT102), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n410_), .A2(new_n457_), .A3(KEYINPUT97), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(new_n458_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n502_), .A2(new_n434_), .B1(new_n469_), .B2(new_n382_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n500_), .B1(new_n503_), .B2(new_n475_), .ZN(new_n504_));
  AND4_X1   g303(.A1(new_n500_), .A2(new_n461_), .A3(new_n470_), .A4(new_n475_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT27), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n380_), .B(new_n483_), .C1(new_n499_), .C2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G78gat), .B(G106gat), .Z(new_n508_));
  AND2_X1   g307(.A1(new_n354_), .A2(KEYINPUT29), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT84), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(G233gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n510_), .A2(G233gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(G228gat), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n509_), .A2(new_n410_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n354_), .A2(KEYINPUT29), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n486_), .A2(new_n487_), .A3(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n519_), .A2(KEYINPUT90), .A3(new_n515_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT90), .B1(new_n519_), .B2(new_n515_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n508_), .B(new_n517_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n354_), .A2(KEYINPUT29), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G22gat), .B(G50gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT28), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n523_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n527_), .A2(KEYINPUT91), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n491_), .A2(new_n492_), .A3(new_n509_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n530_), .B1(new_n531_), .B2(new_n514_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n519_), .A2(KEYINPUT90), .A3(new_n515_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n508_), .B1(new_n534_), .B2(new_n517_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n508_), .ZN(new_n536_));
  AOI211_X1 g335(.A(new_n536_), .B(new_n516_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n529_), .B1(new_n538_), .B2(new_n528_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n516_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT92), .B1(new_n540_), .B2(new_n508_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n517_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n536_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n527_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n507_), .A2(new_n539_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n475_), .A2(KEYINPUT32), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n377_), .A2(new_n379_), .B1(new_n503_), .B2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n497_), .B1(new_n495_), .B2(new_n382_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(new_n548_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n480_), .A2(new_n482_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n356_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n355_), .A2(new_n367_), .A3(new_n361_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n376_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT33), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n379_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n366_), .A2(KEYINPUT33), .A3(new_n378_), .A4(new_n371_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n552_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n542_), .A2(new_n536_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(new_n528_), .A3(new_n522_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n522_), .A2(new_n528_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n526_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n551_), .B(new_n561_), .C1(new_n565_), .C2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G227gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n329_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G15gat), .B(G43gat), .Z(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n569_), .A2(new_n570_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n572_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n569_), .A2(new_n570_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G71gat), .B(G99gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n431_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT76), .B(KEYINPUT30), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  AND3_X1   g380(.A1(new_n573_), .A2(new_n577_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n547_), .A2(new_n567_), .A3(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n546_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n479_), .A2(KEYINPUT102), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n503_), .A2(new_n500_), .A3(new_n475_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n481_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n550_), .B2(new_n475_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n591_), .A2(new_n483_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n587_), .A2(new_n592_), .A3(new_n380_), .A4(new_n584_), .ZN(new_n593_));
  AOI211_X1 g392(.A(new_n254_), .B(new_n316_), .C1(new_n586_), .C2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT68), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n249_), .A2(new_n595_), .A3(new_n272_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n249_), .B2(new_n272_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT34), .Z(new_n600_));
  INV_X1    g399(.A(KEYINPUT35), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n272_), .B2(new_n235_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n598_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(G134gat), .ZN(new_n607_));
  INV_X1    g406(.A(G162gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT36), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT71), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n604_), .A2(KEYINPUT69), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT69), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n614_), .B(new_n603_), .C1(new_n272_), .C2(new_n235_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n613_), .B(new_n615_), .C1(new_n597_), .C2(new_n596_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n616_), .A2(KEYINPUT70), .A3(new_n602_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT70), .B1(new_n616_), .B2(new_n602_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n605_), .B(new_n612_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT72), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n602_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT70), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n616_), .A2(KEYINPUT70), .A3(new_n602_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n626_), .A2(KEYINPUT72), .A3(new_n605_), .A4(new_n612_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n621_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n605_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n610_), .A2(KEYINPUT36), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n611_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT37), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n611_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n626_), .B2(new_n605_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n621_), .A2(new_n627_), .B1(new_n636_), .B2(new_n630_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT37), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n634_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n291_), .B(new_n232_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(G127gat), .B(G155gat), .Z(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(G183gat), .B(G211gat), .Z(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT17), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n642_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n649_), .B2(new_n642_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n639_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n594_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n380_), .B(KEYINPUT103), .Z(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n209_), .A3(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT38), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n637_), .A2(new_n653_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n594_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n380_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n662_), .ZN(G1324gat));
  OAI21_X1  g462(.A(G8gat), .B1(new_n661_), .B2(new_n592_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n592_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n656_), .A2(new_n210_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n661_), .B2(new_n585_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT41), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n655_), .A2(G15gat), .A3(new_n585_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1326gat));
  OAI21_X1  g473(.A(G22gat), .B1(new_n661_), .B2(new_n587_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT42), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n587_), .A2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n655_), .B2(new_n677_), .ZN(G1327gat));
  NAND2_X1  g477(.A1(new_n586_), .A2(new_n593_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n639_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT43), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n679_), .A2(new_n682_), .A3(new_n639_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n316_), .A2(new_n254_), .A3(new_n652_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n684_), .A2(new_n685_), .A3(KEYINPUT44), .A4(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n682_), .B1(new_n679_), .B2(new_n639_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n628_), .A2(KEYINPUT37), .A3(new_n631_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT37), .B1(new_n628_), .B2(new_n631_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT43), .B(new_n691_), .C1(new_n586_), .C2(new_n593_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT44), .B(new_n686_), .C1(new_n688_), .C2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT107), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n687_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n686_), .B1(new_n688_), .B2(new_n692_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n699_));
  OAI211_X1 g498(.A(KEYINPUT105), .B(new_n686_), .C1(new_n688_), .C2(new_n692_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n695_), .A2(new_n701_), .A3(new_n657_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G29gat), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n637_), .A2(new_n653_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT108), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n594_), .A2(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n706_), .A2(G29gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n380_), .B2(new_n707_), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n695_), .A2(new_n701_), .A3(new_n667_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G36gat), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n706_), .A2(G36gat), .A3(new_n592_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT45), .Z(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n710_), .A2(KEYINPUT46), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND3_X1  g516(.A1(new_n695_), .A2(new_n701_), .A3(new_n584_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G43gat), .ZN(new_n719_));
  INV_X1    g518(.A(new_n706_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n216_), .A3(new_n584_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(KEYINPUT47), .A3(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1330gat));
  NOR2_X1   g525(.A1(new_n565_), .A2(new_n566_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n720_), .A2(new_n224_), .A3(new_n727_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n695_), .A2(new_n701_), .A3(new_n727_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n224_), .ZN(G1331gat));
  INV_X1    g529(.A(new_n316_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(new_n253_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n679_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n654_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n657_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n734_), .A2(G57gat), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n380_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n733_), .A2(new_n737_), .A3(new_n660_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(G57gat), .B2(new_n738_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT109), .Z(G1332gat));
  NAND2_X1  g539(.A1(new_n733_), .A2(new_n660_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G64gat), .B1(new_n741_), .B2(new_n592_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT48), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n592_), .A2(G64gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n734_), .B2(new_n744_), .ZN(G1333gat));
  OAI21_X1  g544(.A(G71gat), .B1(new_n741_), .B2(new_n585_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT49), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n585_), .A2(G71gat), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT110), .Z(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n734_), .B2(new_n749_), .ZN(G1334gat));
  OAI21_X1  g549(.A(G78gat), .B1(new_n741_), .B2(new_n587_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT50), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n587_), .A2(G78gat), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT111), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n734_), .B2(new_n754_), .ZN(G1335gat));
  AND2_X1   g554(.A1(new_n733_), .A2(new_n705_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n657_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n732_), .A2(new_n653_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT112), .Z(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n737_), .A2(G85gat), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT113), .Z(new_n762_));
  AOI21_X1  g561(.A(new_n757_), .B1(new_n760_), .B2(new_n762_), .ZN(G1336gat));
  AOI21_X1  g562(.A(G92gat), .B1(new_n756_), .B2(new_n667_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT114), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n667_), .A2(G92gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n760_), .B2(new_n766_), .ZN(G1337gat));
  NAND2_X1  g566(.A1(new_n760_), .A2(new_n584_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G99gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n756_), .A2(new_n256_), .A3(new_n584_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n756_), .A2(new_n257_), .A3(new_n727_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n760_), .A2(new_n727_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(G106gat), .ZN(new_n776_));
  AOI211_X1 g575(.A(KEYINPUT52), .B(new_n257_), .C1(new_n760_), .C2(new_n727_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n773_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1339gat));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n250_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n232_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT116), .B1(new_n785_), .B2(new_n246_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n784_), .A2(new_n238_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n237_), .A2(new_n231_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n206_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n252_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n252_), .A3(KEYINPUT117), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n309_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n253_), .A2(KEYINPUT115), .A3(new_n306_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT115), .B1(new_n253_), .B2(new_n306_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n294_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n289_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(G230gat), .A3(G233gat), .ZN(new_n801_));
  INV_X1    g600(.A(new_n290_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n288_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n803_), .A2(KEYINPUT55), .A3(new_n287_), .A4(new_n293_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n801_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n305_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n794_), .B1(new_n797_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT57), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n812_), .A2(new_n637_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n814_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n253_), .A2(new_n306_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n253_), .A2(KEYINPUT115), .A3(new_n306_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n806_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n806_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n819_), .B(new_n820_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n794_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n816_), .B1(new_n825_), .B2(new_n632_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n815_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n821_), .A2(new_n828_), .B1(new_n793_), .B2(new_n792_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n809_), .A2(KEYINPUT119), .A3(new_n810_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n306_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n829_), .A2(new_n830_), .A3(KEYINPUT58), .A4(new_n306_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n833_), .B(new_n834_), .C1(new_n690_), .C2(new_n689_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n827_), .A2(new_n835_), .A3(KEYINPUT120), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT120), .B1(new_n827_), .B2(new_n835_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n652_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n691_), .A2(new_n254_), .A3(new_n652_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT54), .B1(new_n839_), .B2(new_n316_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n654_), .A2(new_n841_), .A3(new_n254_), .A4(new_n731_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT121), .B1(new_n838_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n833_), .A2(new_n834_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n691_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n814_), .B1(new_n812_), .B2(new_n637_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n825_), .A2(new_n632_), .A3(new_n816_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n845_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n827_), .A2(new_n835_), .A3(KEYINPUT120), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n653_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n840_), .A2(new_n842_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  NOR4_X1   g655(.A1(new_n735_), .A2(new_n667_), .A3(new_n727_), .A4(new_n585_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n844_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(G113gat), .B1(new_n859_), .B2(new_n253_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n653_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n855_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n857_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n858_), .B2(KEYINPUT59), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n865_), .A2(new_n253_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n860_), .B1(new_n866_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n731_), .B2(KEYINPUT60), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n859_), .B(new_n869_), .C1(KEYINPUT60), .C2(new_n868_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n865_), .A2(new_n316_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n868_), .ZN(G1341gat));
  AOI21_X1  g671(.A(G127gat), .B1(new_n859_), .B2(new_n652_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n865_), .A2(G127gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n652_), .ZN(G1342gat));
  AOI21_X1  g674(.A(G134gat), .B1(new_n859_), .B2(new_n637_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT122), .B(G134gat), .Z(new_n877_));
  NOR2_X1   g676(.A1(new_n691_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n865_), .B2(new_n878_), .ZN(G1343gat));
  AND3_X1   g678(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n854_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n587_), .A2(new_n584_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n592_), .A3(new_n657_), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(KEYINPUT123), .Z(new_n885_));
  NAND3_X1  g684(.A1(new_n882_), .A2(new_n253_), .A3(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g686(.A1(new_n882_), .A2(new_n316_), .A3(new_n885_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g688(.A1(new_n882_), .A2(new_n652_), .A3(new_n885_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  AND4_X1   g691(.A1(G162gat), .A2(new_n882_), .A3(new_n639_), .A4(new_n885_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n882_), .A2(new_n637_), .A3(new_n885_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n608_), .B2(new_n894_), .ZN(G1347gat));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n657_), .A2(new_n592_), .A3(new_n585_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n727_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n862_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n254_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n896_), .B1(new_n901_), .B2(new_n203_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n444_), .ZN(new_n903_));
  OAI211_X1 g702(.A(KEYINPUT62), .B(G169gat), .C1(new_n900_), .C2(new_n254_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n902_), .A2(KEYINPUT124), .A3(new_n903_), .A4(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1348gat));
  OAI21_X1  g708(.A(new_n304_), .B1(new_n900_), .B2(new_n731_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n898_), .A2(new_n304_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n844_), .A2(new_n587_), .A3(new_n856_), .A4(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n912_), .B2(new_n731_), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT125), .Z(G1349gat));
  NOR4_X1   g713(.A1(new_n900_), .A2(new_n453_), .A3(new_n451_), .A4(new_n653_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n882_), .A2(new_n587_), .A3(new_n652_), .A4(new_n897_), .ZN(new_n916_));
  INV_X1    g715(.A(G183gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n900_), .B2(new_n691_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n862_), .A2(new_n428_), .A3(new_n899_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n632_), .B2(new_n920_), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n592_), .A2(new_n737_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n844_), .A2(new_n856_), .A3(new_n883_), .A4(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n254_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n924_), .A2(KEYINPUT126), .A3(new_n205_), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT126), .B(G197gat), .Z(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n924_), .B2(new_n926_), .ZN(G1352gat));
  NOR2_X1   g726(.A1(new_n923_), .A2(new_n731_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(new_n301_), .ZN(G1353gat));
  NOR2_X1   g728(.A1(new_n923_), .A2(new_n653_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n930_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931_));
  XOR2_X1   g730(.A(KEYINPUT63), .B(G211gat), .Z(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n930_), .B2(new_n932_), .ZN(G1354gat));
  INV_X1    g732(.A(new_n922_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n880_), .A2(new_n881_), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(G218gat), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n935_), .A2(new_n936_), .A3(new_n637_), .A4(new_n883_), .ZN(new_n937_));
  OAI21_X1  g736(.A(G218gat), .B1(new_n923_), .B2(new_n691_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n937_), .A2(new_n938_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1355gat));
endmodule


