//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G71gat), .B(G78gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n202_), .B(KEYINPUT11), .Z(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(new_n206_), .B2(new_n204_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT9), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n208_), .A2(new_n209_), .A3(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n211_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT10), .B(G99gat), .Z(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n217_), .A2(new_n220_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n219_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n229_), .A2(new_n223_), .A3(new_n224_), .A4(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n214_), .A2(new_n208_), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n226_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n207_), .B(new_n236_), .Z(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT12), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n207_), .A2(new_n236_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n238_), .B1(KEYINPUT12), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G230gat), .A2(G233gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n241_), .B2(new_n237_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT5), .B(G176gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G204gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(G120gat), .B(G148gat), .Z(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT66), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(new_n247_), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT65), .Z(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT13), .ZN(new_n253_));
  XOR2_X1   g052(.A(G43gat), .B(G50gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(G29gat), .B(G36gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G29gat), .B(G36gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(G43gat), .B(G50gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G15gat), .B(G22gat), .ZN(new_n262_));
  INV_X1    g061(.A(G1gat), .ZN(new_n263_));
  INV_X1    g062(.A(G8gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT14), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G1gat), .B(G8gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT72), .Z(new_n270_));
  INV_X1    g069(.A(KEYINPUT15), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n257_), .A2(new_n258_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n254_), .A2(new_n255_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT15), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n268_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n270_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(G229gat), .B2(G233gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G229gat), .A2(G233gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n261_), .A2(new_n268_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n280_), .B1(new_n270_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G113gat), .B(G141gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G169gat), .B(G197gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  OR3_X1    g084(.A1(new_n279_), .A2(new_n282_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n285_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n253_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G8gat), .B(G36gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT93), .ZN(new_n294_));
  XOR2_X1   g093(.A(G64gat), .B(G92gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299_));
  INV_X1    g098(.A(G183gat), .ZN(new_n300_));
  INV_X1    g099(.A(G190gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G169gat), .ZN(new_n305_));
  INV_X1    g104(.A(G176gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n307_), .A2(KEYINPUT24), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(KEYINPUT24), .A3(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n304_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT26), .B(G190gat), .Z(new_n313_));
  INV_X1    g112(.A(KEYINPUT88), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(KEYINPUT25), .B(G183gat), .Z(new_n316_));
  OAI21_X1  g115(.A(new_n312_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n309_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT22), .B(G169gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT89), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n318_), .B1(new_n321_), .B2(new_n306_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n302_), .B(new_n303_), .C1(G183gat), .C2(G190gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT90), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n322_), .A2(KEYINPUT91), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT91), .B1(new_n322_), .B2(new_n325_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n317_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT21), .ZN(new_n329_));
  INV_X1    g128(.A(G204gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(G197gat), .ZN(new_n331_));
  INV_X1    g130(.A(G197gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G204gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n329_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT81), .ZN(new_n335_));
  AND2_X1   g134(.A1(G211gat), .A2(G218gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G211gat), .A2(G218gat), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n334_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n334_), .B2(new_n338_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n331_), .A2(new_n333_), .A3(new_n329_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n338_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n331_), .A2(new_n333_), .A3(KEYINPUT79), .A4(new_n329_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n331_), .A2(new_n333_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT21), .ZN(new_n348_));
  AND4_X1   g147(.A1(new_n342_), .A2(new_n345_), .A3(new_n346_), .A4(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n331_), .A2(new_n333_), .A3(new_n329_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n334_), .B1(new_n350_), .B2(KEYINPUT79), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n342_), .B1(new_n351_), .B2(new_n345_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n341_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n328_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT19), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n316_), .A2(new_n313_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n311_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n319_), .A2(new_n306_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n323_), .A3(new_n309_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n353_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT20), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n354_), .A2(new_n356_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT20), .B1(new_n353_), .B2(new_n361_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT87), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(KEYINPUT87), .B(KEYINPUT20), .C1(new_n353_), .C2(new_n361_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n328_), .A2(new_n353_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n356_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n298_), .B(new_n365_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n298_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n364_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n378_), .A2(KEYINPUT27), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n322_), .A2(new_n325_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n317_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT96), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(KEYINPUT96), .A3(new_n317_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT82), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n353_), .A2(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(KEYINPUT82), .B(new_n341_), .C1(new_n349_), .C2(new_n352_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n356_), .B1(new_n389_), .B2(new_n363_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n370_), .A2(KEYINPUT97), .A3(new_n373_), .A4(new_n371_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n371_), .A2(new_n368_), .A3(new_n373_), .A4(new_n369_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT97), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n375_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(KEYINPUT27), .A3(new_n374_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398_));
  OR2_X1    g197(.A1(G155gat), .A2(G162gat), .ZN(new_n399_));
  INV_X1    g198(.A(G141gat), .ZN(new_n400_));
  INV_X1    g199(.A(G148gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT77), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n402_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G141gat), .A2(G148gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n406_), .B(KEYINPUT2), .Z(new_n407_));
  OAI211_X1 g206(.A(new_n398_), .B(new_n399_), .C1(new_n405_), .C2(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n402_), .A2(new_n406_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n398_), .A2(KEYINPUT1), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT1), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(G155gat), .A3(G162gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n412_), .A3(new_n399_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n409_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n408_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G127gat), .B(G134gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G113gat), .B(G120gat), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n419_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(KEYINPUT75), .A3(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(KEYINPUT75), .B2(new_n420_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n417_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n421_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n408_), .B(new_n425_), .C1(new_n416_), .C2(new_n415_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT4), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT94), .Z(new_n430_));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n424_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n430_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G85gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT0), .B(G57gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n438_), .B(new_n439_), .Z(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n433_), .A2(new_n442_), .A3(new_n435_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(KEYINPUT98), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT98), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n436_), .A2(new_n445_), .A3(new_n440_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n379_), .A2(new_n397_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n417_), .A2(KEYINPUT29), .ZN(new_n450_));
  INV_X1    g249(.A(G228gat), .ZN(new_n451_));
  INV_X1    g250(.A(G233gat), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n450_), .B(new_n353_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n387_), .A2(new_n450_), .A3(new_n388_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n451_), .A2(new_n452_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n454_), .A2(KEYINPUT83), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT83), .B1(new_n454_), .B2(new_n455_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n453_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT84), .ZN(new_n459_));
  XOR2_X1   g258(.A(G78gat), .B(G106gat), .Z(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n462_), .B(new_n453_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT85), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n459_), .A2(new_n466_), .A3(new_n461_), .A4(new_n463_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n417_), .A2(KEYINPUT29), .ZN(new_n468_));
  XOR2_X1   g267(.A(G22gat), .B(G50gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(KEYINPUT78), .B(KEYINPUT28), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT86), .B1(new_n458_), .B2(new_n461_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n454_), .A2(new_n455_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n454_), .A2(KEYINPUT83), .A3(new_n455_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n460_), .A4(new_n453_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n472_), .B1(new_n473_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n465_), .A2(new_n467_), .A3(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(new_n460_), .A3(new_n453_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n460_), .B1(new_n478_), .B2(new_n453_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n472_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n423_), .B(KEYINPUT31), .Z(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT74), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G227gat), .A2(G233gat), .ZN(new_n489_));
  INV_X1    g288(.A(G71gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n361_), .B(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n488_), .B(new_n492_), .Z(new_n493_));
  XOR2_X1   g292(.A(KEYINPUT30), .B(G99gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(G15gat), .B(G43gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n493_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n482_), .A2(new_n486_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n498_), .B1(new_n482_), .B2(new_n486_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n449_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n482_), .A2(new_n486_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n497_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n482_), .A2(new_n486_), .A3(new_n498_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n298_), .A2(KEYINPUT32), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n395_), .A2(new_n506_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n365_), .B(new_n505_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n447_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n442_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n511_), .A2(KEYINPUT33), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n510_), .B(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n430_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n427_), .A2(new_n434_), .ZN(new_n515_));
  OR3_X1    g314(.A1(new_n514_), .A2(new_n440_), .A3(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n513_), .A2(new_n374_), .A3(new_n377_), .A4(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n509_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n503_), .A2(new_n504_), .A3(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n501_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n276_), .A2(new_n236_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n260_), .B(new_n226_), .C1(new_n235_), .C2(new_n234_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n524_), .B(KEYINPUT34), .Z(new_n525_));
  INV_X1    g324(.A(KEYINPUT35), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT67), .B1(new_n522_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n276_), .A2(new_n236_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT67), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n523_), .A4(new_n527_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n525_), .A2(new_n526_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n529_), .A2(new_n534_), .A3(new_n532_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(KEYINPUT36), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G190gat), .B(G218gat), .ZN(new_n539_));
  INV_X1    g338(.A(G162gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT68), .B(G134gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT36), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n536_), .A2(new_n548_), .A3(new_n537_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n529_), .A2(new_n534_), .A3(new_n532_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n534_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n549_), .B(new_n546_), .C1(new_n555_), .C2(new_n545_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(KEYINPUT71), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT37), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(KEYINPUT70), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT70), .ZN(new_n560_));
  INV_X1    g359(.A(new_n556_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n549_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n560_), .B1(new_n563_), .B2(KEYINPUT71), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n551_), .A2(new_n560_), .A3(new_n556_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT37), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n559_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n268_), .B(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(new_n207_), .Z(new_n571_));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(G211gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT16), .B(G183gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n575_), .A2(KEYINPUT17), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n575_), .B(KEYINPUT17), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n568_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n292_), .A2(new_n521_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT99), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n263_), .A3(new_n447_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT38), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n563_), .B(KEYINPUT100), .Z(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n521_), .A2(new_n588_), .A3(new_n580_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n291_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(G1gat), .B1(new_n591_), .B2(new_n448_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n586_), .A2(new_n592_), .ZN(G1324gat));
  NAND2_X1  g392(.A1(new_n379_), .A2(new_n397_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n264_), .B1(new_n590_), .B2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT39), .Z(new_n596_));
  NAND3_X1  g395(.A1(new_n584_), .A2(new_n264_), .A3(new_n594_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g398(.A(G15gat), .B1(new_n591_), .B2(new_n497_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT41), .Z(new_n601_));
  OR3_X1    g400(.A1(new_n583_), .A2(G15gat), .A3(new_n497_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(G1326gat));
  INV_X1    g404(.A(new_n502_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G22gat), .B1(new_n591_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT42), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n606_), .A2(G22gat), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n583_), .B2(new_n609_), .ZN(G1327gat));
  NOR2_X1   g409(.A1(new_n291_), .A2(new_n580_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n501_), .A2(new_n520_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n563_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(G29gat), .B1(new_n616_), .B2(new_n447_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT44), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n612_), .A2(KEYINPUT43), .A3(new_n568_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n567_), .A2(KEYINPUT102), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n621_), .B(new_n559_), .C1(new_n564_), .C2(new_n566_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT43), .B1(new_n612_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n501_), .A2(new_n520_), .A3(new_n620_), .A4(new_n622_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(KEYINPUT103), .A3(KEYINPUT43), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n619_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n611_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n618_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n631_), .A2(G29gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n619_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n627_), .A2(KEYINPUT103), .A3(KEYINPUT43), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT103), .B1(new_n627_), .B2(KEYINPUT43), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n633_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(KEYINPUT44), .A3(new_n611_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(new_n447_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n617_), .B1(new_n632_), .B2(new_n638_), .ZN(G1328gat));
  INV_X1    g438(.A(new_n594_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n615_), .A2(G36gat), .A3(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT45), .Z(new_n642_));
  NAND3_X1  g441(.A1(new_n631_), .A2(new_n594_), .A3(new_n637_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(KEYINPUT104), .A3(G36gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT104), .B1(new_n643_), .B2(G36gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT46), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT46), .B(new_n642_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1329gat));
  XNOR2_X1  g449(.A(KEYINPUT105), .B(G43gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n615_), .B2(new_n497_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT106), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n631_), .A2(G43gat), .A3(new_n498_), .A4(new_n637_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g455(.A1(new_n615_), .A2(G50gat), .A3(new_n606_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n631_), .A2(new_n502_), .A3(new_n637_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n658_), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT107), .B1(new_n658_), .B2(G50gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT108), .B(new_n657_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1331gat));
  INV_X1    g464(.A(new_n253_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n582_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT109), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n612_), .A2(new_n290_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT110), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT110), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n668_), .A2(new_n672_), .A3(new_n669_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n671_), .A2(new_n447_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(G57gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n290_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n666_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(new_n589_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(G57gat), .A3(new_n447_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT111), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n676_), .A2(KEYINPUT111), .A3(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1332gat));
  INV_X1    g484(.A(G64gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n679_), .B2(new_n594_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT48), .Z(new_n688_));
  INV_X1    g487(.A(new_n670_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n686_), .A3(new_n594_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1333gat));
  AOI21_X1  g490(.A(new_n490_), .B1(new_n679_), .B2(new_n498_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n498_), .A2(new_n490_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT113), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n670_), .B2(new_n696_), .ZN(G1334gat));
  INV_X1    g496(.A(G78gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n679_), .B2(new_n502_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT50), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n689_), .A2(new_n698_), .A3(new_n502_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1335gat));
  NOR2_X1   g501(.A1(new_n678_), .A2(new_n580_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n636_), .A2(new_n703_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n704_), .A2(KEYINPUT114), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(KEYINPUT114), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n448_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n703_), .A2(new_n614_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n447_), .A2(new_n212_), .ZN(new_n709_));
  OAI22_X1  g508(.A1(new_n707_), .A2(new_n212_), .B1(new_n708_), .B2(new_n709_), .ZN(G1336gat));
  OAI21_X1  g509(.A(new_n213_), .B1(new_n708_), .B2(new_n640_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT115), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n640_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g513(.A(G99gat), .B1(new_n704_), .B2(new_n497_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n498_), .A2(new_n218_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n708_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g517(.A1(new_n703_), .A2(new_n219_), .A3(new_n502_), .A4(new_n614_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G106gat), .B1(new_n704_), .B2(new_n606_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT52), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(KEYINPUT52), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g523(.A1(new_n594_), .A2(new_n448_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n240_), .B(KEYINPUT116), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(G230gat), .A3(G233gat), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT55), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT117), .B1(new_n242_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n242_), .A2(new_n728_), .ZN(new_n730_));
  OR3_X1    g529(.A1(new_n242_), .A2(KEYINPUT117), .A3(new_n728_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n727_), .A2(new_n729_), .A3(new_n730_), .A4(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n247_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT118), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT56), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(KEYINPUT56), .A3(new_n247_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n734_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n290_), .B(new_n249_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n270_), .A2(new_n281_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n280_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n278_), .B(KEYINPUT119), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n285_), .B(new_n742_), .C1(new_n743_), .C2(new_n280_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT120), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(new_n286_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n252_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n740_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT57), .B1(new_n748_), .B2(new_n613_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT57), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n750_), .B(new_n563_), .C1(new_n740_), .C2(new_n747_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n733_), .A2(new_n735_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT121), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n737_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n732_), .A2(KEYINPUT121), .A3(KEYINPUT56), .A4(new_n247_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(new_n249_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n757_), .A3(new_n746_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT122), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT58), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT58), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(new_n759_), .A3(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n761_), .A2(new_n567_), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n580_), .B1(new_n752_), .B2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n253_), .A2(new_n582_), .A3(new_n677_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n766_), .A2(KEYINPUT54), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(KEYINPUT54), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n499_), .B(new_n725_), .C1(new_n765_), .C2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G113gat), .B1(new_n772_), .B2(new_n290_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(KEYINPUT59), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n748_), .A2(new_n613_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n750_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n748_), .A2(KEYINPUT57), .A3(new_n613_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n764_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n580_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n769_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT59), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n499_), .A4(new_n725_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n774_), .A2(G113gat), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n773_), .B1(new_n784_), .B2(new_n290_), .ZN(G1340gat));
  INV_X1    g584(.A(G120gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n253_), .B2(KEYINPUT60), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n772_), .B(new_n787_), .C1(KEYINPUT60), .C2(new_n786_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n774_), .A2(new_n666_), .A3(new_n783_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n786_), .ZN(G1341gat));
  AND4_X1   g589(.A1(G127gat), .A2(new_n774_), .A3(new_n580_), .A4(new_n783_), .ZN(new_n791_));
  AOI21_X1  g590(.A(G127gat), .B1(new_n772_), .B2(new_n580_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1342gat));
  AND4_X1   g592(.A1(G134gat), .A2(new_n774_), .A3(new_n567_), .A4(new_n783_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G134gat), .B1(new_n772_), .B2(new_n587_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1343gat));
  OAI211_X1 g595(.A(new_n500_), .B(new_n725_), .C1(new_n765_), .C2(new_n770_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n677_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(new_n400_), .ZN(G1344gat));
  NOR2_X1   g598(.A1(new_n797_), .A2(new_n253_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(new_n401_), .ZN(G1345gat));
  XNOR2_X1  g600(.A(KEYINPUT61), .B(G155gat), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n778_), .A2(new_n779_), .B1(new_n768_), .B2(new_n767_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n725_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n503_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n804_), .B1(new_n807_), .B2(new_n580_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n797_), .A2(KEYINPUT123), .A3(new_n779_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n803_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(new_n804_), .A3(new_n580_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT123), .B1(new_n797_), .B2(new_n779_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n802_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(G1346gat));
  AOI21_X1  g613(.A(G162gat), .B1(new_n807_), .B2(new_n587_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n797_), .A2(new_n540_), .A3(new_n623_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1347gat));
  NOR2_X1   g616(.A1(new_n640_), .A2(new_n447_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NOR4_X1   g618(.A1(new_n805_), .A2(new_n677_), .A3(new_n504_), .A4(new_n819_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n820_), .A2(KEYINPUT62), .A3(new_n305_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT62), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n820_), .B2(new_n321_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n781_), .A2(new_n499_), .A3(new_n818_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G169gat), .B1(new_n824_), .B2(new_n677_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n821_), .B1(new_n823_), .B2(new_n825_), .ZN(G1348gat));
  NOR2_X1   g625(.A1(new_n824_), .A2(new_n253_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(new_n306_), .ZN(G1349gat));
  NOR2_X1   g627(.A1(new_n824_), .A2(new_n779_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n316_), .B1(new_n830_), .B2(new_n300_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n830_), .A2(G183gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n829_), .B2(new_n833_), .ZN(G1350gat));
  OAI21_X1  g633(.A(G190gat), .B1(new_n824_), .B2(new_n568_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n588_), .A2(new_n315_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n824_), .B2(new_n836_), .ZN(G1351gat));
  NOR3_X1   g636(.A1(new_n805_), .A2(new_n503_), .A3(new_n819_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n290_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n838_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n677_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT125), .B(G197gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n840_), .B1(new_n842_), .B2(new_n843_), .ZN(G1352gat));
  NOR2_X1   g643(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n845_));
  AND2_X1   g644(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n838_), .B(new_n666_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n841_), .A2(new_n253_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n845_), .ZN(G1353gat));
  XNOR2_X1  g648(.A(KEYINPUT63), .B(G211gat), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n841_), .A2(new_n779_), .A3(new_n850_), .ZN(new_n851_));
  AOI211_X1 g650(.A(KEYINPUT63), .B(G211gat), .C1(new_n838_), .C2(new_n580_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1354gat));
  AND2_X1   g652(.A1(new_n567_), .A2(G218gat), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n781_), .A2(new_n500_), .A3(new_n818_), .A4(new_n854_), .ZN(new_n855_));
  NOR4_X1   g654(.A1(new_n805_), .A2(new_n588_), .A3(new_n503_), .A4(new_n819_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(G218gat), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT127), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT127), .B(new_n855_), .C1(new_n856_), .C2(G218gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1355gat));
endmodule


