//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT36), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(G99gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT10), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT10), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G99gat), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT64), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT64), .B1(new_n209_), .B2(new_n211_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n207_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  AND3_X1   g013(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT65), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  INV_X1    g020(.A(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT9), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n218_), .A2(KEYINPUT65), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n220_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n214_), .A2(new_n217_), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G29gat), .B(G36gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G43gat), .B(G50gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n232_), .B(new_n233_), .C1(G99gat), .C2(G106gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n208_), .B(new_n207_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT6), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(KEYINPUT67), .A3(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n236_), .A2(new_n238_), .A3(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n223_), .A2(new_n218_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n231_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n223_), .A2(new_n231_), .A3(new_n218_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(new_n236_), .B2(new_n217_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n227_), .B(new_n230_), .C1(new_n246_), .C2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G232gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT34), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT35), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n227_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n244_), .A2(new_n245_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT8), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n259_));
  INV_X1    g058(.A(new_n248_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT69), .B1(new_n246_), .B2(new_n248_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n256_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n230_), .B(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n255_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n252_), .A2(new_n253_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n255_), .B(new_n269_), .C1(new_n263_), .C2(new_n265_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n206_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT76), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT77), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT37), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT36), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n204_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n268_), .A2(new_n270_), .A3(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .A4(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT74), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n268_), .A2(new_n281_), .A3(new_n270_), .A4(new_n277_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n268_), .A2(new_n270_), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT75), .B1(new_n284_), .B2(new_n205_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n286_));
  AOI211_X1 g085(.A(new_n286_), .B(new_n206_), .C1(new_n268_), .C2(new_n270_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n274_), .B1(new_n283_), .B2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n259_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n246_), .A2(KEYINPUT69), .A3(new_n248_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n227_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n265_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n269_), .B1(new_n294_), .B2(new_n255_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n270_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n205_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT76), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n284_), .A2(new_n299_), .A3(new_n205_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n298_), .A2(new_n274_), .A3(new_n278_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT77), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n279_), .B1(new_n289_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT78), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT78), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n279_), .B(new_n305_), .C1(new_n289_), .C2(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n227_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G57gat), .B(G64gat), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(KEYINPUT11), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(KEYINPUT11), .ZN(new_n311_));
  XOR2_X1   g110(.A(G71gat), .B(G78gat), .Z(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n311_), .A2(new_n312_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n308_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT71), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n322_), .A3(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n261_), .A2(new_n262_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n315_), .B1(new_n324_), .B2(new_n227_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n321_), .A2(new_n323_), .B1(new_n325_), .B2(KEYINPUT12), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n258_), .A2(new_n260_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(new_n227_), .A3(new_n315_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G230gat), .A2(G233gat), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n326_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n292_), .A2(KEYINPUT12), .A3(new_n316_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n322_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n334_));
  AOI211_X1 g133(.A(KEYINPUT71), .B(new_n318_), .C1(new_n308_), .C2(new_n316_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n333_), .B(new_n331_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT72), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n332_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n329_), .A2(new_n339_), .A3(new_n317_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n308_), .A2(KEYINPUT68), .A3(new_n316_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n330_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n338_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G120gat), .B(G148gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(G204gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT5), .B(G176gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n349_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n338_), .A2(new_n344_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT13), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(KEYINPUT13), .A3(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G15gat), .B(G22gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT79), .ZN(new_n359_));
  INV_X1    g158(.A(G1gat), .ZN(new_n360_));
  INV_X1    g159(.A(G8gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT14), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT80), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G1gat), .B(G8gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(new_n230_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G229gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n366_), .A2(new_n265_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n230_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n368_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G113gat), .B(G141gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G169gat), .B(G197gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT81), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n374_), .B(new_n378_), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n357_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n366_), .B(new_n315_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G231gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT17), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G127gat), .B(G155gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G211gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(KEYINPUT16), .B(G183gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  OR3_X1    g189(.A1(new_n385_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(KEYINPUT17), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n385_), .A2(new_n392_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G113gat), .B(G120gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G127gat), .B(G134gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n399_), .A2(new_n400_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n399_), .A2(new_n400_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(KEYINPUT85), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT2), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n410_));
  OAI22_X1  g209(.A1(new_n407_), .A2(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n408_), .B2(new_n407_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n410_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT88), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n418_), .A2(KEYINPUT1), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n418_), .A2(KEYINPUT1), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n415_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G141gat), .B(G148gat), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n419_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n403_), .A2(new_n406_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n422_), .A2(new_n424_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(new_n401_), .A3(new_n419_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n427_), .B1(new_n426_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n396_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n426_), .A2(new_n395_), .A3(new_n430_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(new_n221_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT0), .B(G57gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n432_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT27), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G211gat), .B(G218gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT92), .ZN(new_n444_));
  INV_X1    g243(.A(G197gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(G204gat), .ZN(new_n446_));
  INV_X1    g245(.A(G204gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(G197gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT21), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT91), .B1(new_n447_), .B2(G197gat), .ZN(new_n450_));
  MUX2_X1   g249(.A(new_n450_), .B(KEYINPUT91), .S(new_n446_), .Z(new_n451_));
  OAI211_X1 g250(.A(new_n444_), .B(new_n449_), .C1(new_n451_), .C2(KEYINPUT21), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT92), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n443_), .B(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n451_), .A3(KEYINPUT21), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G183gat), .A2(G190gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT23), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT23), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(G183gat), .A3(G190gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  OR3_X1    g260(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(G169gat), .ZN(new_n465_));
  INV_X1    g264(.A(G176gat), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n466_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(KEYINPUT24), .A3(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT82), .B(G190gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT26), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT25), .B(G183gat), .ZN(new_n474_));
  INV_X1    g273(.A(G190gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n474_), .B1(KEYINPUT26), .B2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n464_), .B(new_n470_), .C1(new_n473_), .C2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n461_), .B1(new_n471_), .B2(G183gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT22), .B(G169gat), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n467_), .B1(new_n479_), .B2(new_n466_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n456_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n472_), .A2(G190gat), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n476_), .A2(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n463_), .A2(KEYINPUT93), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n463_), .A2(KEYINPUT93), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n470_), .A4(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n480_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G183gat), .A2(G190gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n488_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n483_), .B(KEYINPUT20), .C1(new_n492_), .C2(new_n456_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G226gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT19), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n456_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n456_), .A2(new_n482_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT20), .A4(new_n495_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G8gat), .B(G36gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT95), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G64gat), .B(G92gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n442_), .B1(new_n501_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n493_), .A2(new_n495_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT20), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n510_), .B1(new_n495_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n507_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT97), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n509_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n501_), .A2(new_n508_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n497_), .A2(new_n507_), .A3(new_n500_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT27), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n515_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT86), .B1(new_n403_), .B2(new_n406_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT31), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n403_), .A2(KEYINPUT86), .A3(new_n406_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G15gat), .B(G43gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n477_), .A2(new_n529_), .A3(new_n481_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n529_), .B1(new_n477_), .B2(new_n481_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n482_), .A2(KEYINPUT30), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n530_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n528_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n532_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n536_), .A2(new_n535_), .A3(new_n530_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n528_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n538_), .A2(G227gat), .A3(G233gat), .A4(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G227gat), .A2(G233gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n542_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n541_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n527_), .A2(KEYINPUT87), .A3(new_n543_), .A4(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n543_), .A3(KEYINPUT87), .ZN(new_n549_));
  INV_X1    g348(.A(new_n526_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G22gat), .B(G50gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G78gat), .B(G106gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT28), .B1(new_n425_), .B2(KEYINPUT29), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT29), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n429_), .A2(new_n559_), .A3(new_n560_), .A4(new_n419_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n425_), .A2(KEYINPUT29), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n558_), .A2(new_n561_), .A3(new_n562_), .A4(new_n456_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n558_), .A2(new_n561_), .B1(new_n562_), .B2(new_n456_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G228gat), .A2(G233gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT90), .Z(new_n567_));
  NOR3_X1   g366(.A1(new_n564_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n567_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n558_), .A2(new_n561_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n562_), .A2(new_n456_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n569_), .B1(new_n572_), .B2(new_n563_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n557_), .B1(new_n568_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n567_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n556_), .A3(new_n576_), .ZN(new_n577_));
  AND4_X1   g376(.A1(new_n548_), .A2(new_n553_), .A3(new_n574_), .A4(new_n577_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n548_), .A2(new_n553_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n441_), .B(new_n520_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n432_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT33), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n517_), .A2(new_n518_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n426_), .A2(new_n396_), .A3(new_n430_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n437_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT96), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n395_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(KEYINPUT96), .A3(new_n437_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n432_), .A2(KEYINPUT33), .A3(new_n433_), .A4(new_n438_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n583_), .A2(new_n584_), .A3(new_n591_), .A4(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT32), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n501_), .B1(new_n594_), .B2(new_n507_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n512_), .A2(KEYINPUT32), .A3(new_n508_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n595_), .B(new_n596_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n548_), .A2(new_n553_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n574_), .A2(new_n577_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n580_), .A2(new_n601_), .ZN(new_n602_));
  AND4_X1   g401(.A1(new_n307_), .A2(new_n381_), .A3(new_n394_), .A4(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT98), .ZN(new_n604_));
  INV_X1    g403(.A(new_n441_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n360_), .A3(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n381_), .A2(new_n602_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n394_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n272_), .A2(new_n278_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n611_), .A2(KEYINPUT101), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(KEYINPUT101), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n609_), .A2(new_n610_), .A3(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n616_), .A2(new_n605_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n606_), .A2(new_n607_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(KEYINPUT100), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(KEYINPUT100), .ZN(new_n620_));
  OAI221_X1 g419(.A(new_n608_), .B1(new_n360_), .B2(new_n617_), .C1(new_n619_), .C2(new_n620_), .ZN(G1324gat));
  XNOR2_X1  g420(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n520_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n361_), .B1(new_n616_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT39), .Z(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n604_), .A2(new_n361_), .A3(new_n624_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n627_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n623_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n628_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT40), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n622_), .A3(new_n629_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n599_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n616_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT41), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n604_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1326gat));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n600_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n616_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT42), .Z(new_n646_));
  NOR2_X1   g445(.A1(new_n600_), .A2(G22gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT104), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n604_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT105), .Z(G1327gat));
  NAND2_X1  g450(.A1(new_n615_), .A2(new_n610_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n609_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT107), .ZN(new_n654_));
  INV_X1    g453(.A(G29gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n605_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n602_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT43), .ZN(new_n658_));
  INV_X1    g457(.A(new_n306_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n297_), .A2(new_n286_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n271_), .A2(KEYINPUT75), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n280_), .A4(new_n282_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT37), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(KEYINPUT77), .A3(new_n301_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n305_), .B1(new_n664_), .B2(new_n279_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n659_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n602_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n658_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n610_), .A3(new_n381_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n669_), .A2(KEYINPUT44), .A3(new_n610_), .A4(new_n381_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n605_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT106), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n656_), .B1(new_n676_), .B2(new_n655_), .ZN(G1328gat));
  NAND3_X1  g476(.A1(new_n672_), .A2(new_n624_), .A3(new_n673_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT108), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n672_), .A2(new_n680_), .A3(new_n624_), .A4(new_n673_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(G36gat), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n654_), .A2(new_n683_), .A3(new_n624_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT45), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n682_), .A2(new_n685_), .A3(KEYINPUT46), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1329gat));
  INV_X1    g489(.A(G43gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n654_), .A2(new_n691_), .A3(new_n638_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n674_), .A2(new_n638_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n691_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n692_), .B(KEYINPUT47), .C1(new_n693_), .C2(new_n691_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1330gat));
  INV_X1    g497(.A(G50gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n654_), .A2(new_n699_), .A3(new_n644_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n674_), .A2(new_n644_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n703_), .B2(new_n699_), .ZN(G1331gat));
  INV_X1    g503(.A(new_n357_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n379_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(new_n602_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n707_), .A2(new_n307_), .A3(new_n394_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G57gat), .B1(new_n708_), .B2(new_n605_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n707_), .A2(new_n394_), .A3(new_n614_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n605_), .A2(G57gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(G1332gat));
  INV_X1    g511(.A(G64gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n708_), .A2(new_n713_), .A3(new_n624_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n710_), .A2(new_n624_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G64gat), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n716_), .A2(KEYINPUT110), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(KEYINPUT110), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n717_), .A2(new_n718_), .A3(KEYINPUT48), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n714_), .B1(new_n721_), .B2(new_n722_), .ZN(G1333gat));
  INV_X1    g522(.A(G71gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n710_), .B2(new_n638_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n708_), .A2(new_n724_), .A3(new_n638_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1334gat));
  INV_X1    g528(.A(G78gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n710_), .B2(new_n644_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT50), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n708_), .A2(new_n730_), .A3(new_n644_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1335gat));
  AND3_X1   g533(.A1(new_n707_), .A2(new_n610_), .A3(new_n615_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n605_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n658_), .A2(new_n668_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(KEYINPUT112), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n705_), .A2(new_n394_), .A3(new_n379_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(KEYINPUT112), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n742_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n441_), .A2(new_n221_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT114), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n736_), .B1(new_n745_), .B2(new_n747_), .ZN(G1336gat));
  NAND3_X1  g547(.A1(new_n735_), .A2(new_n222_), .A3(new_n624_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n520_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(new_n222_), .ZN(G1337gat));
  OAI21_X1  g550(.A(G99gat), .B1(new_n741_), .B2(new_n599_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n735_), .B(new_n638_), .C1(new_n213_), .C2(new_n212_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g554(.A1(new_n669_), .A2(new_n610_), .A3(new_n644_), .A4(new_n706_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(G106gat), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT52), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n735_), .A2(new_n207_), .A3(new_n644_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g560(.A(new_n579_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n379_), .A2(new_n352_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT55), .B1(new_n332_), .B2(new_n337_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n336_), .B2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n326_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n331_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n333_), .B(new_n329_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n321_), .A2(new_n323_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n774_), .A2(KEYINPUT115), .A3(new_n329_), .A4(new_n333_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n330_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n765_), .A2(new_n770_), .A3(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n764_), .B1(new_n777_), .B2(new_n351_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n768_), .A2(new_n769_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n327_), .B1(new_n326_), .B2(new_n331_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n336_), .A2(KEYINPUT72), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n767_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT115), .B1(new_n326_), .B2(new_n329_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n334_), .A2(new_n335_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT12), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n263_), .A2(new_n785_), .A3(new_n315_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n329_), .ZN(new_n787_));
  NOR4_X1   g586(.A1(new_n784_), .A2(new_n786_), .A3(new_n772_), .A4(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n342_), .B1(new_n783_), .B2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n779_), .A2(new_n782_), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n349_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n763_), .B1(new_n778_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n371_), .A2(new_n372_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT117), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n371_), .A2(new_n795_), .A3(new_n372_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n368_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n367_), .A2(new_n369_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n377_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n374_), .A2(new_n377_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n614_), .B1(new_n792_), .B2(new_n802_), .ZN(new_n803_));
  XOR2_X1   g602(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n343_), .B(new_n349_), .C1(new_n332_), .C2(new_n337_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n801_), .B2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n352_), .A2(KEYINPUT119), .A3(new_n799_), .A4(new_n800_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n349_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n349_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n810_), .B(KEYINPUT58), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n666_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT57), .B(new_n614_), .C1(new_n792_), .C2(new_n802_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n805_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n610_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n307_), .A2(new_n394_), .A3(new_n380_), .A4(new_n705_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT54), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n762_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n624_), .A2(new_n441_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G113gat), .B1(new_n826_), .B2(new_n379_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT59), .B1(new_n823_), .B2(new_n824_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n380_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n827_), .B1(new_n833_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g633(.A(new_n357_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n705_), .B2(G120gat), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n826_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G120gat), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1341gat));
  AOI21_X1  g640(.A(G127gat), .B1(new_n826_), .B2(new_n394_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n610_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g643(.A(G134gat), .B1(new_n826_), .B2(new_n615_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n307_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g646(.A1(new_n820_), .A2(new_n822_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n848_), .A2(new_n578_), .A3(new_n824_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n379_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n357_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n394_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1346gat));
  AND2_X1   g655(.A1(new_n666_), .A2(G162gat), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n849_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G162gat), .B1(new_n849_), .B2(new_n615_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT120), .B1(new_n858_), .B2(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n520_), .A2(new_n605_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n848_), .A2(new_n379_), .A3(new_n579_), .A4(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n465_), .B1(new_n867_), .B2(KEYINPUT62), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n867_), .A2(KEYINPUT62), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n823_), .A2(new_n865_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n379_), .A3(new_n479_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n866_), .B(new_n868_), .C1(new_n867_), .C2(KEYINPUT62), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n871_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT122), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n871_), .A2(new_n873_), .A3(new_n874_), .A4(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1348gat));
  NAND2_X1  g678(.A1(new_n872_), .A2(new_n357_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g680(.A1(new_n872_), .A2(new_n394_), .A3(new_n474_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n823_), .A2(new_n394_), .A3(new_n865_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G183gat), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n882_), .A2(new_n883_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n883_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1350gat));
  INV_X1    g687(.A(new_n872_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G190gat), .B1(new_n889_), .B2(new_n307_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n872_), .B(new_n615_), .C1(KEYINPUT26), .C2(new_n475_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n484_), .ZN(G1351gat));
  AND2_X1   g691(.A1(new_n848_), .A2(new_n578_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(new_n379_), .A3(new_n865_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n894_), .A2(new_n895_), .A3(new_n445_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n894_), .B2(new_n445_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n894_), .A2(new_n445_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(G1352gat));
  AND2_X1   g698(.A1(new_n893_), .A2(new_n865_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n357_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g701(.A(KEYINPUT63), .ZN(new_n903_));
  INV_X1    g702(.A(G211gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n394_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n905_), .A2(new_n906_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n893_), .A2(new_n865_), .A3(new_n907_), .A4(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n903_), .A2(new_n904_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1354gat));
  NAND2_X1  g710(.A1(new_n900_), .A2(new_n615_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT126), .B(G218gat), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n307_), .A2(new_n913_), .ZN(new_n914_));
  AOI22_X1  g713(.A1(new_n912_), .A2(new_n913_), .B1(new_n900_), .B2(new_n914_), .ZN(G1355gat));
endmodule


