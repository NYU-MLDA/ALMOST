//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n993_, new_n995_,
    new_n997_, new_n998_, new_n1000_, new_n1001_, new_n1002_, new_n1004_,
    new_n1005_, new_n1006_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT23), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G183gat), .A3(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n209_), .A2(KEYINPUT84), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n205_), .A2(new_n207_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n212_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT84), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220_));
  OAI21_X1  g019(.A(G169gat), .B1(new_n220_), .B2(KEYINPUT82), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT82), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT22), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT83), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n221_), .A2(new_n224_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n221_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n228_));
  AOI22_X1  g027(.A1(new_n228_), .A2(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n219_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT85), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT25), .B(G183gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT26), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT80), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT26), .B(G190gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n232_), .B(new_n235_), .C1(new_n236_), .C2(KEYINPUT80), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G169gat), .A2(G176gat), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n239_), .A2(KEYINPUT24), .A3(new_n240_), .A4(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n237_), .A2(new_n209_), .A3(new_n243_), .A4(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n230_), .A2(new_n231_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n231_), .B1(new_n230_), .B2(new_n246_), .ZN(new_n248_));
  INV_X1    g047(.A(G218gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G211gat), .ZN(new_n250_));
  INV_X1    g049(.A(G211gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G218gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT97), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT97), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT21), .ZN(new_n258_));
  INV_X1    g057(.A(G197gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT95), .ZN(new_n260_));
  INV_X1    g059(.A(G204gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(KEYINPUT95), .A2(G204gat), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n259_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G197gat), .A2(G204gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n258_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n258_), .B1(G197gat), .B2(G204gat), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n267_), .A2(KEYINPUT96), .A3(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT96), .B1(new_n267_), .B2(new_n268_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n257_), .B(new_n266_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n264_), .A2(new_n265_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n272_), .A2(KEYINPUT21), .A3(new_n256_), .A4(new_n254_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n247_), .A2(new_n248_), .A3(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n271_), .A2(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n209_), .A2(new_n212_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT22), .B(G169gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n226_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n244_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n242_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n282_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n211_), .A2(KEYINPUT26), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n210_), .A2(KEYINPUT25), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G183gat), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n234_), .A2(new_n284_), .A3(new_n285_), .A4(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(new_n245_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT98), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT98), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n283_), .A2(new_n291_), .A3(new_n245_), .A4(new_n288_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n281_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT20), .B1(new_n276_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n204_), .B1(new_n275_), .B2(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G8gat), .B(G36gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT18), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n274_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n204_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT20), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n276_), .B2(new_n293_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n295_), .A2(new_n299_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT101), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n299_), .B(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n213_), .A2(new_n218_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n228_), .A2(KEYINPUT83), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n244_), .A3(new_n227_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n246_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT85), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n230_), .A2(new_n231_), .A3(new_n246_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n276_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n280_), .A2(new_n289_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT20), .B1(new_n274_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n204_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n313_), .A3(new_n276_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT20), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n290_), .A2(new_n292_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n280_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n319_), .B1(new_n321_), .B2(new_n274_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n322_), .A3(new_n301_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n307_), .B1(new_n317_), .B2(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(KEYINPUT27), .B(new_n305_), .C1(new_n324_), .C2(KEYINPUT102), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT102), .ZN(new_n326_));
  AOI211_X1 g125(.A(new_n326_), .B(new_n307_), .C1(new_n317_), .C2(new_n323_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n202_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n307_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n323_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n316_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n301_), .B1(new_n300_), .B2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n329_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n326_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n324_), .A2(KEYINPUT102), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n318_), .A2(new_n322_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n337_), .A2(new_n204_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n338_), .B2(new_n299_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n334_), .A2(KEYINPUT103), .A3(new_n335_), .A4(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n328_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n312_), .A2(KEYINPUT30), .A3(new_n313_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G71gat), .B(G99gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(G43gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G227gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(G15gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n348_), .B(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT31), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT31), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n346_), .A2(new_n354_), .A3(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n343_), .A2(new_n345_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT86), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G127gat), .B(G134gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G113gat), .B(G120gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n361_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT87), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(KEYINPUT87), .A3(new_n364_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n358_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n368_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n357_), .A2(KEYINPUT86), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n356_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n375_));
  AND2_X1   g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(KEYINPUT91), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT88), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT88), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(G141gat), .A3(G148gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT2), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n389_));
  INV_X1    g188(.A(G141gat), .ZN(new_n390_));
  INV_X1    g189(.A(G148gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n378_), .B(new_n381_), .C1(new_n388_), .C2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n380_), .B1(new_n377_), .B2(KEYINPUT1), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n398_), .A2(KEYINPUT89), .A3(G155gat), .A4(G162gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n380_), .B2(KEYINPUT1), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(G141gat), .A2(G148gat), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n383_), .A2(new_n385_), .A3(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n402_), .A2(KEYINPUT90), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT90), .B1(new_n402_), .B2(new_n404_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n365_), .B(new_n396_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n381_), .A2(new_n378_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n395_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n387_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n402_), .A2(new_n404_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n402_), .A2(KEYINPUT90), .A3(new_n404_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n410_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(KEYINPUT4), .B(new_n407_), .C1(new_n415_), .C2(new_n371_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n396_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n369_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n416_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n369_), .A2(new_n418_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n407_), .A3(new_n420_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G85gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT0), .B(G57gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n422_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n353_), .A2(new_n370_), .A3(new_n355_), .A4(new_n372_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n374_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n438_), .B(new_n396_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT92), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n413_), .A2(new_n414_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT92), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(new_n438_), .A4(new_n396_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n437_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G22gat), .B(G50gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n440_), .A2(new_n443_), .A3(new_n437_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n446_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n440_), .A2(new_n443_), .A3(new_n437_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n449_), .B1(new_n450_), .B2(new_n444_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT94), .B1(new_n271_), .B2(new_n273_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(G106gat), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n274_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G106gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n453_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n438_), .B1(new_n441_), .B2(new_n396_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n460_), .A2(new_n276_), .A3(G78gat), .ZN(new_n461_));
  INV_X1    g260(.A(G78gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n418_), .A2(KEYINPUT29), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(new_n274_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n455_), .B(new_n459_), .C1(new_n461_), .C2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(G78gat), .B1(new_n460_), .B2(new_n276_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n463_), .A2(new_n462_), .A3(new_n274_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n458_), .B1(new_n457_), .B2(new_n453_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n452_), .A2(G106gat), .A3(new_n454_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n466_), .B(new_n467_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  AND4_X1   g269(.A1(new_n448_), .A2(new_n451_), .A3(new_n465_), .A4(new_n470_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n448_), .A2(new_n451_), .B1(new_n465_), .B2(new_n470_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT99), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n305_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n338_), .A2(KEYINPUT99), .A3(new_n299_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n295_), .A2(new_n304_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n299_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n475_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n336_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n341_), .A2(new_n435_), .A3(new_n473_), .A4(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n433_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n483_), .B1(new_n336_), .B2(new_n480_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n431_), .A2(new_n432_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT32), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n338_), .B1(new_n486_), .B2(new_n478_), .ZN(new_n487_));
  OAI211_X1 g286(.A(KEYINPUT32), .B(new_n299_), .C1(new_n330_), .C2(new_n332_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT33), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n423_), .A2(new_n407_), .A3(new_n421_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n491_), .A2(new_n430_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n432_), .A2(new_n490_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n422_), .A2(new_n424_), .A3(KEYINPUT33), .A4(new_n429_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n495_), .A2(KEYINPUT100), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(KEYINPUT100), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n494_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n489_), .B1(new_n498_), .B2(new_n480_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n484_), .A2(new_n341_), .B1(new_n499_), .B2(new_n473_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n374_), .A2(new_n434_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n482_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT104), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT77), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G29gat), .B(G36gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G43gat), .B(G50gat), .Z(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G1gat), .B(G8gat), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516_));
  INV_X1    g315(.A(G1gat), .ZN(new_n517_));
  INV_X1    g316(.A(G8gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n514_), .A2(new_n519_), .A3(new_n516_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n505_), .B1(new_n513_), .B2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n512_), .A2(new_n522_), .A3(KEYINPUT77), .A4(new_n521_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n513_), .A2(KEYINPUT15), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n512_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n523_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT78), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n526_), .A2(new_n530_), .A3(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G113gat), .B(G141gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT79), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G169gat), .B(G197gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n513_), .A2(new_n523_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n526_), .A2(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n533_), .B(new_n537_), .C1(new_n539_), .C2(new_n531_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n537_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n526_), .A2(new_n530_), .A3(new_n532_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n531_), .B1(new_n526_), .B2(new_n538_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n503_), .A2(new_n504_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n504_), .B1(new_n503_), .B2(new_n546_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(G85gat), .ZN(new_n551_));
  INV_X1    g350(.A(G92gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n553_), .A2(KEYINPUT67), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT6), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT6), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(G99gat), .A3(G106gat), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n561_));
  INV_X1    g360(.A(G99gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n458_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n555_), .B1(new_n560_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT8), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n557_), .A2(new_n559_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(new_n564_), .A3(new_n563_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT8), .A3(new_n555_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT10), .B(G99gat), .Z(new_n573_));
  AOI22_X1  g372(.A1(new_n573_), .A2(new_n458_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT66), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n553_), .A2(KEYINPUT9), .A3(new_n554_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(G85gat), .A3(G92gat), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n575_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n554_), .A2(KEYINPUT9), .ZN(new_n580_));
  NOR2_X1   g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n575_), .B(new_n578_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n574_), .B1(new_n579_), .B2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n584_), .A2(KEYINPUT70), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(KEYINPUT70), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n572_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT12), .ZN(new_n588_));
  XOR2_X1   g387(.A(KEYINPUT68), .B(G71gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(G57gat), .B(G64gat), .ZN(new_n590_));
  OAI22_X1  g389(.A1(new_n589_), .A2(G78gat), .B1(new_n590_), .B2(KEYINPUT11), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT68), .B(G71gat), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n462_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT69), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n590_), .B2(KEYINPUT11), .ZN(new_n595_));
  INV_X1    g394(.A(G64gat), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(G57gat), .ZN(new_n597_));
  INV_X1    g396(.A(G57gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(G64gat), .ZN(new_n599_));
  AND4_X1   g398(.A1(new_n594_), .A2(new_n597_), .A3(new_n599_), .A4(KEYINPUT11), .ZN(new_n600_));
  OAI22_X1  g399(.A1(new_n591_), .A2(new_n593_), .B1(new_n595_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n597_), .A2(new_n599_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT11), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n602_), .A2(new_n603_), .B1(new_n592_), .B2(new_n462_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT69), .B1(new_n602_), .B2(new_n603_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n590_), .A2(new_n594_), .A3(KEYINPUT11), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n589_), .A2(G78gat), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .A4(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n588_), .B1(new_n601_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n587_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n584_), .A2(new_n568_), .A3(new_n571_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n601_), .A2(new_n608_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT64), .B(KEYINPUT65), .Z(new_n614_));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n611_), .A2(new_n612_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT71), .B1(new_n618_), .B2(new_n588_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT71), .ZN(new_n620_));
  AOI211_X1 g419(.A(new_n620_), .B(KEYINPUT12), .C1(new_n611_), .C2(new_n612_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n610_), .B(new_n617_), .C1(new_n619_), .C2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n611_), .A2(new_n612_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n616_), .B1(new_n623_), .B2(new_n613_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT5), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n626_), .B(new_n627_), .Z(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n622_), .A2(new_n624_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT72), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n622_), .A2(KEYINPUT72), .A3(new_n624_), .A4(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n622_), .A2(new_n624_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n635_), .B2(new_n629_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT13), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT34), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT35), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT73), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(KEYINPUT73), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n527_), .A2(new_n529_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n584_), .B(KEYINPUT70), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(new_n572_), .ZN(new_n648_));
  OAI22_X1  g447(.A1(new_n611_), .A2(new_n513_), .B1(KEYINPUT35), .B2(new_n640_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n644_), .B(new_n645_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n646_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n587_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n649_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n652_), .A2(KEYINPUT73), .A3(new_n643_), .A4(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n650_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G134gat), .B(G162gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(KEYINPUT36), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n658_), .A2(KEYINPUT36), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n655_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT74), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n655_), .A2(new_n662_), .A3(new_n659_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n655_), .B2(new_n659_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT37), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(G231gat), .A2(G233gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n523_), .B(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(new_n612_), .Z(new_n670_));
  XOR2_X1   g469(.A(G127gat), .B(G155gat), .Z(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT16), .ZN(new_n672_));
  XNOR2_X1  g471(.A(G183gat), .B(G211gat), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT17), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n670_), .A2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT76), .Z(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n670_), .A2(new_n674_), .A3(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n661_), .B(KEYINPUT37), .C1(new_n664_), .C2(new_n663_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n667_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n638_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n550_), .A2(KEYINPUT105), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT105), .B1(new_n550_), .B2(new_n684_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT38), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n485_), .A2(KEYINPUT106), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n485_), .A2(KEYINPUT106), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n517_), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n687_), .A2(new_n688_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n499_), .A2(new_n473_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n328_), .A2(new_n340_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n483_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n481_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n448_), .A2(new_n451_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n465_), .A2(new_n470_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n448_), .A2(new_n451_), .A3(new_n465_), .A4(new_n470_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AOI221_X4 g502(.A(new_n703_), .B1(new_n480_), .B2(new_n336_), .C1(new_n328_), .C2(new_n340_), .ZN(new_n704_));
  AOI22_X1  g503(.A1(new_n698_), .A2(new_n501_), .B1(new_n704_), .B2(new_n435_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n665_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n636_), .B(KEYINPUT13), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n546_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n680_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G1gat), .B1(new_n712_), .B2(new_n433_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n688_), .B1(new_n687_), .B2(new_n692_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n693_), .A2(new_n713_), .A3(new_n714_), .ZN(G1324gat));
  NAND2_X1  g514(.A1(new_n341_), .A2(new_n481_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n685_), .A2(new_n518_), .A3(new_n716_), .A4(new_n686_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n716_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G8gat), .B1(new_n712_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT39), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT40), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n717_), .A2(KEYINPUT40), .A3(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1325gat));
  OAI21_X1  g524(.A(G15gat), .B1(new_n712_), .B2(new_n501_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT41), .Z(new_n727_));
  OR2_X1    g526(.A1(new_n501_), .A2(G15gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n687_), .B2(new_n728_), .ZN(G1326gat));
  OAI21_X1  g528(.A(G22gat), .B1(new_n712_), .B2(new_n473_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT42), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n473_), .A2(G22gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n687_), .B2(new_n732_), .ZN(G1327gat));
  NAND2_X1  g532(.A1(new_n710_), .A2(new_n706_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n550_), .A2(new_n638_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G29gat), .B1(new_n735_), .B2(new_n485_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n709_), .A2(new_n680_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n667_), .A2(new_n681_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n341_), .A2(new_n481_), .A3(new_n696_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n502_), .B1(new_n740_), .B2(new_n694_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n482_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n738_), .B(new_n739_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n738_), .B1(new_n503_), .B2(new_n739_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n737_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT44), .B(new_n737_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n691_), .A2(G29gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n736_), .B1(new_n750_), .B2(new_n751_), .ZN(G1328gat));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n716_), .A3(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G36gat), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n638_), .A2(new_n734_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n718_), .A2(G36gat), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n755_), .B(new_n756_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT45), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT107), .B1(new_n754_), .B2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(KEYINPUT46), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n761_));
  AOI211_X1 g560(.A(KEYINPUT107), .B(new_n761_), .C1(new_n754_), .C2(new_n758_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1329gat));
  NAND3_X1  g562(.A1(new_n750_), .A2(G43gat), .A3(new_n502_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n735_), .A2(new_n502_), .ZN(new_n765_));
  INV_X1    g564(.A(G43gat), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT47), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n764_), .A2(new_n767_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1330gat));
  AOI21_X1  g571(.A(G50gat), .B1(new_n735_), .B2(new_n703_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n703_), .A2(G50gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n750_), .B2(new_n774_), .ZN(G1331gat));
  NOR2_X1   g574(.A1(new_n708_), .A2(new_n546_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n503_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n682_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(new_n598_), .A3(new_n691_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n707_), .A2(new_n680_), .A3(new_n776_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT108), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n707_), .A2(new_n784_), .A3(new_n680_), .A4(new_n776_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(new_n485_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n781_), .B1(new_n787_), .B2(new_n598_), .ZN(G1332gat));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n716_), .ZN(new_n789_));
  XOR2_X1   g588(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(G64gat), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G64gat), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n716_), .A2(new_n596_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT110), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n791_), .A2(new_n792_), .B1(new_n779_), .B2(new_n794_), .ZN(G1333gat));
  OR3_X1    g594(.A1(new_n779_), .A2(G71gat), .A3(new_n501_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n783_), .A2(new_n502_), .A3(new_n785_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n798_), .A3(G71gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G71gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT111), .B(new_n796_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1334gat));
  NAND2_X1  g604(.A1(new_n703_), .A2(new_n462_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT112), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n780_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n783_), .A2(new_n703_), .A3(new_n785_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(G78gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n809_), .B2(G78gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT113), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n808_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1335gat));
  NAND2_X1  g616(.A1(new_n776_), .A2(new_n710_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n739_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT43), .B1(new_n705_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n818_), .B1(new_n820_), .B2(new_n743_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G85gat), .B1(new_n822_), .B2(new_n433_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n777_), .A2(new_n710_), .A3(new_n706_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n551_), .A3(new_n691_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n826_), .ZN(G1336gat));
  OAI21_X1  g626(.A(G92gat), .B1(new_n822_), .B2(new_n718_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n825_), .A2(new_n552_), .A3(new_n716_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1337gat));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(KEYINPUT51), .ZN(new_n832_));
  OAI21_X1  g631(.A(G99gat), .B1(new_n822_), .B2(new_n501_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n825_), .A2(new_n502_), .A3(new_n573_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(KEYINPUT51), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n835_), .B(new_n836_), .Z(G1338gat));
  INV_X1    g636(.A(new_n818_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n703_), .B(new_n838_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840_));
  OAI21_X1  g639(.A(G106gat), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT115), .B1(new_n821_), .B2(new_n703_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT52), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n840_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n821_), .A2(KEYINPUT115), .A3(new_n703_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .A4(G106gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n825_), .A2(new_n458_), .A3(new_n703_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT53), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n848_), .A2(new_n852_), .A3(new_n849_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1339gat));
  NAND2_X1  g653(.A1(new_n546_), .A2(G113gat), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n620_), .B1(new_n623_), .B2(KEYINPUT12), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n618_), .A2(KEYINPUT71), .A3(new_n588_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n610_), .A4(new_n617_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n622_), .A2(KEYINPUT55), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI221_X1 g662(.A(new_n610_), .B1(new_n612_), .B2(new_n611_), .C1(new_n619_), .C2(new_n621_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n616_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n629_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(KEYINPUT117), .A3(new_n868_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n861_), .A2(new_n862_), .B1(new_n616_), .B2(new_n864_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n867_), .B1(new_n870_), .B2(new_n629_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872_));
  INV_X1    g671(.A(new_n868_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n870_), .B2(new_n873_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n869_), .A2(new_n871_), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n634_), .B2(new_n546_), .ZN(new_n877_));
  AOI211_X1 g676(.A(KEYINPUT116), .B(new_n545_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n856_), .B1(new_n875_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n871_), .A2(new_n874_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n869_), .ZN(new_n882_));
  OAI221_X1 g681(.A(KEYINPUT118), .B1(new_n877_), .B2(new_n878_), .C1(new_n881_), .C2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n526_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n532_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n530_), .A2(new_n885_), .ZN(new_n886_));
  OAI221_X1 g685(.A(new_n541_), .B1(new_n884_), .B2(new_n886_), .C1(new_n539_), .C2(new_n885_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n887_), .A2(new_n540_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n636_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n880_), .A2(new_n883_), .A3(new_n889_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n665_), .A2(KEYINPUT57), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT56), .B1(new_n866_), .B2(new_n628_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n870_), .A2(new_n873_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n634_), .B(new_n888_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n739_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n895_), .A2(new_n896_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n892_), .A2(new_n899_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n902_), .B1(new_n890_), .B2(new_n665_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n710_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n683_), .B2(new_n545_), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n638_), .A2(new_n682_), .A3(KEYINPUT54), .A4(new_n546_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n904_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n691_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n716_), .A2(new_n703_), .A3(new_n911_), .A4(new_n501_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(KEYINPUT121), .A3(new_n914_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n914_), .A2(KEYINPUT121), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(KEYINPUT121), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n910_), .A2(new_n912_), .A3(new_n916_), .A4(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n855_), .B1(new_n915_), .B2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n910_), .A2(new_n546_), .A3(new_n912_), .ZN(new_n920_));
  INV_X1    g719(.A(G113gat), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n920_), .A2(KEYINPUT120), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT120), .B1(new_n920_), .B2(new_n921_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n919_), .A2(new_n922_), .A3(new_n923_), .ZN(G1340gat));
  INV_X1    g723(.A(new_n913_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT122), .B(G120gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n708_), .B2(KEYINPUT60), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n925_), .B(new_n927_), .C1(KEYINPUT60), .C2(new_n926_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n708_), .B1(new_n915_), .B2(new_n918_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n926_), .ZN(G1341gat));
  INV_X1    g729(.A(G127gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n925_), .A2(new_n931_), .A3(new_n680_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n710_), .B1(new_n915_), .B2(new_n918_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n931_), .ZN(G1342gat));
  AOI21_X1  g733(.A(G134gat), .B1(new_n925_), .B2(new_n706_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n915_), .A2(new_n918_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n739_), .A2(G134gat), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT123), .Z(new_n938_));
  AOI21_X1  g737(.A(new_n935_), .B1(new_n936_), .B2(new_n938_), .ZN(G1343gat));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n502_), .B1(new_n904_), .B2(new_n909_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n716_), .A2(new_n473_), .A3(new_n911_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n889_), .ZN(new_n944_));
  OAI22_X1  g743(.A1(new_n881_), .A2(new_n882_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n945_), .B2(new_n856_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n706_), .B1(new_n946_), .B2(new_n883_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n892_), .B(new_n899_), .C1(new_n947_), .C2(new_n902_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n908_), .B1(new_n948_), .B2(new_n710_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n942_), .ZN(new_n950_));
  NOR4_X1   g749(.A1(new_n949_), .A2(KEYINPUT124), .A3(new_n502_), .A4(new_n950_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n546_), .B1(new_n943_), .B2(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(G141gat), .ZN(new_n953_));
  OAI211_X1 g752(.A(new_n390_), .B(new_n546_), .C1(new_n943_), .C2(new_n951_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1344gat));
  OAI21_X1  g754(.A(new_n638_), .B1(new_n943_), .B2(new_n951_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(KEYINPUT125), .B(G148gat), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n956_), .A2(new_n958_), .ZN(new_n959_));
  OAI211_X1 g758(.A(new_n638_), .B(new_n957_), .C1(new_n943_), .C2(new_n951_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(G1345gat));
  OAI21_X1  g760(.A(new_n680_), .B1(new_n943_), .B2(new_n951_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(KEYINPUT61), .B(G155gat), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  INV_X1    g763(.A(new_n963_), .ZN(new_n965_));
  OAI211_X1 g764(.A(new_n680_), .B(new_n965_), .C1(new_n943_), .C2(new_n951_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n964_), .A2(new_n966_), .ZN(G1346gat));
  INV_X1    g766(.A(G162gat), .ZN(new_n968_));
  OAI211_X1 g767(.A(new_n968_), .B(new_n706_), .C1(new_n943_), .C2(new_n951_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n941_), .A2(new_n942_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n970_), .A2(KEYINPUT124), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n941_), .A2(new_n940_), .A3(new_n942_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n819_), .B1(new_n971_), .B2(new_n972_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n969_), .B1(new_n973_), .B2(new_n968_), .ZN(G1347gat));
  NOR4_X1   g773(.A1(new_n718_), .A2(new_n703_), .A3(new_n501_), .A4(new_n691_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n890_), .A2(new_n665_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n976_), .A2(new_n901_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n897_), .A2(new_n898_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n978_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n680_), .B1(new_n977_), .B2(new_n979_), .ZN(new_n980_));
  OAI211_X1 g779(.A(new_n546_), .B(new_n975_), .C1(new_n980_), .C2(new_n908_), .ZN(new_n981_));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n981_), .A2(new_n982_), .ZN(new_n983_));
  NAND4_X1  g782(.A1(new_n910_), .A2(KEYINPUT126), .A3(new_n546_), .A4(new_n975_), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n983_), .A2(G169gat), .A3(new_n984_), .ZN(new_n985_));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n985_), .A2(new_n986_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n910_), .A2(new_n975_), .ZN(new_n988_));
  INV_X1    g787(.A(new_n988_), .ZN(new_n989_));
  NAND3_X1  g788(.A1(new_n989_), .A2(new_n278_), .A3(new_n546_), .ZN(new_n990_));
  NAND4_X1  g789(.A1(new_n983_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n984_), .ZN(new_n991_));
  NAND3_X1  g790(.A1(new_n987_), .A2(new_n990_), .A3(new_n991_), .ZN(G1348gat));
  NOR2_X1   g791(.A1(new_n988_), .A2(new_n708_), .ZN(new_n993_));
  XNOR2_X1  g792(.A(new_n993_), .B(new_n226_), .ZN(G1349gat));
  NOR2_X1   g793(.A1(new_n988_), .A2(new_n710_), .ZN(new_n995_));
  MUX2_X1   g794(.A(G183gat), .B(new_n232_), .S(new_n995_), .Z(G1350gat));
  OAI21_X1  g795(.A(G190gat), .B1(new_n988_), .B2(new_n819_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n706_), .A2(new_n236_), .ZN(new_n998_));
  OAI21_X1  g797(.A(new_n997_), .B1(new_n988_), .B2(new_n998_), .ZN(G1351gat));
  NOR2_X1   g798(.A1(new_n718_), .A2(new_n483_), .ZN(new_n1000_));
  OAI211_X1 g799(.A(new_n501_), .B(new_n1000_), .C1(new_n980_), .C2(new_n908_), .ZN(new_n1001_));
  NOR2_X1   g800(.A1(new_n1001_), .A2(new_n545_), .ZN(new_n1002_));
  XNOR2_X1  g801(.A(new_n1002_), .B(new_n259_), .ZN(G1352gat));
  NOR2_X1   g802(.A1(new_n1001_), .A2(new_n708_), .ZN(new_n1004_));
  NOR2_X1   g803(.A1(new_n1004_), .A2(G204gat), .ZN(new_n1005_));
  NAND2_X1  g804(.A1(new_n262_), .A2(new_n263_), .ZN(new_n1006_));
  AOI21_X1  g805(.A(new_n1005_), .B1(new_n1006_), .B2(new_n1004_), .ZN(G1353gat));
  NOR2_X1   g806(.A1(new_n1001_), .A2(new_n710_), .ZN(new_n1008_));
  OR2_X1    g807(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1009_));
  NOR2_X1   g808(.A1(new_n1008_), .A2(new_n1009_), .ZN(new_n1010_));
  XOR2_X1   g809(.A(KEYINPUT63), .B(G211gat), .Z(new_n1011_));
  AOI21_X1  g810(.A(new_n1010_), .B1(new_n1008_), .B2(new_n1011_), .ZN(G1354gat));
  OAI21_X1  g811(.A(G218gat), .B1(new_n1001_), .B2(new_n819_), .ZN(new_n1013_));
  NAND4_X1  g812(.A1(new_n941_), .A2(new_n249_), .A3(new_n706_), .A4(new_n1000_), .ZN(new_n1014_));
  NAND2_X1  g813(.A1(new_n1013_), .A2(new_n1014_), .ZN(new_n1015_));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1016_));
  NAND2_X1  g815(.A1(new_n1015_), .A2(new_n1016_), .ZN(new_n1017_));
  NAND3_X1  g816(.A1(new_n1013_), .A2(KEYINPUT127), .A3(new_n1014_), .ZN(new_n1018_));
  NAND2_X1  g817(.A1(new_n1017_), .A2(new_n1018_), .ZN(G1355gat));
endmodule


