//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n951_, new_n952_, new_n954_, new_n956_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G230gat), .A2(G233gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT10), .B(G99gat), .Z(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n211_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n214_));
  NAND2_X1  g013(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n214_), .A2(G85gat), .A3(G92gat), .A4(new_n215_), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n208_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT6), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT65), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n219_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(KEYINPUT65), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(KEYINPUT6), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n218_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(KEYINPUT66), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n225_), .A2(new_n226_), .A3(new_n218_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n218_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n217_), .A2(new_n228_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT70), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n224_), .A2(KEYINPUT70), .A3(new_n227_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT7), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT7), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT67), .ZN(new_n241_));
  INV_X1    g040(.A(G99gat), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n239_), .A2(new_n241_), .B1(new_n242_), .B2(new_n207_), .ZN(new_n243_));
  AOI211_X1 g042(.A(G99gat), .B(G106gat), .C1(new_n238_), .C2(KEYINPUT7), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n236_), .A2(new_n237_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n211_), .A2(new_n212_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(KEYINPUT69), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(KEYINPUT69), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT8), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n232_), .A2(new_n228_), .A3(new_n245_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n254_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n234_), .B1(new_n252_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT71), .B(G71gat), .ZN(new_n259_));
  INV_X1    g058(.A(G78gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G57gat), .B(G64gat), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n262_), .A2(KEYINPUT11), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n262_), .B(KEYINPUT11), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n264_), .B1(new_n265_), .B2(new_n261_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n257_), .A2(new_n258_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT8), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n268_), .B1(new_n246_), .B2(new_n250_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n253_), .A2(new_n255_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n266_), .B(new_n233_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT72), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n257_), .A2(new_n266_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n205_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n205_), .B1(new_n257_), .B2(new_n266_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n233_), .B1(new_n270_), .B2(new_n269_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n278_));
  INV_X1    g077(.A(new_n266_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n276_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n275_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT73), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n275_), .A2(new_n285_), .A3(new_n282_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G120gat), .B(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT5), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G176gat), .B(G204gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  XOR2_X1   g089(.A(new_n290_), .B(KEYINPUT74), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n284_), .A2(new_n286_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n290_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n275_), .A2(new_n282_), .A3(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(KEYINPUT13), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT13), .B1(new_n293_), .B2(new_n295_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n203_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n298_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(KEYINPUT75), .A3(new_n296_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G29gat), .B(G36gat), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n302_), .A2(KEYINPUT77), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(KEYINPUT77), .ZN(new_n304_));
  XOR2_X1   g103(.A(G43gat), .B(G50gat), .Z(new_n305_));
  OR3_X1    g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n305_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT15), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT80), .B(G8gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT14), .B1(new_n311_), .B2(new_n202_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G15gat), .B(G22gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G8gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT15), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n310_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G229gat), .A2(G233gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT83), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n308_), .B2(new_n319_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n320_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n308_), .A2(new_n319_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n323_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT84), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n330_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n323_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT84), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n327_), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G141gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G169gat), .B(G197gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n332_), .A2(KEYINPUT85), .A3(new_n337_), .A4(new_n341_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n333_), .A2(new_n334_), .B1(new_n322_), .B2(new_n326_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n340_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT85), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n341_), .B1(new_n343_), .B2(new_n336_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n337_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n299_), .A2(new_n301_), .A3(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G127gat), .B(G155gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT16), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G183gat), .B(G211gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G231gat), .A2(G233gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n356_), .B(KEYINPUT81), .Z(new_n357_));
  AND2_X1   g156(.A1(new_n319_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n319_), .A2(new_n357_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n266_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n279_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n355_), .B1(new_n363_), .B2(KEYINPUT17), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(KEYINPUT82), .A3(new_n362_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n355_), .A2(KEYINPUT17), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n277_), .A2(new_n321_), .A3(new_n310_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n257_), .A2(new_n308_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G232gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT35), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n370_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n375_), .A2(new_n376_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n370_), .A2(new_n371_), .A3(new_n381_), .A4(new_n377_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G190gat), .B(G218gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT78), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G134gat), .B(G162gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT36), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n383_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n387_), .B(KEYINPUT36), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n383_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n380_), .A2(KEYINPUT79), .A3(new_n382_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n390_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G141gat), .A2(G148gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT95), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(KEYINPUT95), .B2(KEYINPUT3), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT2), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G155gat), .A2(G162gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(KEYINPUT1), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n412_), .A2(KEYINPUT94), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT1), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n409_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(KEYINPUT94), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n398_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n418_), .A2(new_n404_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n411_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT28), .B1(new_n421_), .B2(KEYINPUT29), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n406_), .A2(new_n410_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT28), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G22gat), .B(G50gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n422_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G78gat), .B(G106gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n432_), .B(KEYINPUT99), .Z(new_n433_));
  OAI22_X1  g232(.A1(new_n430_), .A2(new_n431_), .B1(KEYINPUT100), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n431_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n433_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n429_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n421_), .A2(KEYINPUT29), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT97), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G211gat), .B(G218gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n442_), .B(KEYINPUT96), .Z(new_n443_));
  XNOR2_X1  g242(.A(G197gat), .B(G204gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT21), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT98), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n442_), .B(KEYINPUT96), .ZN(new_n449_));
  INV_X1    g248(.A(new_n446_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n444_), .A2(new_n445_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n447_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(new_n452_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT98), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n421_), .A2(KEYINPUT97), .A3(KEYINPUT29), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n441_), .A2(new_n453_), .A3(new_n455_), .A4(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(G228gat), .A2(G233gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n454_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(new_n458_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n457_), .A2(new_n458_), .B1(new_n439_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n438_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n461_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n434_), .A3(new_n437_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(G71gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(G15gat), .B(G43gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT92), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n469_), .B(KEYINPUT30), .Z(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT89), .B(KEYINPUT23), .ZN(new_n471_));
  AND2_X1   g270(.A1(G183gat), .A2(G190gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(KEYINPUT23), .B2(new_n473_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT25), .B(G183gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT26), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT87), .B1(new_n477_), .B2(G190gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT26), .B(G190gat), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n476_), .B(new_n478_), .C1(new_n479_), .C2(KEYINPUT87), .ZN(new_n480_));
  INV_X1    g279(.A(G169gat), .ZN(new_n481_));
  INV_X1    g280(.A(G176gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT88), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(G169gat), .B2(G176gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT24), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G169gat), .A2(G176gat), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n483_), .A2(new_n485_), .A3(KEYINPUT24), .A4(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n475_), .A2(new_n480_), .A3(new_n488_), .A4(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n471_), .A2(new_n472_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(KEYINPUT23), .B2(new_n472_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(G183gat), .A2(G190gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n489_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT90), .B(G176gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT22), .B(G169gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI22_X1  g297(.A1(new_n493_), .A2(new_n494_), .B1(new_n498_), .B2(KEYINPUT91), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(KEYINPUT91), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n491_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n470_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n470_), .A2(new_n501_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n467_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n504_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n467_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G127gat), .B(G134gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G113gat), .B(G120gat), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G113gat), .B(G120gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(KEYINPUT93), .A3(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT31), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n521_), .A2(KEYINPUT31), .ZN(new_n524_));
  OAI21_X1  g323(.A(G99gat), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n242_), .A3(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n509_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n505_), .A2(new_n508_), .A3(new_n525_), .A4(new_n527_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n465_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n530_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G226gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT19), .ZN(new_n537_));
  INV_X1    g336(.A(new_n498_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n494_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n538_), .B1(new_n539_), .B2(new_n475_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n472_), .A2(KEYINPUT23), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n472_), .B2(new_n471_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n488_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT102), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n542_), .A2(new_n488_), .A3(KEYINPUT102), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n490_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n479_), .B(KEYINPUT101), .Z(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n549_), .B2(new_n476_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n540_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(new_n459_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT20), .B1(new_n501_), .B2(new_n454_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n537_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G8gat), .B(G36gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT18), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G64gat), .B(G92gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  NAND2_X1  g357(.A1(new_n551_), .A2(new_n459_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT20), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n501_), .B2(new_n454_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n537_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n558_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT103), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT103), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n554_), .A2(new_n566_), .A3(new_n563_), .A4(new_n558_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n554_), .A2(new_n563_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n558_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n565_), .A2(new_n567_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT27), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n455_), .A2(new_n453_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n551_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n562_), .B1(new_n574_), .B2(new_n561_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n552_), .A2(new_n553_), .A3(new_n537_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n569_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n564_), .A2(KEYINPUT27), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n571_), .A2(new_n572_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G1gat), .B(G29gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(G85gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT0), .B(G57gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n581_), .B(new_n582_), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n520_), .A2(new_n421_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n423_), .A2(new_n516_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(KEYINPUT4), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G225gat), .A2(G233gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT105), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT4), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n520_), .A2(new_n421_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT104), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT104), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n520_), .A2(new_n421_), .A3(new_n595_), .A4(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n590_), .A2(new_n591_), .A3(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n585_), .A2(new_n586_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n588_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n591_), .B1(new_n590_), .B2(new_n597_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n584_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT107), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n597_), .A2(new_n589_), .A3(new_n587_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT105), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n606_), .A2(new_n583_), .A3(new_n600_), .A4(new_n598_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n604_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n535_), .B(new_n579_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n465_), .A2(new_n533_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n607_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT106), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n597_), .A2(new_n588_), .A3(new_n587_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n583_), .B1(new_n599_), .B2(new_n589_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AND4_X1   g419(.A1(new_n567_), .A2(new_n565_), .A3(new_n570_), .A4(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n607_), .A2(new_n614_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n607_), .A2(KEYINPUT106), .A3(new_n614_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n617_), .A2(new_n621_), .A3(new_n622_), .A4(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n558_), .A2(KEYINPUT32), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n554_), .A2(new_n563_), .A3(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n575_), .A2(new_n576_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n626_), .B1(new_n627_), .B2(new_n625_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n613_), .B1(new_n624_), .B2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n369_), .B(new_n397_), .C1(new_n612_), .C2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n351_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n610_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n608_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n202_), .B1(new_n633_), .B2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT108), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT86), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n342_), .A2(new_n344_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n335_), .A2(new_n327_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n340_), .B1(new_n642_), .B2(KEYINPUT84), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT85), .B1(new_n643_), .B2(new_n337_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n641_), .B2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n349_), .A2(KEYINPUT86), .A3(new_n344_), .A4(new_n342_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n624_), .A2(new_n630_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n613_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n648_), .B1(new_n651_), .B2(new_n611_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT37), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n392_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n390_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n656_), .B1(KEYINPUT37), .B2(new_n396_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n369_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n652_), .A2(new_n299_), .A3(new_n301_), .A4(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n635_), .A2(G1gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n639_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n660_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(KEYINPUT38), .A3(new_n661_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n638_), .A2(new_n663_), .A3(new_n665_), .ZN(G1324gat));
  INV_X1    g465(.A(new_n579_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n311_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT109), .B1(new_n660_), .B2(new_n668_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n607_), .A2(KEYINPUT106), .A3(new_n614_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT106), .B1(new_n607_), .B2(new_n614_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n607_), .A2(new_n614_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n620_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n673_), .A2(new_n571_), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n629_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n611_), .B1(new_n676_), .B2(new_n613_), .ZN(new_n677_));
  AND4_X1   g476(.A1(new_n299_), .A2(new_n677_), .A3(new_n301_), .A4(new_n647_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n679_));
  INV_X1    g478(.A(new_n668_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n659_), .A4(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n669_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT110), .B(KEYINPUT39), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n351_), .A2(new_n632_), .A3(new_n579_), .ZN(new_n684_));
  INV_X1    g483(.A(G8gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n351_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n632_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n667_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n683_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(G8gat), .A3(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n682_), .A2(new_n686_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT112), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT112), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n682_), .A2(new_n686_), .A3(new_n691_), .A4(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT111), .B(KEYINPUT40), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n693_), .A2(new_n695_), .A3(new_n697_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1325gat));
  INV_X1    g500(.A(G15gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n664_), .A2(new_n702_), .A3(new_n531_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT113), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n702_), .B1(new_n633_), .B2(new_n531_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n707_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n703_), .A2(new_n704_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n705_), .A2(new_n708_), .A3(new_n709_), .A4(new_n710_), .ZN(G1326gat));
  INV_X1    g510(.A(G22gat), .ZN(new_n712_));
  INV_X1    g511(.A(new_n465_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n633_), .B2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT42), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n664_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1327gat));
  NOR2_X1   g516(.A1(new_n397_), .A2(new_n369_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n678_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G29gat), .B1(new_n720_), .B2(new_n636_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n657_), .A2(KEYINPUT114), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n656_), .B(new_n723_), .C1(KEYINPUT37), .C2(new_n396_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n677_), .A2(new_n722_), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT43), .ZN(new_n726_));
  INV_X1    g525(.A(new_n657_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(KEYINPUT43), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n677_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n730_), .A2(KEYINPUT44), .A3(new_n687_), .A4(new_n658_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n687_), .A2(new_n658_), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n725_), .A2(KEYINPUT43), .B1(new_n728_), .B2(new_n677_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n731_), .A2(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n636_), .A2(G29gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n721_), .B1(new_n736_), .B2(new_n737_), .ZN(G1328gat));
  NAND3_X1  g537(.A1(new_n731_), .A2(new_n735_), .A3(new_n667_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G36gat), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n579_), .A2(G36gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n719_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n740_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n740_), .A2(new_n744_), .A3(KEYINPUT46), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1329gat));
  NAND4_X1  g548(.A1(new_n731_), .A2(new_n735_), .A3(G43gat), .A4(new_n531_), .ZN(new_n750_));
  INV_X1    g549(.A(G43gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n751_), .B1(new_n719_), .B2(new_n533_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g553(.A1(new_n719_), .A2(G50gat), .A3(new_n465_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n731_), .A2(new_n735_), .A3(new_n713_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G50gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G50gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1331gat));
  INV_X1    g559(.A(new_n677_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(new_n396_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n299_), .A2(new_n301_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n645_), .A2(new_n369_), .A3(new_n646_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n765_), .A2(G57gat), .A3(new_n636_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n763_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n767_), .A2(new_n350_), .A3(new_n761_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n659_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G57gat), .B1(new_n770_), .B2(new_n636_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n771_), .A2(KEYINPUT116), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(KEYINPUT116), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n766_), .B1(new_n772_), .B2(new_n773_), .ZN(G1332gat));
  OR3_X1    g573(.A1(new_n769_), .A2(G64gat), .A3(new_n579_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n765_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G64gat), .B1(new_n776_), .B2(new_n579_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT48), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(KEYINPUT48), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1333gat));
  OR3_X1    g579(.A1(new_n769_), .A2(G71gat), .A3(new_n533_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G71gat), .B1(new_n776_), .B2(new_n533_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(KEYINPUT49), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(KEYINPUT49), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n783_), .B2(new_n784_), .ZN(G1334gat));
  NAND3_X1  g584(.A1(new_n770_), .A2(new_n260_), .A3(new_n713_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G78gat), .B1(new_n776_), .B2(new_n465_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(KEYINPUT50), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(KEYINPUT50), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n786_), .B1(new_n788_), .B2(new_n789_), .ZN(G1335gat));
  NOR3_X1   g589(.A1(new_n767_), .A2(new_n350_), .A3(new_n369_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n730_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792_), .B2(new_n635_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n768_), .A2(new_n718_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n636_), .A2(new_n209_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(G1336gat));
  NOR3_X1   g595(.A1(new_n792_), .A2(new_n210_), .A3(new_n579_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n210_), .B1(new_n794_), .B2(new_n579_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n798_), .A2(KEYINPUT117), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(KEYINPUT117), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n797_), .B1(new_n799_), .B2(new_n800_), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n792_), .B2(new_n533_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n531_), .A2(new_n206_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n794_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g604(.A1(new_n768_), .A2(new_n207_), .A3(new_n713_), .A4(new_n718_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n791_), .A2(new_n730_), .A3(new_n713_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n807_), .A2(G106gat), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n807_), .B2(G106gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT53), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(new_n806_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1339gat));
  XNOR2_X1  g614(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n764_), .B(new_n656_), .C1(KEYINPUT37), .C2(new_n396_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n300_), .A2(new_n296_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n297_), .A2(new_n298_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n816_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n820_), .A2(new_n727_), .A3(new_n764_), .A4(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n295_), .B1(new_n641_), .B2(new_n644_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n271_), .A2(new_n204_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT12), .B1(new_n257_), .B2(new_n266_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT55), .B1(new_n828_), .B2(KEYINPUT120), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n282_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n280_), .A2(new_n281_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n205_), .B1(new_n833_), .B2(new_n273_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n829_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n292_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(KEYINPUT56), .A3(new_n292_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n824_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n333_), .A2(new_n324_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n322_), .A2(new_n330_), .A3(new_n325_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n341_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n344_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT57), .B(new_n397_), .C1(new_n840_), .C2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n397_), .B1(new_n840_), .B2(new_n845_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n295_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n345_), .B2(new_n349_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n835_), .A2(KEYINPUT56), .A3(new_n292_), .ZN(new_n854_));
  AOI21_X1  g653(.A(KEYINPUT56), .B1(new_n835_), .B2(new_n292_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n293_), .A2(new_n295_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n844_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n860_), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n397_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n852_), .A2(new_n844_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT58), .B(new_n862_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n657_), .A3(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n848_), .A2(new_n851_), .A3(new_n861_), .A4(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n823_), .B1(new_n868_), .B2(new_n658_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n635_), .A2(new_n667_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n532_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n869_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(G113gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n350_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n868_), .A2(new_n658_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n823_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n872_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(KEYINPUT59), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n869_), .B2(new_n872_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n648_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n875_), .B1(new_n883_), .B2(new_n874_), .ZN(G1340gat));
  AOI21_X1  g683(.A(new_n767_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT122), .B(G120gat), .Z(new_n886_));
  NAND2_X1  g685(.A1(new_n878_), .A2(new_n879_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n767_), .B2(KEYINPUT60), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(KEYINPUT60), .B2(new_n886_), .ZN(new_n889_));
  OAI22_X1  g688(.A1(new_n885_), .A2(new_n886_), .B1(new_n887_), .B2(new_n889_), .ZN(G1341gat));
  INV_X1    g689(.A(G127gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n658_), .A2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT59), .B1(new_n878_), .B2(new_n879_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n869_), .A2(new_n881_), .A3(new_n872_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n891_), .B1(new_n887_), .B2(new_n658_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n892_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G127gat), .B1(new_n873_), .B2(new_n369_), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT123), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n898_), .A2(new_n902_), .ZN(G1342gat));
  INV_X1    g702(.A(G134gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n873_), .A2(new_n904_), .A3(new_n396_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n727_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n904_), .ZN(G1343gat));
  NOR2_X1   g706(.A1(new_n869_), .A2(new_n534_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n870_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n350_), .ZN(new_n910_));
  OR3_X1    g709(.A1(new_n909_), .A2(G141gat), .A3(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G141gat), .B1(new_n909_), .B2(new_n910_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1344gat));
  NAND3_X1  g712(.A1(new_n908_), .A2(new_n763_), .A3(new_n870_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT124), .B(G148gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1345gat));
  XNOR2_X1  g715(.A(KEYINPUT61), .B(G155gat), .ZN(new_n917_));
  OR3_X1    g716(.A1(new_n909_), .A2(new_n658_), .A3(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n909_), .B2(new_n658_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1346gat));
  INV_X1    g719(.A(new_n909_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n396_), .ZN(new_n922_));
  INV_X1    g721(.A(G162gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n722_), .A2(G162gat), .A3(new_n724_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(KEYINPUT125), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n922_), .A2(new_n923_), .B1(new_n921_), .B2(new_n925_), .ZN(G1347gat));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n636_), .A2(new_n579_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n531_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT126), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n928_), .A2(new_n931_), .A3(new_n531_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n930_), .A2(new_n465_), .A3(new_n932_), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n869_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n910_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n927_), .B1(new_n935_), .B2(new_n481_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n497_), .ZN(new_n937_));
  OAI211_X1 g736(.A(KEYINPUT62), .B(G169gat), .C1(new_n934_), .C2(new_n910_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(G1348gat));
  NOR2_X1   g738(.A1(new_n869_), .A2(new_n933_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n496_), .B1(new_n940_), .B2(new_n763_), .ZN(new_n941_));
  NOR4_X1   g740(.A1(new_n869_), .A2(G176gat), .A3(new_n767_), .A4(new_n933_), .ZN(new_n942_));
  OAI21_X1  g741(.A(KEYINPUT127), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n940_), .A2(new_n482_), .A3(new_n763_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n869_), .A2(new_n767_), .A3(new_n933_), .ZN(new_n946_));
  OAI211_X1 g745(.A(new_n944_), .B(new_n945_), .C1(new_n496_), .C2(new_n946_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n943_), .A2(new_n947_), .ZN(G1349gat));
  NAND2_X1  g747(.A1(new_n940_), .A2(new_n369_), .ZN(new_n949_));
  MUX2_X1   g748(.A(new_n476_), .B(G183gat), .S(new_n949_), .Z(G1350gat));
  OAI21_X1  g749(.A(G190gat), .B1(new_n934_), .B2(new_n727_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n940_), .A2(new_n396_), .A3(new_n549_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1351gat));
  NAND3_X1  g752(.A1(new_n908_), .A2(new_n350_), .A3(new_n928_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g754(.A1(new_n908_), .A2(new_n763_), .A3(new_n928_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g756(.A1(new_n908_), .A2(new_n369_), .A3(new_n928_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(KEYINPUT63), .B(G211gat), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n960_), .B1(new_n958_), .B2(new_n961_), .ZN(G1354gat));
  INV_X1    g761(.A(G218gat), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n908_), .A2(new_n963_), .A3(new_n396_), .A4(new_n928_), .ZN(new_n964_));
  AND3_X1   g763(.A1(new_n908_), .A2(new_n657_), .A3(new_n928_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n964_), .B1(new_n965_), .B2(new_n963_), .ZN(G1355gat));
endmodule


