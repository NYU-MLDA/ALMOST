//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G57gat), .B(G64gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT11), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(KEYINPUT11), .ZN(new_n209_));
  XOR2_X1   g008(.A(G71gat), .B(G78gat), .Z(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n209_), .A2(new_n210_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(KEYINPUT12), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT66), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  AND3_X1   g023(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  INV_X1    g028(.A(G106gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n227_), .A2(new_n231_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n224_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n224_), .B2(new_n236_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(G85gat), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n220_), .A2(KEYINPUT9), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G99gat), .A2(G106gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT10), .B(G99gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n254_), .B2(new_n230_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n247_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n243_), .A2(new_n244_), .B1(KEYINPUT9), .B2(new_n215_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n227_), .B1(G106gat), .B2(new_n253_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT68), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n214_), .B1(new_n240_), .B2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n258_), .A2(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n234_), .A2(new_n235_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n231_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n217_), .A2(new_n223_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT8), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n224_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n264_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n211_), .A2(new_n212_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n263_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n264_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n272_), .B(new_n274_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G230gat), .A2(G233gat), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n262_), .B(new_n273_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n274_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n272_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT67), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(new_n275_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n271_), .A2(KEYINPUT67), .A3(new_n272_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n277_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n206_), .B1(new_n280_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n280_), .A2(new_n287_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(new_n205_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n280_), .A2(new_n287_), .A3(KEYINPUT72), .A4(new_n206_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT13), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n290_), .A2(KEYINPUT13), .A3(new_n295_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT73), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n299_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G229gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G29gat), .B(G36gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G43gat), .B(G50gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G1gat), .B(G8gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(G15gat), .B(G22gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n321_));
  INV_X1    g120(.A(G1gat), .ZN(new_n322_));
  INV_X1    g121(.A(G8gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT14), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n321_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT82), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT82), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(new_n325_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n319_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n331_), .A3(new_n319_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n318_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n334_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n336_), .A2(new_n317_), .A3(new_n332_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n308_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT15), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n316_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(KEYINPUT15), .A3(new_n314_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n334_), .A3(new_n333_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n317_), .B1(new_n336_), .B2(new_n332_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n307_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n338_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G113gat), .B(G141gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT85), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G169gat), .B(G197gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n338_), .A2(new_n346_), .A3(new_n351_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT86), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358_));
  INV_X1    g157(.A(G43gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT30), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(G15gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n361_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT23), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT92), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n369_), .A2(KEYINPUT92), .A3(new_n371_), .A4(new_n372_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G169gat), .ZN(new_n377_));
  INV_X1    g176(.A(G176gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n379_), .A2(KEYINPUT91), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT89), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(KEYINPUT91), .B2(new_n379_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n375_), .A2(new_n376_), .A3(new_n380_), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n366_), .A2(KEYINPUT23), .ZN(new_n385_));
  INV_X1    g184(.A(new_n368_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n385_), .B1(new_n386_), .B2(KEYINPUT23), .ZN(new_n387_));
  NOR3_X1   g186(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n382_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n388_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G183gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(KEYINPUT87), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT25), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT26), .B(G190gat), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n395_), .A2(KEYINPUT88), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT88), .B1(new_n395_), .B2(new_n396_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n387_), .B(new_n392_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n384_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n365_), .A2(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n361_), .A2(new_n364_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n361_), .A2(new_n364_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n402_), .A2(new_n399_), .A3(new_n384_), .A4(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT93), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n401_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT31), .ZN(new_n407_));
  XOR2_X1   g206(.A(G127gat), .B(G134gat), .Z(new_n408_));
  XOR2_X1   g207(.A(G113gat), .B(G120gat), .Z(new_n409_));
  XOR2_X1   g208(.A(new_n408_), .B(new_n409_), .Z(new_n410_));
  INV_X1    g209(.A(KEYINPUT31), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n401_), .A2(new_n404_), .A3(new_n405_), .A4(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n407_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n410_), .B1(new_n407_), .B2(new_n412_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G85gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT0), .B(G57gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422_));
  OR2_X1    g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT3), .ZN(new_n424_));
  INV_X1    g223(.A(G141gat), .ZN(new_n425_));
  INV_X1    g224(.A(G148gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT2), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT94), .B1(G141gat), .B2(G148gat), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n427_), .B(new_n428_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n430_), .A2(new_n429_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n422_), .B(new_n423_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n422_), .A2(KEYINPUT1), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n422_), .A2(KEYINPUT1), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n423_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G141gat), .A2(G148gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n425_), .A2(new_n426_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n410_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n441_), .A2(KEYINPUT4), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n433_), .A2(new_n439_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n408_), .B(new_n409_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(KEYINPUT4), .A3(new_n441_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G225gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n445_), .B2(new_n441_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n421_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n448_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n454_), .A2(new_n420_), .A3(new_n451_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT18), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G64gat), .B(G92gat), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n458_), .B(new_n459_), .Z(new_n460_));
  NAND2_X1  g259(.A1(G226gat), .A2(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT19), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n464_));
  XOR2_X1   g263(.A(G211gat), .B(G218gat), .Z(new_n465_));
  INV_X1    g264(.A(G197gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(G204gat), .ZN(new_n467_));
  INV_X1    g266(.A(G204gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G197gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(KEYINPUT21), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT96), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT96), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n465_), .A2(new_n473_), .A3(KEYINPUT21), .A4(new_n470_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n470_), .A2(KEYINPUT21), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(new_n465_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT95), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n466_), .A3(G204gat), .ZN(new_n479_));
  OAI211_X1 g278(.A(KEYINPUT21), .B(new_n479_), .C1(new_n470_), .C2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n475_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n464_), .B1(new_n400_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n389_), .A2(new_n379_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n387_), .B2(new_n372_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n475_), .A2(new_n481_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n369_), .A2(new_n371_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n388_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT25), .B(G183gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n396_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n391_), .A2(new_n381_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT98), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n488_), .B(new_n489_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n486_), .A2(new_n487_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n463_), .B1(new_n483_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n384_), .A2(new_n399_), .A3(new_n487_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n369_), .A2(new_n489_), .A3(new_n371_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n496_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n494_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n482_), .B1(new_n503_), .B2(new_n485_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(KEYINPUT20), .A3(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(new_n462_), .ZN(new_n506_));
  OAI211_X1 g305(.A(KEYINPUT32), .B(new_n460_), .C1(new_n499_), .C2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT99), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n498_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n486_), .A2(new_n487_), .A3(KEYINPUT99), .A4(new_n497_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n483_), .A2(new_n463_), .A3(new_n509_), .A4(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n505_), .A2(new_n462_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n460_), .A2(KEYINPUT32), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n456_), .A2(new_n507_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT100), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT33), .B1(new_n453_), .B2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n420_), .B1(new_n454_), .B2(new_n451_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT33), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(KEYINPUT100), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n511_), .A2(new_n512_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n460_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n511_), .A2(new_n512_), .A3(new_n460_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n445_), .A2(new_n449_), .A3(new_n441_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n421_), .B(new_n526_), .C1(new_n447_), .C2(new_n449_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n524_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n515_), .B1(new_n521_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G78gat), .B(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT29), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n482_), .B1(new_n443_), .B2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(G228gat), .A2(G233gat), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n534_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n531_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n536_), .A3(new_n531_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n440_), .A2(KEYINPUT29), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G22gat), .B(G50gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT28), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n541_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT97), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n537_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n540_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n538_), .A2(new_n545_), .A3(new_n539_), .A4(new_n544_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n529_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT27), .B1(new_n524_), .B2(new_n525_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n523_), .B1(new_n499_), .B2(new_n506_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n553_), .A2(KEYINPUT27), .A3(new_n525_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n456_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n416_), .B1(new_n551_), .B2(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n413_), .A2(new_n414_), .A3(new_n456_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT27), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n511_), .A2(new_n512_), .A3(new_n460_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n460_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT101), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n553_), .A2(KEYINPUT27), .A3(new_n525_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n559_), .B(new_n550_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n357_), .B1(new_n558_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT79), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT35), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n572_));
  NAND2_X1  g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n271_), .A2(new_n317_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n240_), .A2(new_n261_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n576_), .A2(KEYINPUT76), .A3(new_n343_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT76), .B1(new_n576_), .B2(new_n343_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n575_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n574_), .A2(new_n571_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT77), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n575_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  OAI221_X1 g382(.A(new_n575_), .B1(new_n581_), .B2(new_n580_), .C1(new_n577_), .C2(new_n578_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT78), .ZN(new_n587_));
  XOR2_X1   g386(.A(G134gat), .B(G162gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n570_), .B1(new_n585_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n583_), .A2(new_n584_), .A3(KEYINPUT79), .A4(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n589_), .B(KEYINPUT36), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n585_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n597_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n585_), .B2(KEYINPUT80), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n583_), .A2(new_n584_), .A3(new_n602_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n592_), .A2(new_n594_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n599_), .B1(new_n604_), .B2(KEYINPUT37), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n333_), .A2(new_n334_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n282_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n282_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT83), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n610_), .B(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G127gat), .B(G155gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(KEYINPUT17), .A3(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n619_), .B(KEYINPUT17), .Z(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n620_), .B1(new_n614_), .B2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n605_), .A2(new_n623_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n306_), .A2(new_n569_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n456_), .B(KEYINPUT102), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627_));
  AOI21_X1  g426(.A(G1gat), .B1(new_n627_), .B2(KEYINPUT103), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n626_), .A3(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n627_), .A2(KEYINPUT103), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n604_), .B1(new_n558_), .B2(new_n568_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n300_), .A2(new_n355_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n623_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT104), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(new_n456_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n631_), .B1(new_n637_), .B2(new_n322_), .ZN(G1324gat));
  NOR2_X1   g437(.A1(new_n566_), .A2(new_n567_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n632_), .A2(new_n634_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G8gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT39), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n625_), .A2(new_n323_), .A3(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g444(.A1(new_n625_), .A2(new_n363_), .A3(new_n415_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n636_), .A2(new_n415_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n647_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT41), .B1(new_n647_), .B2(G15gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n646_), .B1(new_n648_), .B2(new_n649_), .ZN(G1326gat));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n625_), .A2(new_n651_), .A3(new_n549_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n636_), .A2(new_n549_), .ZN(new_n653_));
  XOR2_X1   g452(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(G22gat), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n653_), .B2(G22gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(G1327gat));
  INV_X1    g456(.A(new_n623_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n601_), .A2(new_n603_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n595_), .A2(new_n659_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n302_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n569_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G29gat), .B1(new_n663_), .B2(new_n456_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n633_), .A2(new_n658_), .ZN(new_n665_));
  AOI22_X1  g464(.A1(new_n529_), .A2(new_n550_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n568_), .B1(new_n666_), .B2(new_n415_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n605_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(new_n605_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(KEYINPUT106), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672_));
  AOI211_X1 g471(.A(new_n672_), .B(new_n668_), .C1(new_n667_), .C2(new_n605_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT44), .B(new_n665_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n674_), .A2(G29gat), .A3(new_n626_), .ZN(new_n675_));
  AOI22_X1  g474(.A1(new_n660_), .A2(new_n596_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n558_), .B2(new_n568_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n677_), .B2(new_n668_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n670_), .A2(KEYINPUT106), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n669_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT44), .B1(new_n680_), .B2(new_n665_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n664_), .B1(new_n675_), .B2(new_n682_), .ZN(G1328gat));
  NAND2_X1  g482(.A1(new_n674_), .A2(new_n639_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G36gat), .B1(new_n684_), .B2(new_n681_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n639_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n662_), .A2(G36gat), .A3(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT45), .Z(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n685_), .A2(new_n688_), .A3(KEYINPUT46), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  OAI21_X1  g492(.A(new_n359_), .B1(new_n662_), .B2(new_n416_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n674_), .A2(G43gat), .A3(new_n415_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n681_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g496(.A(G50gat), .B1(new_n663_), .B2(new_n549_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n674_), .A2(G50gat), .A3(new_n549_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n682_), .ZN(G1331gat));
  AOI21_X1  g499(.A(new_n355_), .B1(new_n558_), .B2(new_n568_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n701_), .A2(new_n302_), .A3(new_n624_), .ZN(new_n702_));
  INV_X1    g501(.A(G57gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n626_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n623_), .A2(new_n356_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n305_), .A2(new_n632_), .A3(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(new_n456_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n707_), .B2(new_n703_), .ZN(G1332gat));
  INV_X1    g507(.A(G64gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n702_), .A2(new_n709_), .A3(new_n639_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(new_n639_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G64gat), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n712_), .A2(KEYINPUT108), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(KEYINPUT108), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n715_));
  AND3_X1   g514(.A1(new_n713_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n710_), .B1(new_n716_), .B2(new_n717_), .ZN(G1333gat));
  INV_X1    g517(.A(G71gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n706_), .B2(new_n415_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n702_), .A2(new_n719_), .A3(new_n415_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1334gat));
  INV_X1    g523(.A(G78gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n706_), .B2(new_n549_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT50), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n702_), .A2(new_n725_), .A3(new_n549_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n658_), .A2(new_n660_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n305_), .A2(new_n701_), .A3(new_n730_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT110), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(KEYINPUT110), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n218_), .A3(new_n626_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT111), .B1(new_n671_), .B2(new_n673_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n678_), .A2(new_n679_), .A3(new_n737_), .A4(new_n669_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n355_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n302_), .A2(new_n623_), .A3(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(new_n456_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n735_), .B1(new_n744_), .B2(new_n218_), .ZN(G1336gat));
  AOI21_X1  g544(.A(G92gat), .B1(new_n734_), .B2(new_n639_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n241_), .A2(new_n242_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n686_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n743_), .B2(new_n748_), .ZN(G1337gat));
  XNOR2_X1  g548(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n750_));
  INV_X1    g549(.A(new_n742_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n739_), .A2(new_n415_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G99gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n415_), .A2(new_n254_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n750_), .B1(new_n753_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n750_), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n755_), .B(new_n758_), .C1(new_n752_), .C2(G99gat), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1338gat));
  NAND2_X1  g559(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G106gat), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n742_), .A2(new_n550_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n680_), .B2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n766_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n734_), .A2(new_n230_), .A3(new_n549_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n767_), .A2(new_n772_), .A3(new_n768_), .A4(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  NAND2_X1  g573(.A1(new_n300_), .A2(new_n705_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT54), .B1(new_n775_), .B2(new_n605_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n676_), .A2(new_n777_), .A3(new_n300_), .A4(new_n705_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n295_), .A2(new_n355_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n273_), .A2(new_n262_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n279_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n786_), .B2(KEYINPUT55), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(KEYINPUT55), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n273_), .A2(new_n262_), .A3(new_n275_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n273_), .A2(new_n262_), .A3(KEYINPUT115), .A4(new_n275_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n286_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n280_), .A2(KEYINPUT114), .A3(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n787_), .A2(new_n788_), .A3(new_n793_), .A4(new_n795_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n205_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n205_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n781_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT116), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n781_), .B(new_n801_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n307_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n344_), .A2(new_n345_), .A3(new_n308_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n352_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n354_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n290_), .B2(new_n295_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n800_), .A2(new_n802_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n660_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n604_), .A2(new_n811_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n295_), .A2(new_n355_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n796_), .A2(new_n205_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n205_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n814_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n808_), .B1(new_n819_), .B2(new_n801_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n802_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n813_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI211_X1 g623(.A(KEYINPUT117), .B(new_n806_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  INV_X1    g625(.A(new_n806_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n295_), .B2(new_n827_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n825_), .A2(new_n828_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI221_X1 g630(.A(KEYINPUT58), .B1(new_n797_), .B2(new_n798_), .C1(new_n828_), .C2(new_n825_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n605_), .A3(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n809_), .A2(KEYINPUT118), .A3(new_n813_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n812_), .A2(new_n824_), .A3(new_n833_), .A4(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n780_), .B1(new_n835_), .B2(new_n623_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n626_), .ZN(new_n837_));
  NOR4_X1   g636(.A1(new_n639_), .A2(new_n837_), .A3(new_n549_), .A4(new_n416_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(G113gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n355_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(KEYINPUT59), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n357_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n842_), .B1(new_n846_), .B2(new_n841_), .ZN(G1340gat));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n300_), .B2(KEYINPUT60), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n840_), .B(new_n849_), .C1(KEYINPUT60), .C2(new_n848_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n306_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n848_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n840_), .B2(new_n658_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n843_), .A2(new_n845_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(G127gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n658_), .A2(KEYINPUT119), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(G127gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n853_), .B1(new_n854_), .B2(new_n858_), .ZN(G1342gat));
  AOI21_X1  g658(.A(new_n807_), .B1(new_n799_), .B2(KEYINPUT116), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n604_), .B1(new_n860_), .B2(new_n802_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n833_), .B1(new_n861_), .B2(KEYINPUT57), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n809_), .A2(KEYINPUT118), .A3(new_n813_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT118), .B1(new_n809_), .B2(new_n813_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n779_), .B1(new_n865_), .B2(new_n658_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n604_), .A3(new_n838_), .ZN(new_n867_));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(KEYINPUT120), .A3(new_n868_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n676_), .A2(new_n868_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n871_), .A2(new_n872_), .B1(new_n854_), .B2(new_n873_), .ZN(G1343gat));
  XNOR2_X1  g673(.A(KEYINPUT121), .B(G141gat), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877_));
  NOR4_X1   g676(.A1(new_n639_), .A2(new_n837_), .A3(new_n550_), .A4(new_n415_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n836_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n877_), .B1(new_n880_), .B2(new_n355_), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n836_), .A2(KEYINPUT122), .A3(new_n741_), .A4(new_n879_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n876_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n866_), .A2(new_n355_), .A3(new_n878_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT122), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n880_), .A2(new_n877_), .A3(new_n355_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n875_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n887_), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n880_), .A2(new_n305_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g689(.A1(new_n863_), .A2(new_n864_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n862_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n658_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n658_), .B(new_n878_), .C1(new_n893_), .C2(new_n780_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT123), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n866_), .A2(new_n896_), .A3(new_n658_), .A4(new_n878_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT61), .B(G155gat), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n895_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1346gat));
  INV_X1    g700(.A(G162gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n880_), .A2(new_n902_), .A3(new_n604_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n836_), .A2(new_n676_), .A3(new_n879_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n902_), .B2(new_n904_), .ZN(G1347gat));
  INV_X1    g704(.A(G169gat), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(KEYINPUT62), .ZN(new_n908_));
  NOR4_X1   g707(.A1(new_n686_), .A2(new_n549_), .A3(new_n416_), .A4(new_n626_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n866_), .A2(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n910_), .B2(new_n741_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(KEYINPUT124), .A3(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n909_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n836_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n915_), .A2(new_n377_), .A3(new_n355_), .ZN(new_n916_));
  OAI221_X1 g715(.A(new_n908_), .B1(new_n907_), .B2(KEYINPUT62), .C1(new_n910_), .C2(new_n741_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n913_), .A2(new_n916_), .A3(new_n917_), .ZN(G1348gat));
  OAI21_X1  g717(.A(G176gat), .B1(new_n910_), .B2(new_n306_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n915_), .A2(new_n378_), .A3(new_n302_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1349gat));
  NAND2_X1  g720(.A1(new_n915_), .A2(new_n658_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n490_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n393_), .B2(new_n922_), .ZN(G1350gat));
  OAI21_X1  g723(.A(G190gat), .B1(new_n910_), .B2(new_n676_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n915_), .A2(new_n396_), .A3(new_n604_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1351gat));
  NAND2_X1  g726(.A1(new_n416_), .A2(new_n556_), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT125), .Z(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(new_n686_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT126), .B1(new_n836_), .B2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n933_), .B(new_n930_), .C1(new_n893_), .C2(new_n780_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935_), .B2(new_n355_), .ZN(new_n936_));
  AOI211_X1 g735(.A(new_n466_), .B(new_n741_), .C1(new_n932_), .C2(new_n934_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1352gat));
  AOI21_X1  g737(.A(new_n933_), .B1(new_n866_), .B2(new_n930_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n836_), .A2(KEYINPUT126), .A3(new_n931_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n305_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(G204gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n935_), .A2(new_n468_), .A3(new_n305_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1353gat));
  OR2_X1    g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n945_), .B1(new_n935_), .B2(new_n658_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(KEYINPUT63), .B(G211gat), .ZN(new_n947_));
  AOI211_X1 g746(.A(new_n623_), .B(new_n947_), .C1(new_n932_), .C2(new_n934_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n946_), .A2(new_n948_), .ZN(G1354gat));
  NAND2_X1  g748(.A1(new_n935_), .A2(new_n604_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT127), .B(G218gat), .Z(new_n951_));
  NOR2_X1   g750(.A1(new_n676_), .A2(new_n951_), .ZN(new_n952_));
  AOI22_X1  g751(.A1(new_n950_), .A2(new_n951_), .B1(new_n935_), .B2(new_n952_), .ZN(G1355gat));
endmodule


