//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  NOR3_X1   g005(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(G169gat), .B2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n207_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT25), .B(G183gat), .Z(new_n214_));
  INV_X1    g013(.A(KEYINPUT78), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT79), .B(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n216_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G183gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n215_), .B1(KEYINPUT25), .B2(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n206_), .B(new_n213_), .C1(new_n221_), .C2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n210_), .A2(new_n211_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(new_n226_), .B2(new_n211_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT80), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT80), .B1(new_n202_), .B2(KEYINPUT23), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n217_), .A2(new_n222_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n227_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n224_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT30), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237_));
  INV_X1    g036(.A(G113gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G120gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n236_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G15gat), .B(G43gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  NOR2_X1   g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n241_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n236_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n245_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G71gat), .B(G99gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OR3_X1    g053(.A1(new_n246_), .A2(new_n250_), .A3(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n246_), .B2(new_n250_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT83), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(G155gat), .B2(G162gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT83), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT1), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G155gat), .ZN(new_n263_));
  INV_X1    g062(.A(G162gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT82), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT82), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(G155gat), .B2(G162gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n260_), .A2(KEYINPUT83), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n258_), .A2(G155gat), .A3(G162gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n262_), .A2(new_n265_), .A3(new_n267_), .A4(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G141gat), .ZN(new_n273_));
  INV_X1    g072(.A(G148gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT85), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n280_), .A2(new_n282_), .A3(new_n283_), .A4(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT84), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n290_), .A2(KEYINPUT84), .A3(new_n283_), .A4(new_n280_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n265_), .B(new_n267_), .C1(new_n259_), .C2(new_n261_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n278_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  AOI211_X1 g094(.A(KEYINPUT85), .B(new_n293_), .C1(new_n287_), .C2(new_n291_), .ZN(new_n296_));
  OAI211_X1 g095(.A(KEYINPUT93), .B(new_n277_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n247_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n283_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT84), .B1(new_n301_), .B2(new_n290_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n285_), .A2(new_n286_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n294_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT85), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n292_), .A2(new_n278_), .A3(new_n294_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n307_), .A2(KEYINPUT93), .A3(new_n277_), .A4(new_n241_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n298_), .A2(new_n308_), .A3(KEYINPUT4), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n277_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT4), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n247_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n298_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT95), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n298_), .A2(new_n308_), .A3(KEYINPUT95), .A4(new_n310_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G1gat), .B(G29gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G57gat), .B(G85gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n320_), .A2(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n315_), .A2(new_n318_), .A3(new_n325_), .A4(new_n319_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n257_), .A2(new_n329_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n272_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n334_), .A2(KEYINPUT28), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(KEYINPUT28), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G78gat), .B(G106gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(KEYINPUT90), .Z(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n335_), .A2(new_n341_), .A3(new_n336_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G197gat), .B(G204gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT88), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT21), .ZN(new_n346_));
  OR3_X1    g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G211gat), .B(G218gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n346_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  OR4_X1    g149(.A1(new_n345_), .A2(new_n348_), .A3(new_n344_), .A4(new_n346_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n312_), .B2(KEYINPUT29), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n354_));
  INV_X1    g153(.A(G228gat), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n353_), .A2(KEYINPUT89), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT87), .B(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n350_), .A2(new_n351_), .ZN(new_n361_));
  OAI211_X1 g160(.A(KEYINPUT89), .B(new_n361_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n354_), .A2(new_n355_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n362_), .A2(new_n357_), .A3(new_n358_), .A4(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n359_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n353_), .A2(KEYINPUT89), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n360_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n360_), .B2(new_n366_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n343_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n364_), .A2(new_n365_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n364_), .A2(new_n365_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n367_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n342_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n341_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n360_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n374_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n371_), .A2(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(KEYINPUT26), .B(G190gat), .Z(new_n381_));
  OAI221_X1 g180(.A(new_n213_), .B1(new_n214_), .B2(new_n381_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n206_), .B1(G183gat), .B2(G190gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n227_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n361_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n386_), .B(KEYINPUT20), .C1(new_n234_), .C2(new_n361_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n388_), .B(KEYINPUT91), .Z(new_n389_));
  XOR2_X1   g188(.A(new_n389_), .B(KEYINPUT19), .Z(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n234_), .A2(new_n361_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n352_), .A2(new_n384_), .A3(new_n382_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT20), .A4(new_n390_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(G64gat), .B(G92gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n396_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n392_), .A2(new_n401_), .A3(new_n395_), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT27), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n404_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT96), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n352_), .A2(new_n224_), .A3(new_n233_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n408_), .A2(new_n386_), .A3(KEYINPUT20), .A4(new_n390_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT20), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n407_), .B(new_n409_), .C1(new_n410_), .C2(new_n390_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n409_), .A2(new_n407_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n406_), .B1(new_n413_), .B2(new_n402_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n405_), .B1(new_n414_), .B2(KEYINPUT27), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n380_), .A2(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n330_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT97), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n328_), .B(KEYINPUT33), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n403_), .A2(new_n404_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n309_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n298_), .A2(new_n308_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n325_), .B1(new_n422_), .B2(new_n311_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n401_), .A2(KEYINPUT32), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n396_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n413_), .A2(new_n425_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n419_), .A2(new_n424_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n369_), .A2(new_n370_), .A3(new_n343_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n377_), .B1(new_n374_), .B2(new_n378_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n418_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n329_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n434_), .A3(new_n415_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n426_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n329_), .A2(new_n428_), .A3(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n318_), .A2(new_n319_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n438_), .A2(KEYINPUT33), .A3(new_n325_), .A4(new_n315_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n328_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n424_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT97), .A3(new_n380_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n433_), .A2(new_n435_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n417_), .B1(new_n445_), .B2(new_n257_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT7), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G99gat), .A2(G106gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n449_), .A2(new_n452_), .A3(new_n453_), .A4(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G85gat), .B(G92gat), .Z(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT65), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n455_), .A2(KEYINPUT65), .A3(new_n456_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT8), .A3(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT10), .B(G99gat), .Z(new_n462_));
  INV_X1    g261(.A(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n456_), .A2(KEYINPUT9), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT9), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(G85gat), .A3(G92gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n452_), .A2(new_n453_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .A4(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT8), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n457_), .A2(new_n458_), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n461_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G57gat), .B(G64gat), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n474_), .A2(KEYINPUT11), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(KEYINPUT11), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G71gat), .B(G78gat), .ZN(new_n477_));
  OR3_X1    g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n477_), .A3(KEYINPUT11), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n473_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n480_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n472_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G230gat), .A2(G233gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n485_), .B(KEYINPUT64), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT66), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT67), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n490_), .B1(new_n483_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n483_), .A2(new_n491_), .A3(new_n490_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n493_), .A2(new_n486_), .A3(new_n481_), .A4(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT66), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n484_), .A2(new_n496_), .A3(new_n487_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n489_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G120gat), .B(G148gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(G204gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT5), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(new_n211_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT13), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n489_), .A2(new_n495_), .A3(new_n497_), .A4(new_n502_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n505_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G29gat), .B(G36gat), .ZN(new_n511_));
  INV_X1    g310(.A(G43gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(G50gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516_));
  INV_X1    g315(.A(G1gat), .ZN(new_n517_));
  INV_X1    g316(.A(G8gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G1gat), .B(G8gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n515_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n513_), .B(G50gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n526_), .A2(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n515_), .A2(KEYINPUT15), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n531_), .B2(new_n522_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n525_), .B1(new_n524_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G113gat), .B(G141gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(new_n210_), .ZN(new_n535_));
  INV_X1    g334(.A(G197gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT76), .ZN(new_n538_));
  OR3_X1    g337(.A1(new_n533_), .A2(KEYINPUT77), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT77), .B1(new_n533_), .B2(new_n538_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n539_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n510_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT74), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n522_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n480_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G127gat), .B(G155gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G183gat), .B(G211gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n555_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n549_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n557_), .B2(new_n549_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n545_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n446_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n531_), .A2(new_n472_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n473_), .A2(new_n515_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT34), .Z(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT68), .B(KEYINPUT35), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(new_n565_), .A3(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n567_), .A2(new_n568_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n564_), .A2(new_n565_), .A3(new_n573_), .A4(new_n569_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT72), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT69), .B(G190gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT36), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT71), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT72), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n572_), .A2(new_n584_), .A3(new_n574_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n576_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  INV_X1    g386(.A(new_n580_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n572_), .A2(new_n589_), .A3(new_n574_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT73), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n582_), .B1(new_n575_), .B2(KEYINPUT72), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n590_), .B1(new_n594_), .B2(new_n585_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT73), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(new_n587_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT70), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n572_), .A2(new_n599_), .A3(new_n589_), .A4(new_n574_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT37), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n590_), .B1(new_n575_), .B2(new_n583_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n602_), .B2(KEYINPUT70), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n563_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT98), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n563_), .A2(new_n608_), .A3(new_n605_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n607_), .A2(new_n517_), .A3(new_n329_), .A4(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n611_));
  OR3_X1    g410(.A1(new_n610_), .A2(KEYINPUT100), .A3(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n562_), .A2(KEYINPUT101), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n446_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n595_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n562_), .A2(KEYINPUT101), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n517_), .B1(new_n617_), .B2(new_n329_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT100), .B1(new_n610_), .B2(new_n611_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n612_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n612_), .A2(new_n619_), .A3(KEYINPUT102), .A4(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1324gat));
  XNOR2_X1  g424(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT104), .ZN(new_n627_));
  INV_X1    g426(.A(new_n415_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n617_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(G8gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT39), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n607_), .A2(new_n518_), .A3(new_n628_), .A4(new_n609_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n627_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n630_), .A2(KEYINPUT39), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n629_), .B2(G8gat), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n632_), .B(new_n627_), .C1(new_n634_), .C2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n633_), .A2(new_n638_), .ZN(G1325gat));
  INV_X1    g438(.A(new_n617_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G15gat), .B1(new_n640_), .B2(new_n257_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT41), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n607_), .A2(new_n609_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n643_), .A2(G15gat), .A3(new_n257_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1326gat));
  OAI21_X1  g444(.A(G22gat), .B1(new_n640_), .B2(new_n380_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT42), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n380_), .A2(G22gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n643_), .B2(new_n648_), .ZN(G1327gat));
  NOR2_X1   g448(.A1(new_n446_), .A2(new_n615_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n545_), .A2(new_n560_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n329_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n652_), .B(KEYINPUT105), .Z(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  INV_X1    g455(.A(new_n417_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n443_), .A2(KEYINPUT97), .A3(new_n380_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT97), .B1(new_n443_), .B2(new_n380_), .ZN(new_n659_));
  AND4_X1   g458(.A1(new_n434_), .A2(new_n415_), .A3(new_n379_), .A4(new_n371_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n257_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n657_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n603_), .B1(new_n593_), .B2(new_n597_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n656_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n446_), .A2(KEYINPUT43), .A3(new_n605_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n655_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n663_), .A2(new_n656_), .A3(new_n664_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT43), .B1(new_n446_), .B2(new_n605_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n655_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n669_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n434_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n654_), .B1(new_n675_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g475(.A1(new_n669_), .A2(new_n628_), .A3(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n653_), .A2(KEYINPUT45), .A3(new_n679_), .A4(new_n628_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT45), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n650_), .A2(new_n679_), .A3(new_n545_), .A4(new_n560_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n415_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n680_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n678_), .A2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT46), .B1(new_n685_), .B2(KEYINPUT106), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n687_), .B(new_n688_), .C1(new_n678_), .C2(new_n684_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n686_), .A2(new_n689_), .ZN(G1329gat));
  NAND3_X1  g489(.A1(new_n669_), .A2(new_n662_), .A3(new_n673_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n257_), .A2(G43gat), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n691_), .A2(G43gat), .B1(new_n653_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g493(.A1(new_n380_), .A2(new_n514_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n651_), .A2(new_n380_), .A3(new_n652_), .ZN(new_n697_));
  OAI22_X1  g496(.A1(new_n674_), .A2(new_n696_), .B1(G50gat), .B2(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT107), .Z(G1331gat));
  INV_X1    g498(.A(new_n509_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n507_), .ZN(new_n701_));
  NOR4_X1   g500(.A1(new_n446_), .A2(new_n701_), .A3(new_n543_), .A4(new_n560_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n605_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n329_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n615_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(new_n434_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(G57gat), .B2(new_n707_), .ZN(G1332gat));
  OAI21_X1  g507(.A(G64gat), .B1(new_n706_), .B2(new_n415_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT48), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n415_), .A2(G64gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n703_), .B2(new_n711_), .ZN(G1333gat));
  OAI21_X1  g511(.A(G71gat), .B1(new_n706_), .B2(new_n257_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT109), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n713_), .B(new_n715_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n257_), .A2(G71gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n703_), .B2(new_n717_), .ZN(G1334gat));
  OAI21_X1  g517(.A(G78gat), .B1(new_n706_), .B2(new_n380_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n380_), .A2(G78gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n703_), .B2(new_n721_), .ZN(G1335gat));
  NAND3_X1  g521(.A1(new_n510_), .A2(new_n544_), .A3(new_n560_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n651_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n329_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n672_), .A2(KEYINPUT110), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n670_), .A2(new_n727_), .A3(new_n671_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n723_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(new_n329_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n725_), .B1(new_n730_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g530(.A(G92gat), .B1(new_n724_), .B2(new_n628_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n729_), .A2(new_n628_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G92gat), .ZN(G1337gat));
  INV_X1    g533(.A(G99gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n729_), .B2(new_n662_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n724_), .A2(new_n462_), .A3(new_n662_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OR3_X1    g539(.A1(new_n736_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n738_), .B1(new_n736_), .B2(new_n740_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1338gat));
  NAND3_X1  g542(.A1(new_n724_), .A2(new_n463_), .A3(new_n432_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n723_), .A2(new_n380_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n672_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n747_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT112), .B(new_n749_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n745_), .B1(new_n751_), .B2(G106gat), .ZN(new_n752_));
  NOR4_X1   g551(.A1(new_n748_), .A2(new_n750_), .A3(KEYINPUT52), .A4(new_n463_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n744_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n744_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1339gat));
  NAND3_X1  g557(.A1(new_n416_), .A2(new_n329_), .A3(new_n662_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n543_), .A2(new_n560_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n701_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n701_), .A2(KEYINPUT113), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n761_), .B1(new_n767_), .B2(new_n605_), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT114), .B(new_n664_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n760_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n766_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT113), .B1(new_n701_), .B2(new_n762_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n605_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT114), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n767_), .A2(new_n761_), .A3(new_n605_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(KEYINPUT54), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n770_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT118), .ZN(new_n778_));
  INV_X1    g577(.A(new_n495_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n493_), .A2(new_n481_), .A3(new_n494_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n487_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n781_), .B2(KEYINPUT55), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n780_), .A2(new_n783_), .A3(new_n487_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n503_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT56), .B(new_n503_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n524_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n532_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n537_), .C1(new_n790_), .C2(new_n523_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n541_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n506_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n789_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(KEYINPUT117), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n794_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT58), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n798_), .A2(new_n664_), .A3(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n541_), .A2(new_n792_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n781_), .A2(KEYINPUT55), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n495_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n784_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n502_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  XOR2_X1   g608(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n810_));
  OAI21_X1  g609(.A(new_n788_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n543_), .A2(new_n506_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n805_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n803_), .B1(new_n814_), .B2(new_n595_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n803_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n810_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n785_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n812_), .B1(new_n818_), .B2(new_n788_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n615_), .B(new_n816_), .C1(new_n819_), .C2(new_n805_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n778_), .B1(new_n802_), .B2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n798_), .A2(new_n664_), .A3(new_n801_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n823_), .A2(KEYINPUT118), .A3(new_n820_), .A4(new_n815_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n560_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n759_), .B1(new_n777_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G113gat), .B1(new_n826_), .B2(new_n543_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n560_), .B1(new_n802_), .B2(new_n821_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n774_), .A2(new_n775_), .A3(KEYINPUT54), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT54), .B1(new_n774_), .B2(new_n775_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n759_), .A2(KEYINPUT59), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n543_), .B(new_n833_), .C1(new_n826_), .C2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n827_), .B1(new_n836_), .B2(G113gat), .ZN(G1340gat));
  OAI211_X1 g636(.A(new_n510_), .B(new_n833_), .C1(new_n826_), .C2(new_n834_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n839_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(G120gat), .A3(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n240_), .B1(new_n701_), .B2(KEYINPUT60), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n826_), .B(new_n843_), .C1(KEYINPUT60), .C2(new_n240_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1341gat));
  OAI211_X1 g644(.A(new_n561_), .B(new_n833_), .C1(new_n826_), .C2(new_n834_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G127gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n777_), .A2(new_n825_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n759_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OR3_X1    g649(.A1(new_n850_), .A2(G127gat), .A3(new_n560_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT120), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n847_), .A2(new_n851_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1342gat));
  INV_X1    g655(.A(G134gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n850_), .B2(new_n615_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT121), .B(G134gat), .Z(new_n859_));
  OAI211_X1 g658(.A(new_n833_), .B(new_n859_), .C1(new_n826_), .C2(new_n834_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n860_), .B2(new_n605_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n858_), .B(KEYINPUT122), .C1(new_n860_), .C2(new_n605_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1343gat));
  AOI211_X1 g664(.A(new_n380_), .B(new_n628_), .C1(new_n777_), .C2(new_n825_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n662_), .A2(new_n434_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n544_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n273_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n701_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n274_), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n868_), .A2(new_n560_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT123), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n873_), .B(new_n875_), .ZN(G1346gat));
  NOR3_X1   g675(.A1(new_n868_), .A2(new_n264_), .A3(new_n605_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n866_), .A2(new_n595_), .A3(new_n867_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n264_), .B2(new_n878_), .ZN(G1347gat));
  NAND2_X1  g678(.A1(new_n330_), .A2(new_n628_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n777_), .B2(new_n828_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n380_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G169gat), .B1(new_n882_), .B2(new_n544_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n882_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n226_), .A3(new_n543_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n884_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n885_), .A2(new_n887_), .A3(new_n888_), .ZN(G1348gat));
  OAI21_X1  g688(.A(new_n211_), .B1(new_n882_), .B2(new_n701_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n432_), .B1(new_n777_), .B2(new_n825_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n880_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n891_), .A2(G176gat), .A3(new_n510_), .A4(new_n892_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n890_), .A2(new_n893_), .ZN(G1349gat));
  AND2_X1   g693(.A1(new_n561_), .A2(new_n214_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n561_), .A3(new_n892_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n886_), .A2(new_n895_), .B1(new_n896_), .B2(new_n222_), .ZN(G1350gat));
  INV_X1    g696(.A(new_n381_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n881_), .A2(new_n595_), .A3(new_n380_), .A4(new_n898_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n831_), .A2(new_n664_), .A3(new_n380_), .A4(new_n892_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n900_), .A2(new_n901_), .A3(G190gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n900_), .B2(G190gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n899_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT125), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n906_), .B(new_n899_), .C1(new_n902_), .C2(new_n903_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1351gat));
  AOI21_X1  g707(.A(new_n329_), .B1(new_n777_), .B2(new_n825_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n662_), .A2(new_n380_), .A3(new_n415_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n544_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n536_), .ZN(G1352gat));
  INV_X1    g712(.A(new_n911_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n510_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g715(.A1(new_n911_), .A2(new_n560_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT126), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT127), .ZN(new_n922_));
  OR2_X1    g721(.A1(new_n921_), .A2(KEYINPUT127), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n919_), .A2(new_n922_), .A3(new_n923_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n917_), .A2(KEYINPUT127), .A3(new_n921_), .A4(new_n918_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1354gat));
  AOI21_X1  g725(.A(G218gat), .B1(new_n914_), .B2(new_n595_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n914_), .A2(G218gat), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n664_), .B2(new_n928_), .ZN(G1355gat));
endmodule


