//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n593_, new_n594_,
    new_n595_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_;
  NOR2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(G155gat), .ZN(new_n205_));
  INV_X1    g004(.A(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT89), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n209_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT90), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n203_), .B(new_n204_), .C1(new_n211_), .C2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n208_), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n202_), .B(KEYINPUT3), .Z(new_n216_));
  XOR2_X1   g015(.A(new_n204_), .B(KEYINPUT2), .Z(new_n217_));
  OAI211_X1 g016(.A(new_n215_), .B(new_n207_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G113gat), .B(G120gat), .Z(new_n220_));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n219_), .B(new_n222_), .Z(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT4), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G225gat), .A2(G233gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n219_), .A2(new_n222_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n224_), .B(new_n226_), .C1(KEYINPUT4), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n225_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G1gat), .B(G29gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G85gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT0), .B(G57gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n232_), .B(new_n233_), .Z(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n228_), .A2(new_n229_), .A3(new_n234_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT20), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT23), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(G183gat), .A3(G190gat), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n242_), .A2(KEYINPUT85), .ZN(new_n243_));
  INV_X1    g042(.A(G183gat), .ZN(new_n244_));
  INV_X1    g043(.A(G190gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT23), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(KEYINPUT85), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(G183gat), .B2(G190gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT96), .ZN(new_n250_));
  INV_X1    g049(.A(G169gat), .ZN(new_n251_));
  INV_X1    g050(.A(G176gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT22), .B(G169gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n254_), .B2(new_n252_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT94), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT25), .B(G183gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n246_), .A2(new_n242_), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT95), .B(KEYINPUT24), .Z(new_n262_));
  INV_X1    g061(.A(new_n253_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n251_), .A2(new_n252_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n262_), .A2(new_n264_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n260_), .A2(new_n261_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n256_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G197gat), .B(G204gat), .Z(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT21), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT92), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n269_), .A2(KEYINPUT21), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n271_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n240_), .B1(new_n268_), .B2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n248_), .B1(KEYINPUT24), .B2(new_n264_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT86), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n263_), .A2(KEYINPUT24), .A3(new_n264_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n281_));
  OR3_X1    g080(.A1(new_n281_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT84), .B1(new_n281_), .B2(G190gat), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n284_), .B(new_n259_), .C1(KEYINPUT26), .C2(new_n245_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n279_), .A2(new_n280_), .A3(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n261_), .B1(G183gat), .B2(G190gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n255_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n277_), .B1(new_n289_), .B2(new_n276_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT19), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n292_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n268_), .A2(new_n276_), .ZN(new_n295_));
  AOI211_X1 g094(.A(new_n240_), .B(new_n295_), .C1(new_n289_), .C2(new_n276_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n293_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G8gat), .B(G36gat), .ZN(new_n298_));
  INV_X1    g097(.A(G92gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT18), .B(G64gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT32), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n239_), .B1(new_n297_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n296_), .A2(new_n294_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n290_), .A2(new_n292_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(new_n304_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT97), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n308_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(new_n302_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n224_), .B(new_n225_), .C1(KEYINPUT4), .C2(new_n227_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n223_), .A2(new_n226_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n313_), .A2(new_n235_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n303_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n312_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n237_), .B(KEYINPUT33), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n306_), .A2(new_n310_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G227gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n222_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n289_), .B(KEYINPUT87), .Z(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT30), .B(G99gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n289_), .B(KEYINPUT87), .ZN(new_n326_));
  INV_X1    g125(.A(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G15gat), .B(G43gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT31), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G71gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n325_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n322_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n335_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(new_n321_), .A3(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT88), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n336_), .A2(new_n338_), .A3(KEYINPUT88), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT93), .ZN(new_n344_));
  INV_X1    g143(.A(new_n219_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT28), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G22gat), .B(G50gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n350_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n344_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n276_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n355_));
  AND2_X1   g154(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(G228gat), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n355_), .B(new_n358_), .Z(new_n359_));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n354_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n351_), .A2(new_n352_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n359_), .A2(new_n360_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n364_), .B2(new_n353_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n366_), .B2(new_n361_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n319_), .A2(new_n343_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n343_), .A2(new_n368_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n312_), .B1(new_n302_), .B2(new_n297_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT27), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT27), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n312_), .B2(new_n316_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n367_), .A2(new_n339_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n371_), .A2(new_n377_), .A3(new_n239_), .A4(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n370_), .A2(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(G43gat), .B(G50gat), .Z(new_n381_));
  XNOR2_X1  g180(.A(G29gat), .B(G36gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT15), .Z(new_n384_));
  NAND2_X1  g183(.A1(G99gat), .A2(G106gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT6), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT10), .B(G99gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT64), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n387_), .B(new_n388_), .C1(new_n391_), .C2(G106gat), .ZN(new_n392_));
  OR2_X1    g191(.A1(G85gat), .A2(G92gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(G92gat), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT66), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT9), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n396_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT67), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n299_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT66), .B1(new_n409_), .B2(KEYINPUT9), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(KEYINPUT67), .A3(new_n396_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n392_), .B1(new_n406_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G85gat), .A2(G92gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT7), .ZN(new_n416_));
  INV_X1    g215(.A(G99gat), .ZN(new_n417_));
  INV_X1    g216(.A(G106gat), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .A4(KEYINPUT68), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT68), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n420_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n387_), .A2(new_n388_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n393_), .B(new_n415_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(KEYINPUT69), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(KEYINPUT69), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT8), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT8), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(KEYINPUT69), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n425_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n384_), .B1(new_n414_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT73), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G232gat), .A2(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT34), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT75), .B1(new_n434_), .B2(KEYINPUT35), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n414_), .A2(new_n430_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n383_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n432_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(KEYINPUT35), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G190gat), .B(G218gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(new_n206_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT74), .B(G134gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n445_), .B(KEYINPUT36), .Z(new_n446_));
  OR2_X1    g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n441_), .B1(KEYINPUT36), .B2(new_n445_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT76), .B(KEYINPUT37), .Z(new_n450_));
  OR2_X1    g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n450_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G127gat), .B(G155gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(G211gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT16), .B(G183gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G15gat), .B(G22gat), .Z(new_n458_));
  NAND2_X1  g257(.A1(G1gat), .A2(G8gat), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(KEYINPUT14), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT77), .ZN(new_n461_));
  XOR2_X1   g260(.A(G1gat), .B(G8gat), .Z(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT77), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n460_), .B(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n462_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G231gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT78), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n468_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G57gat), .B(G64gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT11), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G71gat), .B(G78gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n473_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n472_), .A2(KEYINPUT11), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n475_), .B1(new_n478_), .B2(new_n474_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n471_), .B(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n457_), .B1(new_n481_), .B2(KEYINPUT17), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(KEYINPUT17), .B2(new_n457_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT79), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n483_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n453_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT80), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n391_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n423_), .B1(new_n490_), .B2(new_n418_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT67), .B1(new_n412_), .B2(new_n396_), .ZN(new_n492_));
  AOI211_X1 g291(.A(new_n405_), .B(new_n395_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n424_), .A2(KEYINPUT69), .A3(new_n428_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n428_), .B1(new_n424_), .B2(KEYINPUT69), .ZN(new_n496_));
  OAI22_X1  g295(.A1(new_n495_), .A2(new_n496_), .B1(KEYINPUT69), .B2(new_n424_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n497_), .A3(new_n480_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G230gat), .A2(G233gat), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n498_), .A2(KEYINPUT71), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT71), .B1(new_n498_), .B2(new_n499_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n479_), .B(new_n504_), .C1(new_n414_), .C2(new_n430_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n480_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT12), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(KEYINPUT70), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n505_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT72), .B1(new_n502_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT71), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n414_), .A2(new_n430_), .A3(new_n479_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n499_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n498_), .A2(KEYINPUT71), .A3(new_n499_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT72), .ZN(new_n517_));
  INV_X1    g316(.A(new_n509_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n510_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n513_), .B1(new_n512_), .B2(new_n506_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT5), .B(G176gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G204gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G120gat), .B(G148gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n522_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n520_), .A2(new_n521_), .A3(new_n527_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(KEYINPUT13), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(KEYINPUT13), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT81), .B(G113gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT82), .B(G141gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n463_), .A2(new_n467_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n384_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n468_), .A2(new_n437_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n383_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n546_), .B2(new_n544_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n540_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n468_), .B(new_n383_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n549_), .B(new_n539_), .C1(new_n550_), .C2(new_n543_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(KEYINPUT83), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT83), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n553_), .B(new_n540_), .C1(new_n545_), .C2(new_n547_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n534_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n380_), .A2(new_n489_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT98), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT98), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n380_), .A2(new_n489_), .A3(new_n560_), .A4(new_n557_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n562_), .A2(G1gat), .A3(new_n239_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT38), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT99), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n563_), .A2(new_n564_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n449_), .B1(new_n370_), .B2(new_n379_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n557_), .A3(new_n486_), .ZN(new_n569_));
  OAI21_X1  g368(.A(G1gat), .B1(new_n569_), .B2(new_n239_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT99), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n563_), .A2(new_n571_), .A3(new_n564_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n566_), .A2(new_n567_), .A3(new_n570_), .A4(new_n572_), .ZN(G1324gat));
  NOR2_X1   g372(.A1(new_n377_), .A2(G8gat), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n559_), .A2(new_n561_), .A3(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n568_), .A2(new_n557_), .A3(new_n486_), .A4(new_n376_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT39), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(new_n577_), .A3(G8gat), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n577_), .B1(new_n576_), .B2(G8gat), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n575_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT101), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT101), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n575_), .B(new_n582_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n581_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(G1325gat));
  INV_X1    g386(.A(new_n343_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G15gat), .B1(new_n569_), .B2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT41), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n562_), .A2(G15gat), .A3(new_n588_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(G1326gat));
  OAI21_X1  g391(.A(G22gat), .B1(new_n569_), .B2(new_n367_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT42), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n367_), .A2(G22gat), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n594_), .B1(new_n562_), .B2(new_n595_), .ZN(G1327gat));
  INV_X1    g395(.A(new_n449_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n370_), .B2(new_n379_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n534_), .A2(new_n556_), .A3(new_n486_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(G29gat), .B1(new_n600_), .B2(new_n238_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n453_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT43), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT102), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n367_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n378_), .A2(new_n239_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n376_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n602_), .B(new_n604_), .C1(new_n607_), .C2(new_n369_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n453_), .B1(new_n370_), .B2(new_n379_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n603_), .A2(KEYINPUT102), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n599_), .B(new_n608_), .C1(new_n609_), .C2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT44), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n613_), .A2(KEYINPUT103), .A3(new_n614_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT103), .B1(new_n613_), .B2(new_n614_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n618_), .A2(new_n239_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n601_), .B1(new_n620_), .B2(G29gat), .ZN(G1328gat));
  OAI211_X1 g420(.A(new_n376_), .B(new_n615_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G36gat), .ZN(new_n623_));
  INV_X1    g422(.A(G36gat), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n598_), .A2(new_n624_), .A3(new_n376_), .A4(new_n599_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT45), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT46), .ZN(new_n629_));
  AOI22_X1  g428(.A1(new_n623_), .A2(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  AOI211_X1 g430(.A(new_n631_), .B(new_n626_), .C1(new_n622_), .C2(G36gat), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(G1329gat));
  AND2_X1   g432(.A1(new_n600_), .A2(new_n343_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(G43gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n339_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G43gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n635_), .B1(new_n618_), .B2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g438(.A(G50gat), .B1(new_n618_), .B2(new_n367_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n367_), .A2(G50gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT105), .Z(new_n642_));
  NAND2_X1  g441(.A1(new_n600_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(G1331gat));
  AND2_X1   g443(.A1(new_n489_), .A2(new_n534_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT106), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n555_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n647_), .B(new_n380_), .C1(new_n646_), .C2(new_n645_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n239_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n568_), .A2(new_n556_), .A3(new_n534_), .A4(new_n486_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n238_), .ZN(new_n652_));
  MUX2_X1   g451(.A(new_n649_), .B(new_n652_), .S(G57gat), .Z(G1332gat));
  NOR2_X1   g452(.A1(new_n377_), .A2(G64gat), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n648_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G64gat), .B1(new_n650_), .B2(new_n377_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT48), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n656_), .A2(KEYINPUT107), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1333gat));
  INV_X1    g462(.A(G71gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n651_), .B2(new_n343_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n666_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n343_), .A2(new_n664_), .ZN(new_n669_));
  OAI22_X1  g468(.A1(new_n667_), .A2(new_n668_), .B1(new_n648_), .B2(new_n669_), .ZN(G1334gat));
  OAI21_X1  g469(.A(G78gat), .B1(new_n650_), .B2(new_n367_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT50), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n367_), .A2(G78gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n648_), .B2(new_n673_), .ZN(G1335gat));
  INV_X1    g473(.A(new_n486_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n534_), .A2(new_n556_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n598_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT109), .ZN(new_n679_));
  AOI21_X1  g478(.A(G85gat), .B1(new_n679_), .B2(new_n238_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n609_), .A2(new_n612_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n608_), .A3(new_n677_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n239_), .A2(new_n408_), .A3(new_n407_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1336gat));
  AOI21_X1  g484(.A(G92gat), .B1(new_n679_), .B2(new_n376_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n682_), .A2(new_n299_), .A3(new_n377_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1337gat));
  NAND3_X1  g487(.A1(new_n679_), .A2(new_n490_), .A3(new_n636_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G99gat), .B1(new_n682_), .B2(new_n588_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT111), .Z(new_n693_));
  XNOR2_X1  g492(.A(new_n691_), .B(new_n693_), .ZN(G1338gat));
  OAI21_X1  g493(.A(G106gat), .B1(new_n682_), .B2(new_n367_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n679_), .A2(new_n418_), .A3(new_n368_), .ZN(new_n699_));
  OAI211_X1 g498(.A(G106gat), .B(new_n696_), .C1(new_n682_), .C2(new_n367_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT53), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT53), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n698_), .A2(new_n703_), .A3(new_n699_), .A4(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1339gat));
  INV_X1    g504(.A(KEYINPUT119), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT57), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT114), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n555_), .A2(new_n710_), .A3(new_n529_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n555_), .B2(new_n529_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT55), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n502_), .A2(KEYINPUT72), .A3(new_n509_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n517_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT115), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n499_), .B1(new_n518_), .B2(new_n498_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n502_), .A2(new_n509_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(KEYINPUT55), .B2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n520_), .A2(KEYINPUT115), .A3(new_n714_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n719_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n724_), .A2(KEYINPUT56), .A3(new_n526_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT56), .B1(new_n724_), .B2(new_n526_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n713_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n550_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n543_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n542_), .A2(new_n544_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n729_), .B(new_n540_), .C1(new_n543_), .C2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n551_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n531_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n449_), .B(new_n709_), .C1(new_n727_), .C2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n711_), .A2(new_n712_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n724_), .A2(new_n526_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT56), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n724_), .A2(KEYINPUT56), .A3(new_n526_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n597_), .B(new_n737_), .C1(new_n743_), .C2(new_n733_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n735_), .B1(new_n709_), .B2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n530_), .A2(new_n732_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT58), .B(new_n746_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT118), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n741_), .A2(new_n742_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT118), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(KEYINPUT58), .A4(new_n746_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n746_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT116), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n746_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n754_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n752_), .A2(new_n758_), .A3(new_n602_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n486_), .B1(new_n745_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n534_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n675_), .A2(new_n555_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT54), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n761_), .A2(new_n453_), .A3(new_n762_), .A4(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(KEYINPUT54), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n636_), .B(new_n367_), .C1(new_n760_), .C2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n376_), .A2(new_n239_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT120), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n752_), .A2(new_n758_), .A3(new_n602_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n597_), .B(new_n708_), .C1(new_n743_), .C2(new_n733_), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n449_), .B(new_n736_), .C1(new_n727_), .C2(new_n734_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n708_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n675_), .B1(new_n772_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n766_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n765_), .B(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n368_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT120), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n636_), .A4(new_n769_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n771_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(G113gat), .B1(new_n782_), .B2(new_n555_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT121), .ZN(new_n784_));
  OAI21_X1  g583(.A(G113gat), .B1(new_n556_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT59), .B1(new_n768_), .B2(new_n770_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT59), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n779_), .A2(new_n787_), .A3(new_n636_), .A4(new_n769_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n784_), .A2(G113gat), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n786_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n783_), .B1(new_n785_), .B2(new_n790_), .ZN(G1340gat));
  NAND3_X1  g590(.A1(new_n786_), .A2(new_n788_), .A3(new_n534_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT122), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT122), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n786_), .A2(new_n788_), .A3(new_n794_), .A4(new_n534_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(G120gat), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(G120gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n761_), .B2(KEYINPUT60), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n782_), .B(new_n798_), .C1(KEYINPUT60), .C2(new_n797_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n799_), .ZN(G1341gat));
  AOI21_X1  g599(.A(G127gat), .B1(new_n782_), .B2(new_n486_), .ZN(new_n801_));
  AND4_X1   g600(.A1(G127gat), .A2(new_n786_), .A3(new_n486_), .A4(new_n788_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1342gat));
  AOI21_X1  g602(.A(G134gat), .B1(new_n782_), .B2(new_n449_), .ZN(new_n804_));
  AND4_X1   g603(.A1(G134gat), .A2(new_n786_), .A3(new_n602_), .A4(new_n788_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1343gat));
  NAND2_X1  g605(.A1(new_n776_), .A2(new_n778_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n343_), .A2(new_n367_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n769_), .A3(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n556_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT123), .B(G141gat), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(G1344gat));
  NOR2_X1   g611(.A1(new_n809_), .A2(new_n761_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g613(.A1(new_n809_), .A2(new_n675_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT61), .B(G155gat), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n815_), .B(new_n816_), .Z(G1346gat));
  AND2_X1   g616(.A1(new_n807_), .A2(new_n808_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n818_), .A2(G162gat), .A3(new_n602_), .A4(new_n769_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n206_), .B1(new_n809_), .B2(new_n597_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT124), .ZN(G1347gat));
  NAND2_X1  g621(.A1(new_n779_), .A2(new_n343_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n377_), .A2(new_n238_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT62), .B(G169gat), .C1(new_n827_), .C2(new_n556_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n823_), .A2(new_n556_), .A3(new_n825_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n251_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n254_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n831_), .A3(new_n832_), .ZN(G1348gat));
  NAND2_X1  g632(.A1(new_n826_), .A2(new_n534_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g634(.A(G183gat), .B1(new_n827_), .B2(new_n675_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n826_), .A2(new_n486_), .A3(new_n259_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1350gat));
  OAI21_X1  g637(.A(G190gat), .B1(new_n827_), .B2(new_n453_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n449_), .A2(new_n258_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT125), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n827_), .B2(new_n841_), .ZN(G1351gat));
  NAND2_X1  g641(.A1(new_n818_), .A2(new_n824_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n556_), .ZN(new_n844_));
  INV_X1    g643(.A(G197gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1352gat));
  OAI22_X1  g645(.A1(new_n843_), .A2(new_n761_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT127), .Z(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  OAI221_X1 g650(.A(new_n849_), .B1(KEYINPUT126), .B2(G204gat), .C1(new_n843_), .C2(new_n761_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1353gat));
  NOR2_X1   g652(.A1(new_n843_), .A2(new_n675_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n855_));
  AND2_X1   g654(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n854_), .B2(new_n855_), .ZN(G1354gat));
  INV_X1    g657(.A(new_n843_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n859_), .A2(G218gat), .A3(new_n602_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G218gat), .B1(new_n859_), .B2(new_n449_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1355gat));
endmodule


