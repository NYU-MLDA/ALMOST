//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G190gat), .B(G218gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G232gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT34), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT35), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n211_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  INV_X1    g022(.A(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT9), .A3(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n226_), .A2(KEYINPUT9), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n218_), .A2(new_n222_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G43gat), .B(G50gat), .Z(new_n230_));
  INV_X1    g029(.A(G36gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G29gat), .ZN(new_n232_));
  INV_X1    g031(.A(G29gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G36gat), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n232_), .A2(new_n234_), .A3(KEYINPUT69), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT69), .B1(new_n232_), .B2(new_n234_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n230_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n233_), .A2(G36gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n231_), .A2(G29gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n232_), .A2(new_n234_), .A3(KEYINPUT69), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n237_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n246_));
  INV_X1    g045(.A(G99gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n220_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT64), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n251_), .A2(new_n246_), .A3(new_n247_), .A4(new_n220_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n249_), .A2(new_n218_), .A3(new_n250_), .A4(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT8), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n225_), .A2(new_n226_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n229_), .B(new_n245_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n213_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT71), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n253_), .A2(new_n255_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT8), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n267_), .A2(KEYINPUT70), .A3(new_n229_), .A4(new_n245_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n262_), .A2(new_n268_), .A3(KEYINPUT71), .A4(new_n213_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n237_), .A2(new_n244_), .A3(KEYINPUT15), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT15), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n235_), .A2(new_n236_), .A3(new_n230_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n243_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n256_), .A2(new_n257_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n229_), .B(KEYINPUT65), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n270_), .B(new_n274_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n269_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n212_), .B1(new_n263_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT72), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281_));
  INV_X1    g080(.A(new_n229_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n282_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT70), .B1(new_n283_), .B2(new_n245_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n281_), .B1(new_n260_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(new_n269_), .A3(new_n277_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(new_n212_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n280_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n261_), .A2(new_n262_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n277_), .B1(new_n211_), .B2(new_n210_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n207_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n286_), .A2(new_n287_), .A3(new_n212_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n287_), .B1(new_n286_), .B2(new_n212_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n207_), .B(new_n293_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n206_), .B1(new_n294_), .B2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n205_), .A2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n301_), .B(KEYINPUT74), .Z(new_n302_));
  NAND3_X1  g101(.A1(new_n289_), .A2(new_n293_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n299_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G113gat), .B(G120gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT88), .Z(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT31), .Z(new_n310_));
  AND2_X1   g109(.A1(new_n310_), .A2(KEYINPUT89), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT23), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G183gat), .A3(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT24), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319_));
  MUX2_X1   g118(.A(new_n318_), .B(KEYINPUT24), .S(new_n319_), .Z(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT85), .B(G190gat), .ZN(new_n321_));
  MUX2_X1   g120(.A(G190gat), .B(new_n321_), .S(KEYINPUT26), .Z(new_n322_));
  XOR2_X1   g121(.A(KEYINPUT25), .B(G183gat), .Z(new_n323_));
  OAI211_X1 g122(.A(new_n316_), .B(new_n320_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G176gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT86), .B1(new_n326_), .B2(G169gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT22), .B(G169gat), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n325_), .B(new_n327_), .C1(new_n328_), .C2(KEYINPUT86), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n313_), .A2(new_n315_), .A3(KEYINPUT87), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(KEYINPUT87), .B2(new_n315_), .ZN(new_n331_));
  INV_X1    g130(.A(G183gat), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n321_), .A2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n317_), .B(new_n329_), .C1(new_n331_), .C2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n324_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G227gat), .A2(G233gat), .ZN(new_n336_));
  INV_X1    g135(.A(G15gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT30), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n335_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341_));
  INV_X1    g140(.A(G43gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n340_), .B(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n311_), .A2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n310_), .A2(KEYINPUT89), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n344_), .B1(new_n311_), .B2(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(G197gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(G204gat), .ZN(new_n350_));
  INV_X1    g149(.A(G204gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(G197gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT21), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G211gat), .B(G218gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT95), .B1(new_n349_), .B2(G204gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT95), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n351_), .A3(G197gat), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n355_), .B(new_n357_), .C1(G197gat), .C2(new_n351_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n353_), .B(new_n354_), .C1(new_n358_), .C2(KEYINPUT21), .ZN(new_n359_));
  INV_X1    g158(.A(new_n354_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(KEYINPUT21), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT1), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G155gat), .A3(G162gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT91), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n363_), .B1(G155gat), .B2(G162gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n366_), .A2(KEYINPUT90), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT90), .B1(new_n366_), .B2(new_n367_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n365_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  OR2_X1    g169(.A1(G141gat), .A2(G148gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n371_), .A2(KEYINPUT3), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT2), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n371_), .A2(KEYINPUT3), .B1(new_n376_), .B2(new_n372_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT92), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n378_), .A2(new_n379_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n375_), .A2(new_n377_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n367_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n374_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n362_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G78gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n362_), .A2(KEYINPUT94), .B1(G228gat), .B2(G233gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(G22gat), .B(G50gat), .Z(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n387_), .A2(new_n388_), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n387_), .A2(new_n388_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n394_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n394_), .B1(new_n399_), .B2(new_n397_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n391_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT96), .B(G106gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n389_), .B(G78gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n397_), .A2(new_n399_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n394_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n408_), .A3(new_n400_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n403_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n404_), .B1(new_n403_), .B2(new_n409_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n335_), .A2(new_n362_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n316_), .B1(G183gat), .B2(G190gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n328_), .A2(new_n325_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n317_), .A3(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(KEYINPUT26), .B(G190gat), .Z(new_n418_));
  OAI21_X1  g217(.A(new_n320_), .B1(new_n323_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n417_), .B1(new_n419_), .B2(new_n331_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT20), .B1(new_n420_), .B2(new_n362_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT19), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n414_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n362_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n426_), .A2(KEYINPUT20), .ZN(new_n427_));
  INV_X1    g226(.A(new_n362_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(new_n334_), .A3(new_n324_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n423_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G8gat), .B(G36gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT18), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n433_), .B(new_n434_), .Z(new_n435_));
  NAND3_X1  g234(.A1(new_n425_), .A2(new_n431_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n435_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n423_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n439_), .B2(new_n424_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n385_), .B(new_n308_), .C1(new_n370_), .C2(new_n373_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G225gat), .A2(G233gat), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n442_), .B(new_n444_), .C1(new_n309_), .C2(new_n387_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G29gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(G85gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT0), .B(G57gat), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n447_), .B(new_n448_), .Z(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n445_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT98), .Z(new_n452_));
  OAI211_X1 g251(.A(new_n442_), .B(KEYINPUT4), .C1(new_n309_), .C2(new_n387_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT97), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n309_), .A2(new_n387_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n453_), .A2(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n309_), .A2(new_n387_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n458_), .A2(KEYINPUT97), .A3(KEYINPUT4), .A4(new_n442_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n443_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n441_), .B1(new_n452_), .B2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n443_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n444_), .B1(new_n458_), .B2(new_n442_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n449_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  OAI211_X1 g265(.A(KEYINPUT33), .B(new_n449_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n435_), .A2(KEYINPUT32), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n439_), .A2(new_n424_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n414_), .B1(KEYINPUT99), .B2(new_n421_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n421_), .A2(KEYINPUT99), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n423_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n430_), .A2(new_n423_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n470_), .B1(new_n477_), .B2(new_n469_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n464_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n462_), .A2(new_n449_), .A3(new_n463_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n412_), .B1(new_n468_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n403_), .A2(new_n409_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n404_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OR3_X1    g284(.A1(new_n462_), .A2(new_n449_), .A3(new_n463_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n403_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n485_), .A2(new_n464_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n435_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n436_), .A2(KEYINPUT27), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT100), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n438_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n437_), .B1(new_n492_), .B2(new_n475_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT100), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(KEYINPUT27), .A4(new_n436_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT27), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n441_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n491_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n488_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n348_), .B1(new_n482_), .B2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n498_), .A2(new_n412_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n486_), .A2(new_n464_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n502_), .A2(new_n348_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n305_), .B1(new_n500_), .B2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G127gat), .B(G155gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT16), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G183gat), .B(G211gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G57gat), .B(G64gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n511_));
  XOR2_X1   g310(.A(G71gat), .B(G78gat), .Z(new_n512_));
  OR2_X1    g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n512_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n513_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G8gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT14), .ZN(new_n519_));
  INV_X1    g318(.A(G8gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT78), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT78), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G8gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n519_), .B1(new_n524_), .B2(G1gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(G15gat), .B(G22gat), .Z(new_n526_));
  OAI21_X1  g325(.A(new_n518_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT78), .B(G8gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(new_n528_), .B2(new_n202_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n526_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n517_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n516_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT79), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n533_), .B(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n509_), .B1(new_n536_), .B2(KEYINPUT80), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT17), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(new_n536_), .B2(new_n509_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n283_), .A2(new_n516_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n283_), .A2(new_n516_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n542_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT66), .B(KEYINPUT12), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n283_), .B2(new_n516_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n542_), .B1(new_n283_), .B2(new_n516_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n513_), .B(KEYINPUT12), .C1(new_n515_), .C2(new_n514_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n552_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT68), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n555_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT13), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n274_), .A2(new_n270_), .A3(new_n531_), .A4(new_n527_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT81), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n565_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n237_), .A2(new_n244_), .A3(KEYINPUT81), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n532_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT82), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n564_), .A2(new_n568_), .A3(new_n569_), .A4(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT82), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n566_), .A2(new_n567_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n532_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n570_), .B1(new_n576_), .B2(new_n568_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n571_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT83), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G113gat), .B(G141gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G169gat), .B(G197gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n581_), .B(new_n582_), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(KEYINPUT83), .B(new_n571_), .C1(new_n573_), .C2(new_n577_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n580_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT84), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n578_), .A2(new_n587_), .A3(new_n583_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n586_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n505_), .A2(new_n541_), .A3(new_n563_), .A4(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n591_), .A2(KEYINPUT103), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(KEYINPUT103), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n202_), .B1(new_n594_), .B2(new_n502_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n303_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n299_), .A2(new_n598_), .A3(KEYINPUT77), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT77), .ZN(new_n600_));
  INV_X1    g399(.A(new_n206_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n293_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT76), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n603_), .B2(new_n297_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n604_), .B2(new_n597_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n602_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT75), .B1(new_n606_), .B2(new_n601_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT75), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(new_n608_), .A3(new_n206_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n609_), .A3(new_n303_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n599_), .A2(new_n605_), .B1(KEYINPUT37), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n541_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n563_), .A2(new_n590_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n500_), .B2(new_n504_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT101), .Z(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n202_), .A3(new_n502_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n595_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n617_), .A2(KEYINPUT38), .A3(new_n202_), .A4(new_n502_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(G1324gat));
  NAND3_X1  g424(.A1(new_n617_), .A2(new_n528_), .A3(new_n498_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  INV_X1    g426(.A(new_n498_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n591_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n629_), .B2(G8gat), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(new_n627_), .A3(G8gat), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n626_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n626_), .B(KEYINPUT40), .C1(new_n630_), .C2(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1325gat));
  INV_X1    g435(.A(new_n348_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n637_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G15gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT104), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n641_), .A3(G15gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT41), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(KEYINPUT41), .A3(new_n642_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n613_), .A2(new_n337_), .A3(new_n637_), .A4(new_n615_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(G1326gat));
  INV_X1    g447(.A(G22gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n594_), .B2(new_n412_), .ZN(new_n650_));
  XOR2_X1   g449(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n613_), .A2(new_n649_), .A3(new_n412_), .A4(new_n615_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1327gat));
  NAND2_X1  g453(.A1(new_n500_), .A2(new_n504_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n611_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT43), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n611_), .A2(new_n655_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n614_), .A2(new_n541_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(KEYINPUT44), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT44), .B1(new_n660_), .B2(new_n661_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n502_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G29gat), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n304_), .A2(new_n541_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n615_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n502_), .A2(new_n233_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT106), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n667_), .B1(new_n670_), .B2(new_n672_), .ZN(G1328gat));
  NAND3_X1  g472(.A1(new_n669_), .A2(new_n231_), .A3(new_n498_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT45), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n662_), .A2(new_n663_), .A3(new_n628_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(new_n231_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT46), .B(new_n675_), .C1(new_n676_), .C2(new_n231_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  AOI21_X1  g480(.A(G43gat), .B1(new_n669_), .B2(new_n637_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n348_), .A2(new_n342_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n664_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(G1330gat));
  AOI21_X1  g485(.A(G50gat), .B1(new_n669_), .B2(new_n412_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n412_), .A2(G50gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n664_), .B2(new_n688_), .ZN(G1331gat));
  NOR2_X1   g488(.A1(new_n563_), .A2(new_n590_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n655_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n613_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n666_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n563_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n590_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n505_), .A2(new_n541_), .A3(new_n694_), .A4(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G57gat), .B1(new_n666_), .B2(KEYINPUT107), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n697_), .B1(KEYINPUT107), .B2(G57gat), .ZN(new_n698_));
  OAI22_X1  g497(.A1(new_n693_), .A2(G57gat), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT108), .ZN(G1332gat));
  OAI21_X1  g499(.A(G64gat), .B1(new_n696_), .B2(new_n628_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT48), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n628_), .A2(G64gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n692_), .B2(new_n703_), .ZN(G1333gat));
  OAI21_X1  g503(.A(G71gat), .B1(new_n696_), .B2(new_n348_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT49), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n348_), .A2(G71gat), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT109), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n692_), .B2(new_n708_), .ZN(G1334gat));
  INV_X1    g508(.A(new_n412_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G78gat), .B1(new_n696_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT50), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n412_), .A2(new_n390_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n692_), .B2(new_n713_), .ZN(G1335gat));
  NAND2_X1  g513(.A1(new_n690_), .A2(new_n612_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G85gat), .B1(new_n717_), .B2(new_n666_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n691_), .A2(new_n668_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n502_), .A2(new_n223_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(G1336gat));
  OAI21_X1  g520(.A(G92gat), .B1(new_n717_), .B2(new_n628_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n498_), .A2(new_n224_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n719_), .B2(new_n723_), .ZN(G1337gat));
  AND3_X1   g523(.A1(new_n637_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n691_), .A2(new_n668_), .A3(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT110), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n247_), .B1(new_n716_), .B2(new_n637_), .ZN(new_n728_));
  OAI22_X1  g527(.A1(new_n727_), .A2(new_n728_), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n729_));
  NAND2_X1  g528(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT112), .Z(new_n731_));
  XNOR2_X1  g530(.A(new_n729_), .B(new_n731_), .ZN(G1338gat));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n716_), .A2(new_n412_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(G106gat), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT52), .B(new_n220_), .C1(new_n716_), .C2(new_n412_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n412_), .A2(new_n220_), .ZN(new_n737_));
  OAI22_X1  g536(.A1(new_n735_), .A2(new_n736_), .B1(new_n719_), .B2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g538(.A(KEYINPUT121), .ZN(new_n740_));
  NOR2_X1   g539(.A1(KEYINPUT120), .A2(G113gat), .ZN(new_n741_));
  AND2_X1   g540(.A1(KEYINPUT120), .A2(G113gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n590_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n610_), .A2(KEYINPUT37), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n576_), .A2(new_n568_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n583_), .B1(new_n745_), .B2(new_n570_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n564_), .A2(new_n568_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n570_), .B2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n589_), .B2(new_n588_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT116), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT116), .B(new_n748_), .C1(new_n589_), .C2(new_n588_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n555_), .A2(new_n561_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n554_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n549_), .A2(new_n543_), .A3(new_n553_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n542_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n549_), .A2(new_n550_), .A3(KEYINPUT55), .A4(new_n553_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n561_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(KEYINPUT56), .A3(new_n561_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n754_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n753_), .A2(KEYINPUT58), .A3(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT58), .B1(new_n753_), .B2(new_n765_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT77), .B1(new_n299_), .B2(new_n598_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n604_), .A2(new_n600_), .A3(new_n597_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n744_), .B(new_n768_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n761_), .A2(KEYINPUT114), .A3(new_n762_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n754_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n590_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n760_), .A2(KEYINPUT56), .A3(new_n561_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT56), .B1(new_n760_), .B2(new_n561_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(KEYINPUT114), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT115), .B1(new_n774_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n763_), .A2(new_n779_), .A3(new_n764_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n578_), .A2(new_n583_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT84), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n578_), .A2(new_n587_), .A3(new_n583_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n754_), .B1(new_n784_), .B2(new_n586_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n780_), .A2(new_n785_), .A3(new_n786_), .A4(new_n772_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT116), .B1(new_n784_), .B2(new_n748_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n752_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n562_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n778_), .A2(KEYINPUT117), .A3(new_n787_), .A4(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n299_), .A2(KEYINPUT117), .A3(new_n303_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n792_), .A3(KEYINPUT57), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n771_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n695_), .A2(new_n541_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT113), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n563_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT54), .B1(new_n611_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n744_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n799_), .A2(new_n563_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n612_), .A2(new_n797_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n501_), .A2(new_n502_), .A3(new_n637_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT59), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n807_), .ZN(new_n809_));
  XOR2_X1   g608(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n801_), .A2(new_n805_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n791_), .A2(new_n792_), .A3(KEYINPUT57), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT57), .B1(new_n791_), .B2(new_n792_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n541_), .B1(new_n815_), .B2(new_n771_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n809_), .B(new_n811_), .C1(new_n812_), .C2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n808_), .A2(new_n817_), .A3(KEYINPUT119), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n797_), .A2(new_n612_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n801_), .A2(new_n805_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n807_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n811_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n743_), .B1(new_n818_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G113gat), .B1(new_n821_), .B2(new_n590_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n740_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n825_), .ZN(new_n827_));
  NOR4_X1   g626(.A1(new_n806_), .A2(KEYINPUT119), .A3(new_n807_), .A4(new_n810_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n822_), .B1(new_n821_), .B2(new_n811_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n808_), .B2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT121), .B(new_n827_), .C1(new_n830_), .C2(new_n743_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n826_), .A2(new_n831_), .ZN(G1340gat));
  OAI21_X1  g631(.A(G120gat), .B1(new_n830_), .B2(new_n563_), .ZN(new_n833_));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n563_), .B2(KEYINPUT60), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n821_), .B(new_n835_), .C1(KEYINPUT60), .C2(new_n834_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(G1341gat));
  OAI21_X1  g636(.A(G127gat), .B1(new_n830_), .B2(new_n612_), .ZN(new_n838_));
  INV_X1    g637(.A(G127gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n821_), .A2(new_n839_), .A3(new_n541_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1342gat));
  OAI21_X1  g640(.A(G134gat), .B1(new_n830_), .B2(new_n802_), .ZN(new_n842_));
  INV_X1    g641(.A(G134gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n821_), .A2(new_n843_), .A3(new_n305_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1343gat));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  NOR4_X1   g645(.A1(new_n710_), .A2(new_n666_), .A3(new_n498_), .A4(new_n637_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n806_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n819_), .A2(new_n820_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(KEYINPUT122), .A3(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n590_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n694_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n852_), .B2(new_n541_), .ZN(new_n860_));
  AOI211_X1 g659(.A(KEYINPUT123), .B(new_n612_), .C1(new_n849_), .C2(new_n851_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT122), .B1(new_n850_), .B2(new_n847_), .ZN(new_n863_));
  AOI211_X1 g662(.A(new_n846_), .B(new_n848_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n541_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT123), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n852_), .A2(new_n859_), .A3(new_n541_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n857_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n862_), .A2(new_n868_), .ZN(G1346gat));
  INV_X1    g668(.A(new_n852_), .ZN(new_n870_));
  OR3_X1    g669(.A1(new_n870_), .A2(G162gat), .A3(new_n304_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G162gat), .B1(new_n870_), .B2(new_n802_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1347gat));
  AOI21_X1  g672(.A(new_n628_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n874_), .A2(new_n710_), .A3(new_n503_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n590_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G169gat), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n875_), .A2(new_n590_), .A3(new_n328_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n876_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .ZN(G1348gat));
  NAND3_X1  g681(.A1(new_n874_), .A2(new_n710_), .A3(new_n503_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n563_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n325_), .ZN(G1349gat));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n612_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n323_), .B1(new_n887_), .B2(new_n332_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n887_), .A2(G183gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n886_), .B2(new_n890_), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n883_), .B2(new_n802_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n304_), .A2(new_n418_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n883_), .B2(new_n893_), .ZN(G1351gat));
  NOR2_X1   g693(.A1(new_n488_), .A2(new_n637_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n498_), .B(new_n895_), .C1(new_n812_), .C2(new_n816_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n874_), .A2(KEYINPUT125), .A3(new_n895_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n695_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n349_), .ZN(G1352gat));
  AOI21_X1  g700(.A(new_n563_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n351_), .A2(KEYINPUT126), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n351_), .A2(KEYINPUT126), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n902_), .B2(new_n904_), .ZN(G1353gat));
  NAND2_X1  g705(.A1(new_n898_), .A2(new_n899_), .ZN(new_n907_));
  OR2_X1    g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  AND4_X1   g708(.A1(new_n541_), .A2(new_n907_), .A3(new_n908_), .A4(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n907_), .B2(new_n541_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1354gat));
  NAND2_X1  g711(.A1(new_n611_), .A2(G218gat), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n913_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n304_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n915_));
  AOI21_X1  g714(.A(G218gat), .B1(new_n915_), .B2(KEYINPUT127), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n896_), .A2(new_n897_), .ZN(new_n917_));
  AOI21_X1  g716(.A(KEYINPUT125), .B1(new_n874_), .B2(new_n895_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n305_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n914_), .B1(new_n916_), .B2(new_n921_), .ZN(G1355gat));
endmodule


