//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT85), .B(G43gat), .Z(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT83), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT83), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n212_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n223_), .A2(new_n214_), .A3(new_n213_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  INV_X1    g024(.A(G183gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT25), .B1(new_n226_), .B2(KEYINPUT81), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(G183gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n225_), .A2(KEYINPUT82), .A3(new_n227_), .A4(new_n230_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n224_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n220_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n210_), .A2(new_n211_), .ZN(new_n237_));
  INV_X1    g036(.A(G190gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n226_), .B2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(new_n223_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT22), .B1(new_n221_), .B2(KEYINPUT84), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n222_), .B(new_n241_), .C1(new_n242_), .C2(KEYINPUT84), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT30), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n220_), .A2(new_n235_), .B1(new_n243_), .B2(new_n240_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT30), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G227gat), .A2(G233gat), .ZN(new_n251_));
  INV_X1    g050(.A(G15gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G71gat), .ZN(new_n254_));
  INV_X1    g053(.A(G99gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n247_), .A2(new_n258_), .A3(new_n249_), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n207_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n264_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(new_n206_), .A3(new_n262_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G197gat), .ZN(new_n269_));
  INV_X1    g068(.A(G204gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT90), .B(G204gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(new_n269_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G211gat), .B(G218gat), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n270_), .A2(KEYINPUT90), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT90), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G204gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(G197gat), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT91), .ZN(new_n281_));
  OAI22_X1  g080(.A1(new_n280_), .A2(new_n281_), .B1(new_n269_), .B2(G204gat), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n272_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT21), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n275_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT92), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(KEYINPUT92), .A3(new_n286_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n276_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G141gat), .ZN(new_n292_));
  INV_X1    g091(.A(G148gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G141gat), .A2(G148gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT1), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT88), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n298_), .B(new_n300_), .C1(KEYINPUT1), .C2(new_n296_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n297_), .A2(KEYINPUT88), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n294_), .B(new_n295_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n294_), .A2(KEYINPUT3), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n294_), .A2(KEYINPUT3), .B1(new_n305_), .B2(new_n295_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT89), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n304_), .A2(new_n306_), .A3(new_n309_), .A4(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n303_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G228gat), .ZN(new_n317_));
  INV_X1    g116(.A(G233gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n291_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n291_), .A2(KEYINPUT93), .ZN(new_n322_));
  INV_X1    g121(.A(new_n276_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n284_), .A2(KEYINPUT92), .A3(new_n286_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT92), .B1(new_n284_), .B2(new_n286_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT93), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n316_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n319_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n321_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G78gat), .B(G106gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT95), .ZN(new_n334_));
  INV_X1    g133(.A(new_n332_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n335_), .B(new_n321_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n333_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT94), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n314_), .A2(new_n315_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G22gat), .B(G50gat), .Z(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT28), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n341_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n337_), .A2(new_n338_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n344_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n316_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n291_), .A2(KEYINPUT93), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n326_), .A2(new_n327_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n349_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n319_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n335_), .B1(new_n353_), .B2(new_n321_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n336_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT95), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n333_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n348_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n268_), .B1(new_n346_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n291_), .A2(new_n248_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G169gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n222_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n223_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT96), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n364_), .A2(new_n239_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(KEYINPUT96), .A3(new_n363_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n216_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT25), .B(G183gat), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n224_), .B1(new_n225_), .B2(new_n368_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n365_), .A2(new_n366_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n360_), .B(KEYINPUT20), .C1(new_n291_), .C2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n291_), .B2(new_n370_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n326_), .B2(new_n245_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G8gat), .B(G36gat), .Z(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT18), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n374_), .A2(new_n383_), .A3(new_n378_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT27), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n314_), .A2(KEYINPUT97), .A3(new_n204_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n204_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT97), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n392_), .B1(new_n313_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n314_), .A2(KEYINPUT4), .A3(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n394_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n396_), .B1(new_n397_), .B2(KEYINPUT4), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n395_), .B1(new_n398_), .B2(new_n391_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G1gat), .B(G29gat), .Z(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT98), .B(G85gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT0), .B(G57gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n399_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n371_), .A2(new_n373_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n373_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n322_), .A2(new_n328_), .A3(new_n370_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n377_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n384_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(KEYINPUT27), .A3(new_n386_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n389_), .A2(new_n406_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n345_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n268_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n265_), .A2(new_n267_), .A3(KEYINPUT87), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n356_), .A2(new_n348_), .A3(new_n357_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n415_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n359_), .A2(new_n414_), .A3(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n398_), .A2(new_n391_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n391_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n424_), .A2(new_n404_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT33), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n399_), .A2(new_n404_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n399_), .A2(KEYINPUT33), .A3(new_n404_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n428_), .A2(new_n385_), .A3(new_n386_), .A4(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n383_), .A2(KEYINPUT32), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n431_), .B(KEYINPUT99), .Z(new_n432_));
  NAND3_X1  g231(.A1(new_n374_), .A2(new_n432_), .A3(new_n378_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT100), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT32), .B(new_n383_), .C1(new_n407_), .C2(new_n410_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n434_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n435_), .A2(new_n405_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n419_), .B1(new_n430_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n415_), .A2(new_n420_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n422_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G230gat), .A2(G233gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(G78gat), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n446_), .ZN(new_n448_));
  INV_X1    g247(.A(G78gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n444_), .ZN(new_n450_));
  INV_X1    g249(.A(G64gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G57gat), .ZN(new_n452_));
  INV_X1    g251(.A(G57gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G64gat), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n452_), .A2(new_n454_), .A3(KEYINPUT11), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT11), .B1(new_n452_), .B2(new_n454_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n447_), .B(new_n450_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n452_), .A2(new_n454_), .A3(KEYINPUT11), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n449_), .B1(new_n448_), .B2(new_n444_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n445_), .A2(new_n446_), .A3(G78gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n457_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n462_), .B1(new_n457_), .B2(new_n461_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT10), .B(G99gat), .Z(new_n467_));
  INV_X1    g266(.A(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G85gat), .B(G92gat), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT9), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G99gat), .A2(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(G99gat), .A3(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G85gat), .ZN(new_n477_));
  INV_X1    g276(.A(G92gat), .ZN(new_n478_));
  OR3_X1    g277(.A1(new_n477_), .A2(new_n478_), .A3(KEYINPUT9), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n469_), .A2(new_n471_), .A3(new_n476_), .A4(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(KEYINPUT65), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT65), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n473_), .A2(new_n475_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n255_), .A3(new_n468_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n482_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n481_), .B1(new_n489_), .B2(new_n470_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n470_), .A2(new_n481_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT64), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n473_), .A2(new_n475_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n486_), .A2(new_n487_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n476_), .A2(KEYINPUT64), .A3(new_n486_), .A4(new_n487_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n491_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n480_), .B1(new_n490_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n466_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n480_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n473_), .A2(new_n475_), .A3(new_n483_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n483_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n494_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n470_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT8), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n491_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n496_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT64), .B1(new_n488_), .B2(new_n476_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n500_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n457_), .A2(new_n461_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT67), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n463_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n443_), .B1(new_n499_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT68), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n498_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT68), .B(new_n480_), .C1(new_n490_), .C2(new_n497_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n511_), .A2(KEYINPUT69), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT69), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n457_), .A2(new_n461_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n519_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n518_), .A3(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n519_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n443_), .B1(new_n466_), .B2(new_n498_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n514_), .A2(KEYINPUT70), .A3(new_n443_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n515_), .B1(new_n527_), .B2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G176gat), .B(G204gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT72), .ZN(new_n535_));
  XOR2_X1   g334(.A(G120gat), .B(G148gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  OR2_X1    g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n539_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n542_), .A2(KEYINPUT13), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(KEYINPUT13), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G29gat), .B(G36gat), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n549_), .A2(KEYINPUT73), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(KEYINPUT73), .ZN(new_n551_));
  XOR2_X1   g350(.A(G43gat), .B(G50gat), .Z(new_n552_));
  OR3_X1    g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G15gat), .B(G22gat), .ZN(new_n554_));
  INV_X1    g353(.A(G1gat), .ZN(new_n555_));
  INV_X1    g354(.A(G8gat), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT14), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G1gat), .B(G8gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n552_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n553_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n553_), .B2(new_n561_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n548_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT77), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(KEYINPUT77), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n553_), .A2(new_n561_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT15), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n560_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n563_), .A2(new_n548_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n566_), .A2(new_n567_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT78), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n571_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n567_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n574_), .B1(new_n575_), .B2(new_n565_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT78), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G113gat), .B(G141gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT79), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G169gat), .B(G197gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  NAND3_X1  g381(.A1(new_n573_), .A2(new_n578_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT80), .B1(new_n572_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n573_), .A2(new_n578_), .A3(KEYINPUT80), .A4(new_n582_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n546_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n442_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n569_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n595_));
  AOI211_X1 g394(.A(KEYINPUT74), .B(new_n595_), .C1(new_n510_), .C2(new_n568_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n591_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n594_), .B1(new_n591_), .B2(new_n596_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  OR4_X1    g400(.A1(KEYINPUT36), .A2(new_n597_), .A3(new_n598_), .A4(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(KEYINPUT36), .Z(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(KEYINPUT75), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n602_), .A2(KEYINPUT75), .A3(KEYINPUT37), .A4(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT76), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n560_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n520_), .A2(new_n522_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n613_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n617_));
  XOR2_X1   g416(.A(G127gat), .B(G155gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT16), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G183gat), .B(G211gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  OR4_X1    g420(.A1(new_n610_), .A2(new_n616_), .A3(new_n617_), .A4(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(KEYINPUT17), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n614_), .A2(new_n513_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n613_), .A2(new_n466_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n609_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n590_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT101), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n555_), .A3(new_n405_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n413_), .B1(new_n440_), .B2(new_n268_), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n634_), .A2(new_n421_), .B1(new_n440_), .B2(new_n439_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n602_), .A2(new_n604_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n635_), .A2(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n546_), .A2(new_n627_), .A3(new_n588_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n406_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n631_), .A2(new_n632_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n633_), .A2(new_n644_), .A3(new_n645_), .ZN(G1324gat));
  NAND2_X1  g445(.A1(new_n389_), .A2(new_n412_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n630_), .A2(new_n556_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  INV_X1    g448(.A(new_n643_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n647_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n647_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT103), .B1(new_n643_), .B2(new_n653_), .ZN(new_n654_));
  AND4_X1   g453(.A1(new_n649_), .A2(new_n652_), .A3(G8gat), .A4(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n643_), .A2(new_n653_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n556_), .B1(new_n656_), .B2(new_n651_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n649_), .B1(new_n657_), .B2(new_n654_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n648_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT40), .B(new_n648_), .C1(new_n655_), .C2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  NAND3_X1  g462(.A1(new_n630_), .A2(new_n252_), .A3(new_n419_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n650_), .A2(new_n419_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n665_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT41), .B1(new_n665_), .B2(G15gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n664_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(G1326gat));
  INV_X1    g469(.A(G22gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n440_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n630_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G22gat), .B1(new_n643_), .B2(new_n440_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(KEYINPUT42), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(KEYINPUT42), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1327gat));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n442_), .B2(new_n609_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n609_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT43), .B(new_n682_), .C1(new_n422_), .C2(new_n441_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n627_), .B(new_n589_), .C1(new_n681_), .C2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT43), .B1(new_n635_), .B2(new_n682_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n442_), .A2(new_n680_), .A3(new_n609_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n689_), .A2(KEYINPUT44), .A3(new_n627_), .A4(new_n589_), .ZN(new_n690_));
  AND4_X1   g489(.A1(G29gat), .A2(new_n686_), .A3(new_n405_), .A4(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n640_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n627_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n590_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n405_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n691_), .A2(new_n696_), .ZN(G1328gat));
  NOR2_X1   g496(.A1(new_n653_), .A2(G36gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n590_), .A2(new_n694_), .A3(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n686_), .A2(new_n647_), .A3(new_n690_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(G36gat), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(KEYINPUT107), .A3(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(KEYINPUT107), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n704_), .A2(KEYINPUT107), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n703_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(new_n268_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n686_), .A2(new_n690_), .A3(G43gat), .A4(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n695_), .A2(new_n419_), .ZN(new_n712_));
  XOR2_X1   g511(.A(KEYINPUT108), .B(G43gat), .Z(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g514(.A(G50gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n695_), .A2(new_n716_), .A3(new_n672_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n686_), .A2(new_n672_), .A3(new_n690_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G50gat), .B1(new_n718_), .B2(new_n719_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1331gat));
  INV_X1    g521(.A(new_n588_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n545_), .A2(new_n723_), .A3(new_n627_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n641_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G57gat), .B1(new_n726_), .B2(new_n406_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n545_), .A2(new_n723_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n442_), .A2(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(new_n628_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n453_), .A3(new_n405_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n731_), .ZN(G1332gat));
  AOI21_X1  g531(.A(new_n451_), .B1(new_n725_), .B2(new_n647_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT48), .Z(new_n734_));
  NAND2_X1  g533(.A1(new_n647_), .A2(new_n451_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT110), .Z(new_n736_));
  NAND2_X1  g535(.A1(new_n730_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(G1333gat));
  INV_X1    g537(.A(G71gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n730_), .A2(new_n739_), .A3(new_n419_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n725_), .A2(new_n419_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G71gat), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(KEYINPUT49), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(KEYINPUT49), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(KEYINPUT111), .B(new_n740_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  AOI21_X1  g548(.A(new_n449_), .B1(new_n725_), .B2(new_n672_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT50), .Z(new_n751_));
  NOR2_X1   g550(.A1(new_n440_), .A2(G78gat), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT112), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n730_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n754_), .ZN(G1335gat));
  AOI21_X1  g554(.A(new_n693_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n728_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n406_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n729_), .A2(new_n694_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(new_n477_), .A3(new_n405_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1336gat));
  OAI21_X1  g560(.A(G92gat), .B1(new_n757_), .B2(new_n653_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n478_), .A3(new_n647_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n756_), .A2(new_n419_), .A3(new_n728_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n710_), .A2(new_n467_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n765_), .A2(G99gat), .B1(new_n759_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n767_), .B(new_n768_), .Z(G1338gat));
  NAND3_X1  g568(.A1(new_n759_), .A2(new_n468_), .A3(new_n672_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n756_), .A2(new_n672_), .A3(new_n728_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(G106gat), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n771_), .B2(G106gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n770_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n770_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n627_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n545_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n545_), .A2(KEYINPUT114), .A3(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n781_), .B1(new_n787_), .B2(new_n682_), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT54), .B(new_n609_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n586_), .A2(new_n541_), .A3(new_n587_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT70), .B1(new_n514_), .B2(new_n443_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n443_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n529_), .B(new_n794_), .C1(new_n510_), .C2(new_n513_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n796_), .B2(new_n526_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n524_), .A2(new_n514_), .A3(new_n525_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n794_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(KEYINPUT115), .A3(new_n794_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n527_), .A2(new_n532_), .A3(KEYINPUT55), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n797_), .A2(new_n801_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n539_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n805_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(KEYINPUT116), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n809_), .B(KEYINPUT56), .C1(new_n804_), .C2(new_n805_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n791_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT117), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n791_), .B(new_n813_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n563_), .A2(new_n547_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n570_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n547_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n817_), .A2(new_n582_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n572_), .A2(new_n584_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n542_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n812_), .A2(new_n814_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n692_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n820_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n811_), .B2(KEYINPUT117), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n640_), .B1(new_n826_), .B2(new_n814_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT57), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n819_), .A2(new_n541_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n807_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n806_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n609_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(KEYINPUT58), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n609_), .B(KEYINPUT119), .C1(new_n831_), .C2(new_n832_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n824_), .A2(new_n828_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n790_), .B1(new_n839_), .B2(new_n627_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n647_), .A2(new_n406_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(new_n440_), .A3(new_n710_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT59), .B1(new_n843_), .B2(KEYINPUT122), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(KEYINPUT122), .B2(new_n843_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n840_), .A2(new_n845_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT123), .B(G113gat), .Z(new_n847_));
  NAND2_X1  g646(.A1(new_n723_), .A2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n838_), .B1(new_n827_), .B2(KEYINPUT57), .ZN(new_n849_));
  AOI211_X1 g648(.A(new_n823_), .B(new_n640_), .C1(new_n826_), .C2(new_n814_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n627_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n788_), .A2(new_n789_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n842_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT121), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(KEYINPUT59), .C1(new_n840_), .C2(new_n842_), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n846_), .B(new_n848_), .C1(new_n855_), .C2(new_n857_), .ZN(new_n858_));
  AOI211_X1 g657(.A(new_n588_), .B(new_n842_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT120), .B1(new_n859_), .B2(G113gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n853_), .A2(new_n723_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862_));
  INV_X1    g661(.A(G113gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n858_), .A2(new_n865_), .ZN(G1340gat));
  INV_X1    g665(.A(G120gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n545_), .B2(KEYINPUT60), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n853_), .B(new_n868_), .C1(KEYINPUT60), .C2(new_n867_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n546_), .B1(new_n840_), .B2(new_n845_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n871_), .B2(new_n867_), .ZN(G1341gat));
  AOI21_X1  g671(.A(G127gat), .B1(new_n853_), .B2(new_n693_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n846_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n693_), .A2(G127gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1342gat));
  AOI21_X1  g675(.A(G134gat), .B1(new_n853_), .B2(new_n640_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n609_), .A2(G134gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n874_), .B2(new_n878_), .ZN(G1343gat));
  NAND2_X1  g678(.A1(new_n851_), .A2(new_n852_), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n440_), .A2(new_n647_), .A3(new_n419_), .A4(new_n406_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n588_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n292_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n545_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n293_), .ZN(G1345gat));
  OAI21_X1  g685(.A(KEYINPUT124), .B1(new_n882_), .B2(new_n627_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n880_), .A2(new_n888_), .A3(new_n693_), .A4(new_n881_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT61), .B(G155gat), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n887_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n882_), .B2(new_n682_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n692_), .A2(G162gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n882_), .B2(new_n895_), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n653_), .A2(new_n405_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n440_), .A2(new_n419_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n880_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G169gat), .B1(new_n899_), .B2(new_n588_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n899_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(new_n723_), .A3(new_n361_), .ZN(new_n904_));
  OAI211_X1 g703(.A(KEYINPUT62), .B(G169gat), .C1(new_n899_), .C2(new_n588_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n902_), .A2(new_n904_), .A3(new_n905_), .ZN(G1348gat));
  NOR2_X1   g705(.A1(new_n899_), .A2(new_n545_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n222_), .ZN(G1349gat));
  NOR3_X1   g707(.A1(new_n899_), .A2(new_n627_), .A3(new_n368_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n903_), .A2(new_n693_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n226_), .B2(new_n910_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n899_), .B2(new_n682_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n640_), .A2(new_n225_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n899_), .B2(new_n913_), .ZN(G1351gat));
  NOR2_X1   g713(.A1(new_n440_), .A2(new_n419_), .ZN(new_n915_));
  AND3_X1   g714(.A1(new_n880_), .A2(new_n897_), .A3(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n723_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT125), .B(G197gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n916_), .B(new_n723_), .C1(KEYINPUT125), .C2(G197gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1352gat));
  NAND2_X1  g720(.A1(new_n916_), .A2(new_n546_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n272_), .ZN(new_n923_));
  AOI21_X1  g722(.A(G204gat), .B1(new_n916_), .B2(new_n546_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1353gat));
  AOI21_X1  g724(.A(new_n627_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n880_), .A2(new_n897_), .A3(new_n915_), .A4(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n927_), .A2(KEYINPUT127), .A3(new_n928_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n928_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n916_), .A2(KEYINPUT126), .A3(new_n933_), .A4(new_n926_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n931_), .A2(new_n932_), .B1(new_n934_), .B2(new_n936_), .ZN(G1354gat));
  INV_X1    g736(.A(G218gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n916_), .A2(new_n938_), .A3(new_n640_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n916_), .A2(new_n609_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n938_), .ZN(G1355gat));
endmodule


