//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT80), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT80), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(G169gat), .B2(G176gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT81), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT82), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .A4(KEYINPUT24), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n209_), .B(KEYINPUT81), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT24), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT82), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT83), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT23), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n217_), .A2(KEYINPUT83), .A3(G183gat), .A4(G190gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n205_), .A2(new_n207_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT24), .ZN(new_n226_));
  OR2_X1    g025(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n225_), .A2(new_n226_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n213_), .A2(new_n216_), .A3(new_n224_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n222_), .A2(new_n218_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(G183gat), .B2(G190gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G169gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT84), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n236_), .B1(new_n203_), .B2(KEYINPUT22), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n204_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n234_), .B(new_n211_), .C1(new_n237_), .C2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G197gat), .B(G204gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT21), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G197gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(G204gat), .ZN(new_n246_));
  INV_X1    g045(.A(G204gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(G197gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT21), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G211gat), .B(G218gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n244_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G211gat), .B(G218gat), .Z(new_n252_));
  OAI211_X1 g051(.A(new_n252_), .B(KEYINPUT21), .C1(new_n246_), .C2(new_n248_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n202_), .B1(new_n241_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT19), .Z(new_n257_));
  OAI21_X1  g056(.A(new_n224_), .B1(G183gat), .B2(G190gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT99), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n214_), .B1(new_n204_), .B2(new_n235_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n224_), .B(KEYINPUT99), .C1(G183gat), .C2(G190gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n254_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n227_), .A2(KEYINPUT97), .A3(new_n228_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT97), .B1(new_n227_), .B2(new_n228_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n230_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n209_), .A2(KEYINPUT24), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT98), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(KEYINPUT98), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n208_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n225_), .A2(new_n226_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n267_), .A2(new_n271_), .A3(new_n233_), .A4(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n263_), .A2(new_n264_), .A3(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n255_), .A2(new_n257_), .A3(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G8gat), .B(G36gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G64gat), .B(G92gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n264_), .B1(new_n263_), .B2(new_n273_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n232_), .A2(new_n264_), .A3(new_n240_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n282_), .A2(new_n202_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n257_), .B(KEYINPUT96), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n275_), .B(new_n281_), .C1(new_n284_), .C2(new_n286_), .ZN(new_n287_));
  NOR4_X1   g086(.A1(new_n282_), .A2(new_n283_), .A3(new_n202_), .A4(new_n285_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n251_), .A2(new_n253_), .A3(KEYINPUT93), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT93), .B1(new_n251_), .B2(new_n253_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(new_n273_), .A3(new_n263_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n257_), .B1(new_n292_), .B2(new_n255_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n280_), .B1(new_n288_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT104), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n287_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n263_), .A2(new_n273_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n202_), .B1(new_n297_), .B2(new_n254_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n283_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n286_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n292_), .A2(new_n255_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n257_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT104), .B1(new_n304_), .B2(new_n280_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT27), .B1(new_n296_), .B2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n286_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n275_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n280_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n287_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT90), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT90), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(G141gat), .A3(G148gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n314_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n319_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT91), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n319_), .A2(KEYINPUT91), .A3(new_n323_), .A4(new_n324_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT92), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n314_), .B(KEYINPUT3), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n316_), .A2(new_n318_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n331_), .B(new_n332_), .C1(KEYINPUT2), .C2(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n320_), .A2(new_n322_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n313_), .B1(new_n329_), .B2(new_n336_), .ZN(new_n337_));
  OAI211_X1 g136(.A(G228gat), .B(G233gat), .C1(new_n337_), .C2(new_n291_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G78gat), .B(G106gat), .Z(new_n339_));
  NAND2_X1  g138(.A1(new_n329_), .A2(new_n336_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT29), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n264_), .B1(G228gat), .B2(G233gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n338_), .A2(new_n339_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n339_), .B1(new_n338_), .B2(new_n343_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n329_), .A2(new_n336_), .A3(new_n313_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G22gat), .B(G50gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT28), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n348_), .B(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n344_), .A2(KEYINPUT94), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n338_), .A2(new_n343_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n339_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT94), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n338_), .A2(new_n343_), .A3(new_n357_), .A4(new_n339_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n353_), .A2(new_n356_), .A3(new_n351_), .A4(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT95), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n346_), .B1(KEYINPUT94), .B2(new_n344_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n358_), .A2(new_n351_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(KEYINPUT95), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n352_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n312_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n367_), .A2(G113gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(G113gat), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n368_), .A2(G120gat), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(G120gat), .B1(new_n368_), .B2(new_n369_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n340_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n370_), .A2(new_n371_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n329_), .A3(new_n336_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT101), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n373_), .A2(KEYINPUT4), .A3(new_n375_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n372_), .A2(new_n340_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n378_), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G1gat), .B(G29gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(G57gat), .B(G85gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n380_), .A2(new_n384_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n372_), .B(KEYINPUT31), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n241_), .A2(KEYINPUT30), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n241_), .A2(KEYINPUT30), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT86), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n241_), .A2(KEYINPUT30), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT86), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n241_), .A2(KEYINPUT30), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G71gat), .B(G99gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT85), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n405_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n398_), .A2(new_n402_), .A3(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(KEYINPUT86), .B(new_n408_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT87), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT88), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n395_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n395_), .A2(new_n413_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n411_), .B(new_n410_), .C1(new_n415_), .C2(KEYINPUT87), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n366_), .A2(new_n393_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n361_), .A2(new_n364_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n352_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n393_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT32), .B(new_n281_), .C1(new_n288_), .C2(new_n293_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n281_), .A2(KEYINPUT32), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n275_), .B(new_n423_), .C1(new_n284_), .C2(new_n286_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n422_), .B(new_n424_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n381_), .A2(new_n379_), .A3(new_n383_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT103), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n389_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n381_), .A2(KEYINPUT103), .A3(new_n379_), .A4(new_n383_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n287_), .A3(new_n309_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT33), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n390_), .A2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n380_), .A2(new_n384_), .A3(KEYINPUT33), .A4(new_n389_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n425_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n421_), .A2(new_n312_), .B1(new_n437_), .B2(new_n365_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n417_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n414_), .A2(KEYINPUT89), .A3(new_n416_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT105), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT105), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n441_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n309_), .A2(new_n310_), .A3(new_n287_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n294_), .A2(new_n295_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n304_), .A2(KEYINPUT104), .A3(new_n280_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n287_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n446_), .B1(new_n449_), .B2(KEYINPUT27), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n450_), .A2(new_n393_), .A3(new_n365_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n437_), .A2(new_n365_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n444_), .B(new_n445_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n418_), .B1(new_n443_), .B2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(G229gat), .A2(G233gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT77), .ZN(new_n456_));
  AND2_X1   g255(.A1(G29gat), .A2(G36gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G29gat), .A2(G36gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(G43gat), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(G29gat), .ZN(new_n460_));
  INV_X1    g259(.A(G36gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G43gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G29gat), .A2(G36gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n459_), .A2(new_n465_), .A3(G50gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(G50gat), .B1(new_n459_), .B2(new_n465_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT14), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT72), .B(G1gat), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n469_), .B1(new_n470_), .B2(G8gat), .ZN(new_n471_));
  INV_X1    g270(.A(G15gat), .ZN(new_n472_));
  INV_X1    g271(.A(G22gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G15gat), .A2(G22gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G1gat), .B(G8gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n471_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n476_), .ZN(new_n480_));
  INV_X1    g279(.A(G1gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT72), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT72), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G1gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n484_), .A3(G8gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT14), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n477_), .B1(new_n480_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n468_), .B1(new_n479_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT76), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n478_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n480_), .A2(new_n486_), .A3(new_n477_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT76), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n468_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n492_), .A2(new_n468_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n456_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  AOI211_X1 g297(.A(KEYINPUT77), .B(new_n496_), .C1(new_n489_), .C2(new_n494_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n455_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT78), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n468_), .B(KEYINPUT15), .ZN(new_n502_));
  INV_X1    g301(.A(new_n492_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(new_n495_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT78), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n507_), .B(new_n455_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n501_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(new_n203_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(new_n245_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n501_), .A2(new_n506_), .A3(new_n508_), .A4(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(KEYINPUT79), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT79), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n509_), .A2(new_n517_), .A3(new_n512_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G190gat), .B(G218gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G134gat), .ZN(new_n522_));
  INV_X1    g321(.A(G162gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT36), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT10), .B(G99gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT64), .B(G106gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(G85gat), .A2(G92gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT9), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT65), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT9), .ZN(new_n537_));
  INV_X1    g336(.A(G85gat), .ZN(new_n538_));
  INV_X1    g337(.A(G92gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n535_), .A2(new_n536_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n536_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n529_), .B(new_n532_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(G99gat), .ZN(new_n544_));
  INV_X1    g343(.A(G106gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(KEYINPUT66), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT7), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n548_), .A2(new_n544_), .A3(new_n545_), .A4(KEYINPUT66), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n532_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n533_), .A2(new_n534_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT67), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT8), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n550_), .A2(new_n553_), .A3(KEYINPUT8), .A4(new_n551_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n543_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n502_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT70), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT34), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT35), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n543_), .A2(new_n555_), .A3(new_n468_), .A4(new_n556_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n558_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n561_), .A2(new_n562_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n526_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n524_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n570_), .A2(KEYINPUT36), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(new_n571_), .A3(new_n568_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n567_), .A2(KEYINPUT71), .A3(new_n571_), .A4(new_n568_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n569_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT37), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G57gat), .B(G64gat), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT11), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT11), .ZN(new_n581_));
  XOR2_X1   g380(.A(G71gat), .B(G78gat), .Z(new_n582_));
  NAND3_X1  g381(.A1(new_n580_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n557_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n585_), .A2(new_n543_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(KEYINPUT12), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n557_), .A2(new_n590_), .A3(new_n586_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n587_), .A2(new_n588_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n594_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(G120gat), .B(G148gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n596_), .B(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n603_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n503_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n492_), .A2(G231gat), .A3(G233gat), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n585_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n585_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT16), .B(G183gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G127gat), .B(G155gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  OAI22_X1  g420(.A1(new_n612_), .A2(new_n613_), .B1(new_n619_), .B2(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT73), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n623_), .A2(KEYINPUT73), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT74), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT74), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n578_), .A2(new_n608_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT75), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n520_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  AOI211_X1 g434(.A(new_n454_), .B(new_n635_), .C1(new_n634_), .C2(new_n633_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n470_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n393_), .A3(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT38), .ZN(new_n639_));
  INV_X1    g438(.A(new_n418_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n438_), .A2(new_n442_), .A3(KEYINPUT105), .ZN(new_n641_));
  INV_X1    g440(.A(new_n393_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n359_), .A2(new_n360_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT95), .B1(new_n362_), .B2(new_n363_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n420_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n312_), .A2(new_n642_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n437_), .A2(new_n365_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n444_), .B1(new_n648_), .B2(new_n445_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n640_), .B1(new_n641_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT108), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n576_), .B(KEYINPUT107), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n651_), .A3(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT108), .B1(new_n454_), .B2(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n520_), .A2(new_n608_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n627_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT106), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n656_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n642_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n639_), .A2(new_n662_), .ZN(G1324gat));
  INV_X1    g462(.A(G8gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n636_), .A2(new_n664_), .A3(new_n450_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n656_), .A2(new_n450_), .A3(new_n660_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(G8gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n666_), .B2(G8gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n671_), .B(new_n665_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1325gat));
  NAND3_X1  g474(.A1(new_n636_), .A2(new_n472_), .A3(new_n442_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n656_), .A2(new_n442_), .A3(new_n660_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n677_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT41), .B1(new_n677_), .B2(G15gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT110), .B(new_n676_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1326gat));
  NAND3_X1  g483(.A1(new_n636_), .A2(new_n473_), .A3(new_n645_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G22gat), .B1(new_n661_), .B2(new_n365_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(KEYINPUT42), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(KEYINPUT42), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n685_), .B1(new_n687_), .B2(new_n688_), .ZN(G1327gat));
  NAND2_X1  g488(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n650_), .A2(new_n577_), .A3(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(new_n454_), .B2(new_n578_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n520_), .A2(new_n608_), .A3(new_n631_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n692_), .A2(new_n695_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n692_), .A2(new_n695_), .A3(KEYINPUT44), .A4(new_n697_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n700_), .A2(G29gat), .A3(new_n393_), .A4(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n574_), .A2(new_n575_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n569_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n454_), .A2(new_n696_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n460_), .B1(new_n707_), .B2(new_n642_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n702_), .A2(new_n708_), .ZN(G1328gat));
  NAND2_X1  g508(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n700_), .A2(new_n450_), .A3(new_n701_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G36gat), .ZN(new_n712_));
  OR2_X1    g511(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n650_), .A2(new_n461_), .A3(new_n576_), .A4(new_n697_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT45), .B1(new_n714_), .B2(new_n312_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n706_), .A2(new_n716_), .A3(new_n461_), .A4(new_n450_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AND4_X1   g518(.A1(new_n710_), .A2(new_n712_), .A3(new_n713_), .A4(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n718_), .B1(new_n711_), .B2(G36gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n710_), .B1(new_n721_), .B2(new_n713_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1329gat));
  INV_X1    g522(.A(new_n417_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n700_), .A2(G43gat), .A3(new_n724_), .A4(new_n701_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n463_), .B1(new_n707_), .B2(new_n445_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n706_), .B2(new_n645_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n700_), .A2(new_n645_), .A3(new_n701_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(G50gat), .ZN(G1331gat));
  NOR2_X1   g530(.A1(new_n520_), .A2(new_n608_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n632_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n454_), .A2(new_n577_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n393_), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n642_), .B(new_n733_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g536(.A(G64gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n734_), .A2(new_n738_), .A3(new_n450_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n733_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n656_), .A2(new_n450_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G64gat), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(KEYINPUT48), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(KEYINPUT48), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n739_), .B1(new_n743_), .B2(new_n744_), .ZN(G1333gat));
  NOR2_X1   g544(.A1(new_n445_), .A2(G71gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT114), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n734_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n656_), .A2(new_n442_), .A3(new_n740_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G71gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT113), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n752_), .A3(G71gat), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n751_), .A2(KEYINPUT49), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT49), .B1(new_n751_), .B2(new_n753_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n748_), .B1(new_n754_), .B2(new_n755_), .ZN(G1334gat));
  INV_X1    g555(.A(G78gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n734_), .A2(new_n757_), .A3(new_n645_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n656_), .A2(new_n645_), .A3(new_n740_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(G78gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT115), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n762_), .A3(G78gat), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n761_), .A2(KEYINPUT50), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT50), .B1(new_n761_), .B2(new_n763_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n758_), .B1(new_n764_), .B2(new_n765_), .ZN(G1335gat));
  NOR3_X1   g565(.A1(new_n632_), .A2(new_n520_), .A3(new_n608_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n650_), .A2(new_n576_), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n393_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT116), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n692_), .A2(new_n695_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n767_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n393_), .A2(G85gat), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT117), .Z(new_n775_));
  AOI21_X1  g574(.A(new_n770_), .B1(new_n773_), .B2(new_n775_), .ZN(G1336gat));
  AOI21_X1  g575(.A(G92gat), .B1(new_n768_), .B2(new_n450_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n772_), .A2(new_n539_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n450_), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n772_), .B2(new_n445_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n768_), .A2(new_n527_), .A3(new_n724_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n768_), .A2(new_n528_), .A3(new_n645_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n692_), .A2(new_n695_), .A3(new_n645_), .A4(new_n767_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(G106gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n785_), .B2(G106gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  XOR2_X1   g588(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1339gat));
  NOR2_X1   g590(.A1(new_n577_), .A2(new_n631_), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n792_), .A2(new_n519_), .A3(new_n608_), .A4(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT120), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n793_), .B1(new_n633_), .B2(new_n520_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n605_), .A2(new_n607_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n798_), .A2(new_n577_), .A3(new_n631_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n799_), .A2(new_n800_), .A3(new_n519_), .A4(new_n794_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n796_), .A2(new_n797_), .A3(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n596_), .A2(new_n602_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n593_), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT55), .B(new_n806_), .C1(new_n589_), .C2(new_n591_), .ZN(new_n807_));
  OAI22_X1  g606(.A1(new_n805_), .A2(new_n807_), .B1(new_n593_), .B2(new_n592_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n602_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT122), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n803_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n498_), .A2(new_n499_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n512_), .B1(new_n813_), .B2(new_n455_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT121), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n504_), .A2(new_n455_), .A3(new_n495_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n817_), .B(new_n512_), .C1(new_n813_), .C2(new_n455_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(new_n515_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n592_), .A2(new_n593_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n594_), .A2(KEYINPUT55), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n592_), .A2(new_n804_), .A3(new_n593_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n821_), .B1(new_n825_), .B2(new_n601_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(KEYINPUT122), .A3(new_n809_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n812_), .A2(new_n820_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n812_), .A2(new_n820_), .A3(new_n827_), .A4(KEYINPUT58), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n577_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n803_), .B1(new_n826_), .B2(new_n809_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n518_), .A3(new_n516_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n819_), .A2(new_n603_), .A3(new_n515_), .ZN(new_n835_));
  AOI211_X1 g634(.A(KEYINPUT57), .B(new_n576_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  INV_X1    g636(.A(new_n803_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT56), .B1(new_n808_), .B2(new_n602_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n810_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n835_), .B1(new_n519_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n837_), .B1(new_n841_), .B2(new_n705_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n832_), .B1(new_n836_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n631_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n802_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n366_), .A2(new_n642_), .A3(new_n417_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n847_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n843_), .A2(KEYINPUT123), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n851_), .B(new_n832_), .C1(new_n836_), .C2(new_n842_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n658_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n849_), .B1(new_n853_), .B2(new_n802_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n848_), .B1(new_n854_), .B2(new_n846_), .ZN(new_n855_));
  INV_X1    g654(.A(G113gat), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n519_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n796_), .A2(new_n801_), .A3(new_n797_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n627_), .B1(new_n843_), .B2(KEYINPUT123), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n852_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n861_), .B2(new_n849_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n854_), .A2(KEYINPUT124), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n520_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n857_), .B1(new_n856_), .B2(new_n865_), .ZN(G1340gat));
  INV_X1    g665(.A(G120gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n608_), .B2(KEYINPUT60), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n864_), .B(new_n868_), .C1(KEYINPUT60), .C2(new_n867_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G120gat), .B1(new_n855_), .B2(new_n608_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1341gat));
  INV_X1    g670(.A(G127gat), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n855_), .A2(new_n872_), .A3(new_n658_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n864_), .A2(new_n632_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n872_), .B2(new_n874_), .ZN(G1342gat));
  INV_X1    g674(.A(G134gat), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n855_), .A2(new_n876_), .A3(new_n578_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n864_), .A2(new_n652_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n876_), .B2(new_n878_), .ZN(G1343gat));
  NOR2_X1   g678(.A1(new_n442_), .A2(new_n365_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n853_), .B2(new_n802_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n450_), .A2(new_n642_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(new_n520_), .A3(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g684(.A1(new_n882_), .A2(new_n798_), .A3(new_n883_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g686(.A1(new_n882_), .A2(new_n883_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n631_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT61), .B(G155gat), .Z(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1346gat));
  NOR3_X1   g690(.A1(new_n888_), .A2(new_n523_), .A3(new_n578_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n882_), .A2(new_n652_), .A3(new_n883_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n523_), .B2(new_n893_), .ZN(G1347gat));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n645_), .B1(new_n802_), .B2(new_n844_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n312_), .A2(new_n393_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n445_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n519_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n895_), .B1(new_n901_), .B2(new_n203_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n235_), .ZN(new_n903_));
  OAI211_X1 g702(.A(KEYINPUT62), .B(G169gat), .C1(new_n900_), .C2(new_n519_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(G1348gat));
  INV_X1    g704(.A(new_n900_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G176gat), .B1(new_n906_), .B2(new_n798_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n861_), .A2(new_n645_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n899_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n909_), .A2(new_n204_), .A3(new_n608_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n907_), .B1(new_n908_), .B2(new_n910_), .ZN(G1349gat));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n645_), .B(new_n909_), .C1(new_n853_), .C2(new_n802_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G183gat), .B1(new_n913_), .B2(new_n632_), .ZN(new_n914_));
  NOR4_X1   g713(.A1(new_n900_), .A2(new_n266_), .A3(new_n265_), .A4(new_n658_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n912_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n265_), .A2(new_n266_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n906_), .A2(new_n917_), .A3(new_n627_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n861_), .A2(new_n645_), .A3(new_n631_), .A4(new_n909_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n918_), .B(KEYINPUT125), .C1(new_n919_), .C2(G183gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n916_), .A2(new_n920_), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n900_), .B2(new_n578_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n652_), .A2(new_n230_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n900_), .B2(new_n923_), .ZN(G1351gat));
  NOR3_X1   g723(.A1(new_n861_), .A2(new_n881_), .A3(new_n898_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n520_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n798_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g728(.A1(new_n853_), .A2(new_n802_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n658_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n930_), .A2(new_n880_), .A3(new_n897_), .A4(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT126), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n882_), .A2(new_n935_), .A3(new_n897_), .A4(new_n931_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n933_), .A2(new_n934_), .A3(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n934_), .B1(new_n933_), .B2(new_n936_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1354gat));
  AOI21_X1  g738(.A(G218gat), .B1(new_n925_), .B2(new_n652_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n577_), .A2(G218gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT127), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n925_), .B2(new_n942_), .ZN(G1355gat));
endmodule


