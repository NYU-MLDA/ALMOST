//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n202_), .B(new_n203_), .C1(new_n206_), .C2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n204_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(new_n203_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n211_), .B(new_n207_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT29), .ZN(new_n217_));
  XOR2_X1   g016(.A(G22gat), .B(G50gat), .Z(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n219_), .A2(new_n221_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n216_), .A2(KEYINPUT29), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G211gat), .B(G218gat), .ZN(new_n227_));
  INV_X1    g026(.A(G204gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(G197gat), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n227_), .B(KEYINPUT21), .C1(KEYINPUT92), .C2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G197gat), .B(G204gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n227_), .A2(KEYINPUT21), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n229_), .A2(KEYINPUT92), .ZN(new_n234_));
  INV_X1    g033(.A(new_n231_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT21), .A4(new_n227_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT91), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT93), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n226_), .A2(new_n238_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n226_), .A2(new_n238_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n241_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G78gat), .B(G106gat), .Z(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n247_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n225_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT94), .B1(new_n246_), .B2(new_n247_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n249_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT90), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n224_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n222_), .A3(KEYINPUT90), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n251_), .B1(new_n253_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G183gat), .A2(G190gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT23), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n263_), .B(new_n264_), .C1(G183gat), .C2(G190gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT22), .B(G169gat), .Z(new_n267_));
  OAI211_X1 g066(.A(new_n265_), .B(new_n266_), .C1(G176gat), .C2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n270_));
  AND2_X1   g069(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n272_));
  OAI22_X1  g071(.A1(new_n269_), .A2(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT83), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT25), .B(G183gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G190gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT24), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT84), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n281_), .A2(G169gat), .A3(G176gat), .ZN(new_n282_));
  INV_X1    g081(.A(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT84), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n280_), .B1(new_n282_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n263_), .A2(new_n264_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT84), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n281_), .B1(G169gat), .B2(G176gat), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(KEYINPUT24), .A4(new_n266_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n268_), .B1(new_n279_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT85), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(KEYINPUT85), .B(new_n268_), .C1(new_n279_), .C2(new_n292_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(new_n237_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n297_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT95), .B1(new_n297_), .B2(KEYINPUT20), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT99), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT19), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n289_), .A2(new_n290_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n287_), .B1(new_n280_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(new_n291_), .A3(new_n273_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n268_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(new_n237_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n300_), .A2(new_n301_), .A3(new_n304_), .A4(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT95), .ZN(new_n313_));
  INV_X1    g112(.A(new_n296_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n306_), .A2(new_n291_), .A3(new_n274_), .A4(new_n278_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT85), .B1(new_n315_), .B2(new_n268_), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n314_), .A2(new_n316_), .A3(new_n238_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT20), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n313_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n297_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n319_), .A2(new_n304_), .A3(new_n311_), .A4(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT99), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n308_), .A2(KEYINPUT98), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n308_), .A2(KEYINPUT98), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n237_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n295_), .A2(new_n296_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n238_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n327_), .A3(KEYINPUT20), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n303_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n312_), .A2(new_n322_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT100), .ZN(new_n331_));
  XOR2_X1   g130(.A(G8gat), .B(G36gat), .Z(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G92gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT18), .B(G64gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT32), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n330_), .A2(new_n331_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n331_), .B1(new_n330_), .B2(new_n337_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n318_), .B1(new_n309_), .B2(new_n237_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n327_), .A2(new_n304_), .A3(new_n340_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n298_), .A2(new_n299_), .A3(new_n310_), .ZN(new_n342_));
  OAI221_X1 g141(.A(new_n341_), .B1(new_n336_), .B2(new_n335_), .C1(new_n342_), .C2(new_n304_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT0), .B(G57gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(G127gat), .B(G134gat), .Z(new_n350_));
  XNOR2_X1  g149(.A(G113gat), .B(G120gat), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n351_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n216_), .A2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(KEYINPUT4), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT96), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n210_), .A2(new_n353_), .A3(new_n352_), .A4(new_n215_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  OR3_X1    g158(.A1(new_n216_), .A2(new_n357_), .A3(new_n354_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AOI211_X1 g160(.A(new_n349_), .B(new_n356_), .C1(new_n361_), .C2(KEYINPUT4), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n349_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n348_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n356_), .B1(new_n361_), .B2(KEYINPUT4), .ZN(new_n366_));
  INV_X1    g165(.A(new_n349_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n363_), .A3(new_n347_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n343_), .A2(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n338_), .A2(new_n339_), .A3(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n341_), .B1(new_n342_), .B2(new_n304_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n335_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n369_), .B1(KEYINPUT97), .B2(KEYINPUT33), .ZN(new_n375_));
  NOR2_X1   g174(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n368_), .A2(new_n363_), .A3(new_n347_), .A4(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n373_), .A2(new_n335_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n347_), .B1(new_n366_), .B2(new_n349_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n361_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n349_), .B2(new_n381_), .ZN(new_n382_));
  AND4_X1   g181(.A1(new_n374_), .A2(new_n378_), .A3(new_n379_), .A4(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n260_), .B1(new_n372_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT101), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n260_), .A2(new_n370_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n330_), .A2(new_n335_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n379_), .A3(KEYINPUT27), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT102), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n379_), .A2(new_n374_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT27), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT102), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n387_), .A2(new_n379_), .A3(new_n393_), .A4(KEYINPUT27), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n386_), .A2(new_n389_), .A3(new_n392_), .A4(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n330_), .A2(new_n337_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT100), .ZN(new_n397_));
  INV_X1    g196(.A(new_n371_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n330_), .A2(new_n331_), .A3(new_n337_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n378_), .A2(new_n379_), .A3(new_n374_), .A4(new_n382_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT101), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n260_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n385_), .A2(new_n395_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT31), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n326_), .B(new_n409_), .Z(new_n410_));
  XNOR2_X1  g209(.A(G71gat), .B(G99gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G15gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n354_), .B(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(KEYINPUT86), .B(G43gat), .Z(new_n414_));
  XOR2_X1   g213(.A(new_n413_), .B(new_n414_), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n410_), .B(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n416_), .B(KEYINPUT88), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT103), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n389_), .A2(new_n416_), .A3(new_n392_), .A4(new_n394_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n259_), .A2(new_n370_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n389_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n424_), .A2(KEYINPUT103), .A3(new_n416_), .A4(new_n421_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n405_), .A2(new_n418_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G15gat), .B(G22gat), .ZN(new_n427_));
  INV_X1    g226(.A(G1gat), .ZN(new_n428_));
  INV_X1    g227(.A(G8gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT14), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G1gat), .B(G8gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G29gat), .B(G36gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G50gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT71), .B(G43gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n439_), .B(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n441_), .B1(new_n444_), .B2(new_n435_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G229gat), .A2(G233gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT81), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT81), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n435_), .B(new_n440_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(new_n447_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n449_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G113gat), .B(G141gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G169gat), .B(G197gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n453_), .B(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n458_), .B(KEYINPUT82), .Z(new_n459_));
  OR3_X1    g258(.A1(new_n426_), .A2(KEYINPUT104), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT66), .ZN(new_n461_));
  INV_X1    g260(.A(G99gat), .ZN(new_n462_));
  INV_X1    g261(.A(G106gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n464_), .A2(KEYINPUT7), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT6), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(KEYINPUT7), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G85gat), .B(G92gat), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT8), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT10), .B(G99gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n463_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(KEYINPUT9), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n477_), .A2(KEYINPUT9), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n475_), .A2(new_n476_), .A3(new_n478_), .A4(new_n467_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT65), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n472_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G57gat), .B(G64gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT11), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(KEYINPUT11), .ZN(new_n484_));
  XOR2_X1   g283(.A(G71gat), .B(G78gat), .Z(new_n485_));
  MUX2_X1   g284(.A(new_n483_), .B(new_n484_), .S(new_n485_), .Z(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT12), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n486_), .B(KEYINPUT67), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(KEYINPUT12), .A3(new_n481_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n481_), .A2(new_n486_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n489_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G230gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT64), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n492_), .A2(new_n487_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n497_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G120gat), .B(G148gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT69), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G176gat), .B(G204gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT70), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n499_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n505_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n499_), .A2(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT13), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  OR3_X1    g311(.A1(new_n507_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT104), .B1(new_n426_), .B2(new_n459_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n460_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT37), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT34), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n439_), .B(new_n442_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n521_), .A2(new_n481_), .ZN(new_n522_));
  OAI211_X1 g321(.A(KEYINPUT35), .B(new_n520_), .C1(new_n522_), .C2(KEYINPUT73), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n481_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(new_n439_), .B2(new_n481_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n525_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n520_), .A2(KEYINPUT35), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G190gat), .B(G218gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(KEYINPUT36), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n526_), .A2(new_n528_), .A3(new_n527_), .A4(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n518_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n529_), .A2(KEYINPUT74), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n526_), .A2(new_n527_), .A3(new_n539_), .A4(new_n528_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(new_n518_), .A3(new_n534_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n541_), .A2(KEYINPUT75), .A3(new_n518_), .A4(new_n534_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n537_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n435_), .B(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n486_), .B(KEYINPUT80), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n551_));
  XNOR2_X1  g350(.A(G127gat), .B(G155gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G183gat), .B(G211gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n555_), .A2(new_n556_), .ZN(new_n558_));
  OR3_X1    g357(.A1(new_n550_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n548_), .A2(new_n490_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n548_), .A2(new_n490_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n562_), .A2(KEYINPUT79), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(KEYINPUT79), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n546_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n517_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n370_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n567_), .A2(G1gat), .A3(new_n568_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n569_), .A2(KEYINPUT38), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(KEYINPUT38), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n514_), .A2(new_n459_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n541_), .A2(new_n534_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n565_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n426_), .A2(new_n575_), .A3(new_n568_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n570_), .B(new_n571_), .C1(new_n428_), .C2(new_n576_), .ZN(G1324gat));
  NOR3_X1   g376(.A1(new_n426_), .A2(new_n575_), .A3(new_n424_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT105), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(G8gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT39), .ZN(new_n581_));
  INV_X1    g380(.A(new_n424_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n517_), .A2(new_n429_), .A3(new_n582_), .A4(new_n566_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT40), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n581_), .A2(KEYINPUT40), .A3(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(G1325gat));
  INV_X1    g387(.A(G15gat), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n426_), .A2(new_n575_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n590_), .B2(new_n417_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT41), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n417_), .A2(new_n589_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n592_), .B1(new_n567_), .B2(new_n593_), .ZN(G1326gat));
  INV_X1    g393(.A(G22gat), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n590_), .B2(new_n259_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT42), .Z(new_n597_));
  NAND2_X1  g396(.A1(new_n259_), .A2(new_n595_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n567_), .B2(new_n598_), .ZN(G1327gat));
  INV_X1    g398(.A(new_n573_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n565_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AND4_X1   g401(.A1(new_n515_), .A2(new_n460_), .A3(new_n516_), .A4(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n604_), .A2(G29gat), .A3(new_n568_), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n544_), .A2(new_n545_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n537_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT43), .B1(new_n426_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT43), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n403_), .B1(new_n402_), .B2(new_n260_), .ZN(new_n613_));
  AOI211_X1 g412(.A(KEYINPUT101), .B(new_n259_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n417_), .B1(new_n615_), .B2(new_n395_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n425_), .A2(new_n423_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n612_), .B(new_n546_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n611_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n572_), .A2(new_n565_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n607_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI211_X1 g423(.A(new_n620_), .B(new_n624_), .C1(new_n611_), .C2(new_n618_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G29gat), .B1(new_n626_), .B2(new_n568_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n605_), .A2(new_n627_), .ZN(G1328gat));
  OAI21_X1  g427(.A(G36gat), .B1(new_n626_), .B2(new_n424_), .ZN(new_n629_));
  INV_X1    g428(.A(G36gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n603_), .A2(new_n630_), .A3(new_n582_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n603_), .A2(new_n630_), .A3(new_n582_), .A4(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n629_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT46), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1329gat));
  INV_X1    g437(.A(G43gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n604_), .B2(new_n418_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT108), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n405_), .A2(new_n418_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n425_), .A2(new_n423_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n612_), .B1(new_n644_), .B2(new_n546_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n426_), .A2(KEYINPUT43), .A3(new_n610_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n621_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n606_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n621_), .B(new_n623_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n639_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n641_), .B1(new_n650_), .B2(new_n416_), .ZN(new_n651_));
  OAI211_X1 g450(.A(G43gat), .B(new_n416_), .C1(new_n622_), .C2(new_n625_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(KEYINPUT108), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n640_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT47), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT47), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n656_), .B(new_n640_), .C1(new_n651_), .C2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1330gat));
  INV_X1    g457(.A(G50gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n603_), .A2(new_n659_), .A3(new_n259_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n620_), .B1(new_n611_), .B2(new_n618_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n649_), .B1(new_n661_), .B2(new_n607_), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT109), .B(new_n659_), .C1(new_n662_), .C2(new_n259_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT109), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n259_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(G50gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n660_), .B1(new_n663_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT110), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT110), .B(new_n660_), .C1(new_n663_), .C2(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1331gat));
  INV_X1    g470(.A(G57gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n514_), .A2(new_n459_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n426_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n566_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n675_), .B2(new_n568_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT111), .Z(new_n677_));
  AND2_X1   g476(.A1(new_n674_), .A2(new_n574_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n568_), .A2(new_n672_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(new_n678_), .B2(new_n679_), .ZN(G1332gat));
  INV_X1    g479(.A(G64gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n678_), .B2(new_n582_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT48), .Z(new_n683_));
  INV_X1    g482(.A(new_n675_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n681_), .A3(new_n582_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1333gat));
  INV_X1    g485(.A(G71gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n678_), .B2(new_n417_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT49), .Z(new_n689_));
  NAND3_X1  g488(.A1(new_n684_), .A2(new_n687_), .A3(new_n417_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1334gat));
  NAND2_X1  g490(.A1(new_n678_), .A2(new_n259_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT113), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(G78gat), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n692_), .B2(G78gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT112), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n696_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT112), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n694_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT50), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OR3_X1    g502(.A1(new_n675_), .A2(G78gat), .A3(new_n260_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n697_), .A2(new_n700_), .A3(KEYINPUT50), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(G1335gat));
  AND2_X1   g505(.A1(new_n674_), .A2(new_n602_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G85gat), .B1(new_n707_), .B2(new_n370_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n673_), .B1(new_n611_), .B2(new_n618_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n565_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(new_n568_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n711_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g511(.A(G92gat), .B1(new_n707_), .B2(new_n582_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n710_), .A2(new_n424_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(G92gat), .ZN(G1337gat));
  NAND3_X1  g514(.A1(new_n707_), .A2(new_n416_), .A3(new_n474_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT114), .Z(new_n717_));
  OAI21_X1  g516(.A(G99gat), .B1(new_n710_), .B2(new_n418_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g519(.A1(new_n707_), .A2(new_n463_), .A3(new_n259_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n709_), .A2(new_n259_), .A3(new_n565_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G106gat), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(KEYINPUT52), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(KEYINPUT52), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n721_), .B(new_n722_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n724_), .B(KEYINPUT52), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n722_), .B1(new_n729_), .B2(new_n721_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1339gat));
  INV_X1    g530(.A(KEYINPUT117), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n497_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n497_), .B2(new_n732_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n493_), .A2(new_n496_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n734_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n506_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT56), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n509_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n453_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n445_), .A2(new_n446_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n457_), .B1(new_n451_), .B2(new_n446_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT118), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n742_), .A2(new_n457_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n497_), .A2(new_n732_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT55), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n497_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n736_), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n506_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n740_), .A2(new_n741_), .A3(new_n746_), .A4(new_n752_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT119), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT58), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n753_), .B2(KEYINPUT119), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n546_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT120), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n753_), .A2(new_n755_), .ZN(new_n760_));
  OAI211_X1 g559(.A(KEYINPUT120), .B(new_n546_), .C1(new_n754_), .C2(new_n756_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n458_), .B(KEYINPUT82), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n763_), .A2(new_n741_), .A3(new_n752_), .A4(new_n740_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n510_), .A2(new_n746_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n573_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT57), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n601_), .B1(new_n762_), .B2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n610_), .A2(new_n459_), .A3(new_n515_), .A4(new_n601_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT116), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n566_), .A2(new_n772_), .A3(new_n459_), .A4(new_n515_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(KEYINPUT54), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n770_), .A2(KEYINPUT116), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n370_), .B(new_n260_), .C1(new_n769_), .C2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(new_n420_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n763_), .ZN(new_n780_));
  INV_X1    g579(.A(G113gat), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n762_), .A2(new_n768_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n565_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n774_), .A2(new_n776_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n259_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT59), .ZN(new_n787_));
  INV_X1    g586(.A(new_n420_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n370_), .A4(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT59), .B1(new_n778_), .B2(new_n420_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(G113gat), .A4(new_n763_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n782_), .A2(new_n791_), .ZN(G1340gat));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n790_), .A3(new_n514_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(G120gat), .ZN(new_n794_));
  INV_X1    g593(.A(G120gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n515_), .B2(KEYINPUT60), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n779_), .B(new_n796_), .C1(KEYINPUT60), .C2(new_n795_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(G1341gat));
  AOI21_X1  g597(.A(G127gat), .B1(new_n779_), .B2(new_n601_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n789_), .A2(new_n790_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n601_), .A2(G127gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(G1342gat));
  AOI21_X1  g601(.A(G134gat), .B1(new_n779_), .B2(new_n573_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n546_), .A2(G134gat), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(KEYINPUT121), .Z(new_n805_));
  AOI21_X1  g604(.A(new_n803_), .B1(new_n800_), .B2(new_n805_), .ZN(G1343gat));
  NOR3_X1   g605(.A1(new_n582_), .A2(new_n568_), .A3(new_n260_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n418_), .B(new_n807_), .C1(new_n769_), .C2(new_n777_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(new_n459_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n515_), .ZN(new_n811_));
  XOR2_X1   g610(.A(new_n811_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g611(.A1(new_n808_), .A2(new_n565_), .ZN(new_n813_));
  XOR2_X1   g612(.A(KEYINPUT61), .B(G155gat), .Z(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(G1346gat));
  INV_X1    g614(.A(G162gat), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n808_), .A2(new_n816_), .A3(new_n610_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n808_), .B2(new_n600_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n818_), .A2(KEYINPUT122), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(KEYINPUT122), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n817_), .B1(new_n819_), .B2(new_n820_), .ZN(G1347gat));
  NOR2_X1   g620(.A1(new_n424_), .A2(new_n370_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n786_), .A2(new_n417_), .A3(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT62), .B(G169gat), .C1(new_n823_), .C2(new_n459_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT62), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n417_), .B(new_n260_), .C1(new_n769_), .C2(new_n777_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n822_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n826_), .A2(new_n459_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n825_), .B1(new_n828_), .B2(new_n283_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n828_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n824_), .B(new_n829_), .C1(new_n267_), .C2(new_n830_), .ZN(G1348gat));
  XOR2_X1   g630(.A(KEYINPUT123), .B(G176gat), .Z(new_n832_));
  NOR3_X1   g631(.A1(new_n823_), .A2(new_n515_), .A3(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n826_), .A2(new_n827_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n514_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(KEYINPUT123), .A2(G176gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n833_), .B1(new_n835_), .B2(new_n836_), .ZN(G1349gat));
  OAI21_X1  g636(.A(G183gat), .B1(new_n823_), .B2(new_n565_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n834_), .A2(new_n275_), .A3(new_n601_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1350gat));
  OAI21_X1  g639(.A(G190gat), .B1(new_n823_), .B2(new_n610_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n834_), .A2(new_n276_), .A3(new_n573_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1351gat));
  OAI211_X1 g642(.A(new_n418_), .B(new_n259_), .C1(new_n769_), .C2(new_n777_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n827_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n763_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g646(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(new_n514_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT125), .B1(new_n850_), .B2(G204gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT126), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n845_), .A2(new_n514_), .A3(new_n848_), .A4(new_n852_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1353gat));
  NOR3_X1   g655(.A1(new_n844_), .A2(new_n565_), .A3(new_n827_), .ZN(new_n857_));
  OR2_X1    g656(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT63), .B(G211gat), .Z(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n857_), .B2(new_n860_), .ZN(G1354gat));
  XOR2_X1   g660(.A(KEYINPUT127), .B(G218gat), .Z(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n845_), .B2(new_n573_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n845_), .A2(new_n862_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n546_), .B2(new_n864_), .ZN(G1355gat));
endmodule


