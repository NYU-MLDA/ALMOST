//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n839_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(G1gat), .A2(G8gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(KEYINPUT14), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT80), .ZN(new_n205_));
  XOR2_X1   g004(.A(G1gat), .B(G8gat), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n205_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G29gat), .B(G36gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n211_), .A2(new_n212_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n210_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n211_), .A2(new_n212_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(new_n209_), .A3(new_n213_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n208_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n205_), .B(new_n206_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n216_), .A2(KEYINPUT15), .A3(new_n218_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT15), .B1(new_n216_), .B2(new_n218_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n221_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n222_), .A2(new_n219_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n221_), .B2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G141gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G169gat), .B(G197gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G176gat), .ZN(new_n243_));
  INV_X1    g042(.A(G169gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT92), .B1(new_n244_), .B2(KEYINPUT22), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G169gat), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n243_), .B(new_n245_), .C1(new_n246_), .C2(KEYINPUT92), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT23), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT23), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(G183gat), .A3(G190gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G183gat), .ZN(new_n254_));
  INV_X1    g053(.A(G190gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n247_), .A2(new_n248_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT90), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n251_), .A2(KEYINPUT90), .A3(G183gat), .A4(G190gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT89), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n249_), .A2(new_n262_), .A3(KEYINPUT23), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n249_), .B2(KEYINPUT23), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n260_), .B(new_n261_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT91), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT88), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(new_n244_), .A3(new_n243_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT88), .B1(G169gat), .B2(G176gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(new_n266_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n255_), .A2(KEYINPUT26), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT25), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(G183gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n254_), .A2(KEYINPUT25), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT86), .ZN(new_n279_));
  OR3_X1    g078(.A1(new_n275_), .A2(KEYINPUT86), .A3(G183gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n277_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G190gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT87), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n268_), .A2(KEYINPUT24), .A3(new_n269_), .A4(new_n248_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n273_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n266_), .B1(new_n265_), .B2(new_n272_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n258_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G71gat), .B(G99gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(G43gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n289_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G113gat), .B(G120gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G134gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G127gat), .ZN(new_n296_));
  INV_X1    g095(.A(G127gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G134gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n298_), .A3(KEYINPUT95), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT95), .B1(new_n296_), .B2(new_n298_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n294_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n298_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT95), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(new_n299_), .A3(new_n293_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n302_), .A2(new_n306_), .A3(KEYINPUT96), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT96), .B1(new_n302_), .B2(new_n306_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n292_), .B(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT94), .B(G15gat), .Z(new_n311_));
  NAND2_X1  g110(.A1(G227gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT93), .B(KEYINPUT30), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT97), .B(KEYINPUT31), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n310_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n310_), .A2(new_n317_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G141gat), .ZN(new_n321_));
  INV_X1    g120(.A(G148gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT3), .ZN(new_n324_));
  OR3_X1    g123(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n324_), .A2(new_n325_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  OR2_X1    g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(KEYINPUT1), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n332_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n331_), .A2(KEYINPUT1), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n323_), .B(new_n326_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n338_), .A2(KEYINPUT29), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT28), .ZN(new_n340_));
  XOR2_X1   g139(.A(G197gat), .B(G204gat), .Z(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(KEYINPUT21), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(KEYINPUT21), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G211gat), .B(G218gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n343_), .A2(new_n344_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(KEYINPUT29), .B2(new_n338_), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n340_), .B(new_n348_), .Z(new_n349_));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT98), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G228gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G22gat), .B(G50gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n349_), .B(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G1gat), .B(G29gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT105), .B(KEYINPUT0), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G57gat), .B(G85gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OAI211_X1 g161(.A(KEYINPUT102), .B(new_n338_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n338_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(new_n306_), .A3(new_n302_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT103), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n338_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT102), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n365_), .A3(new_n363_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(KEYINPUT4), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n362_), .B(new_n372_), .C1(new_n377_), .C2(new_n368_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n345_), .A2(new_n346_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n265_), .A2(new_n256_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n246_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n248_), .B1(new_n381_), .B2(G176gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n283_), .A2(new_n278_), .A3(new_n274_), .A4(new_n276_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n286_), .A2(new_n384_), .A3(KEYINPUT99), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT99), .B1(new_n286_), .B2(new_n384_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n272_), .A2(new_n253_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n379_), .B1(new_n383_), .B2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(KEYINPUT20), .C1(new_n289_), .C2(new_n379_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT19), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT100), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n289_), .A2(new_n379_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n388_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n380_), .A2(new_n382_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n347_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n395_), .A2(KEYINPUT20), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n392_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n393_), .A2(new_n394_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT18), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  NAND2_X1  g204(.A1(new_n390_), .A2(new_n392_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT100), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n401_), .A2(KEYINPUT101), .A3(new_n405_), .A4(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n399_), .A2(new_n400_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n390_), .A2(new_n394_), .A3(new_n392_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n407_), .A2(new_n409_), .A3(new_n405_), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT101), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n407_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n405_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AND4_X1   g215(.A1(new_n378_), .A2(new_n408_), .A3(new_n413_), .A4(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT104), .ZN(new_n418_));
  INV_X1    g217(.A(new_n368_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n418_), .B1(new_n377_), .B2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n373_), .B1(new_n366_), .B2(new_n371_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT104), .B(new_n368_), .C1(new_n421_), .C2(new_n375_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT106), .B1(new_n376_), .B2(new_n368_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT106), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n366_), .A2(new_n424_), .A3(new_n419_), .A4(new_n371_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n420_), .A2(new_n422_), .A3(new_n361_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT107), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT33), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(KEYINPUT107), .A3(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n417_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n420_), .A2(new_n422_), .A3(new_n426_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n362_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n427_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n399_), .A2(new_n400_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n390_), .A2(new_n392_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT108), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n401_), .A2(new_n407_), .A3(new_n440_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT108), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n438_), .A2(new_n443_), .A3(KEYINPUT32), .A4(new_n405_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n435_), .A2(new_n441_), .A3(new_n442_), .A4(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n356_), .B1(new_n432_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n408_), .A2(new_n413_), .A3(new_n416_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT109), .B(KEYINPUT27), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT27), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(new_n438_), .B2(new_n415_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n447_), .A2(new_n449_), .B1(new_n411_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n435_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n356_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n320_), .B1(new_n446_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n452_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(new_n356_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n435_), .A2(new_n320_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n242_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT13), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G230gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G57gat), .B(G64gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT11), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT70), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n463_), .A2(KEYINPUT11), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G71gat), .B(G78gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n464_), .B(KEYINPUT70), .ZN(new_n471_));
  INV_X1    g270(.A(new_n469_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT10), .B(G99gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT64), .ZN(new_n476_));
  INV_X1    g275(.A(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(KEYINPUT65), .B(G85gat), .Z(new_n480_));
  INV_X1    g279(.A(G92gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n479_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT66), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n483_), .A2(KEYINPUT66), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT6), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n478_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT7), .ZN(new_n490_));
  INV_X1    g289(.A(G99gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n477_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n488_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT8), .ZN(new_n495_));
  XOR2_X1   g294(.A(G85gat), .B(G92gat), .Z(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n493_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT68), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT68), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n492_), .A2(new_n501_), .A3(new_n493_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n487_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(KEYINPUT67), .A2(KEYINPUT6), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n507_), .A2(G99gat), .A3(G106gat), .A4(new_n503_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n500_), .A2(new_n502_), .A3(new_n506_), .A4(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n495_), .B1(new_n509_), .B2(new_n496_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT69), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n497_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  AOI211_X1 g311(.A(KEYINPUT69), .B(new_n495_), .C1(new_n509_), .C2(new_n496_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n474_), .B(new_n489_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n462_), .B1(new_n515_), .B2(KEYINPUT71), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n489_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n474_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT71), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n514_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT72), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT12), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n517_), .A2(new_n518_), .A3(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n527_), .A2(new_n462_), .A3(new_n529_), .A4(new_n514_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G120gat), .B(G148gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G176gat), .B(G204gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n522_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n522_), .B2(new_n530_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n461_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n522_), .A2(new_n530_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n535_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n522_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(KEYINPUT13), .A3(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n220_), .B(new_n489_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT78), .B1(new_n547_), .B2(new_n548_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n502_), .A2(new_n508_), .A3(new_n506_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n501_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n496_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT8), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT69), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n510_), .A2(new_n511_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n497_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n225_), .B1(new_n559_), .B2(new_n489_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n549_), .B1(new_n552_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n226_), .A2(new_n517_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n549_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n562_), .A2(new_n563_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT76), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT36), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT77), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n561_), .A2(new_n564_), .A3(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(KEYINPUT37), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n565_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n561_), .A2(KEYINPUT79), .A3(new_n564_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n580_), .A3(new_n570_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n575_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n577_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n518_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n474_), .A2(G231gat), .A3(G233gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n222_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n208_), .A3(new_n588_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n590_), .A2(KEYINPUT81), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT81), .B1(new_n590_), .B2(new_n591_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT16), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n598_));
  NOR4_X1   g397(.A1(new_n592_), .A2(new_n593_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n597_), .B(KEYINPUT17), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n590_), .A2(new_n591_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT83), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n585_), .A2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n460_), .A2(new_n544_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(G1gat), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n435_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n582_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n539_), .A2(new_n543_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n605_), .A2(new_n614_), .A3(new_n242_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n453_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n609_), .A2(new_n610_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(new_n617_), .A3(new_n618_), .ZN(G1324gat));
  INV_X1    g418(.A(G8gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n607_), .A2(new_n620_), .A3(new_n456_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G8gat), .B1(new_n616_), .B2(new_n452_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(KEYINPUT39), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(KEYINPUT39), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n621_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g425(.A(G15gat), .B1(new_n616_), .B2(new_n320_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT41), .Z(new_n628_));
  INV_X1    g427(.A(G15gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n320_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n607_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(G1326gat));
  XOR2_X1   g431(.A(new_n356_), .B(KEYINPUT110), .Z(new_n633_));
  OAI21_X1  g432(.A(G22gat), .B1(new_n616_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(G22gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT111), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n607_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(G1327gat));
  NOR3_X1   g438(.A1(new_n614_), .A2(new_n604_), .A3(new_n582_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n460_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n435_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n614_), .A2(new_n604_), .A3(new_n242_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n455_), .A2(new_n459_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(new_n585_), .ZN(new_n647_));
  AOI211_X1 g446(.A(KEYINPUT43), .B(new_n584_), .C1(new_n455_), .C2(new_n459_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n644_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT44), .B(new_n644_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n435_), .A2(G29gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n643_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  NAND3_X1  g454(.A1(new_n651_), .A2(new_n456_), .A3(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G36gat), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n641_), .A2(G36gat), .A3(new_n452_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT45), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n657_), .A2(new_n660_), .A3(KEYINPUT46), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1329gat));
  NAND4_X1  g464(.A1(new_n651_), .A2(G43gat), .A3(new_n630_), .A4(new_n652_), .ZN(new_n666_));
  INV_X1    g465(.A(G43gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(new_n641_), .B2(new_n320_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g469(.A1(new_n651_), .A2(G50gat), .A3(new_n356_), .A4(new_n652_), .ZN(new_n671_));
  INV_X1    g470(.A(G50gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n672_), .B1(new_n641_), .B2(new_n633_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT112), .ZN(G1331gat));
  NOR2_X1   g474(.A1(new_n544_), .A2(new_n241_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n646_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(new_n606_), .ZN(new_n678_));
  INV_X1    g477(.A(G57gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n435_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n544_), .A2(new_n605_), .A3(new_n241_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n613_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G57gat), .B1(new_n683_), .B2(new_n453_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n680_), .A2(new_n684_), .ZN(G1332gat));
  NOR2_X1   g484(.A1(new_n452_), .A2(G64gat), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT113), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n678_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G64gat), .B1(new_n683_), .B2(new_n452_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(KEYINPUT48), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(KEYINPUT48), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(G1333gat));
  INV_X1    g491(.A(G71gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n682_), .B2(new_n630_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n678_), .A2(new_n693_), .A3(new_n630_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1334gat));
  INV_X1    g497(.A(G78gat), .ZN(new_n699_));
  INV_X1    g498(.A(new_n633_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n682_), .B2(new_n700_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT50), .Z(new_n702_));
  NAND3_X1  g501(.A1(new_n678_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1335gat));
  OR2_X1    g503(.A1(new_n647_), .A2(new_n648_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n676_), .A2(new_n605_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT115), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n708_), .A2(new_n453_), .A3(new_n480_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n677_), .A2(new_n605_), .A3(new_n612_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n435_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1336gat));
  OAI21_X1  g511(.A(G92gat), .B1(new_n708_), .B2(new_n452_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(new_n481_), .A3(new_n456_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT116), .ZN(G1337gat));
  OAI21_X1  g515(.A(G99gat), .B1(new_n708_), .B2(new_n320_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n710_), .A2(new_n630_), .A3(new_n476_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(G1338gat));
  NAND3_X1  g520(.A1(new_n710_), .A2(new_n477_), .A3(new_n356_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n356_), .B(new_n707_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G106gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G106gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g527(.A(new_n474_), .B1(new_n559_), .B2(new_n489_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n529_), .B(new_n514_), .C1(new_n729_), .C2(new_n525_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n462_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT120), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n530_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n515_), .B1(new_n519_), .B2(new_n526_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n736_), .A2(KEYINPUT55), .A3(new_n462_), .A4(new_n529_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT120), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n730_), .A2(new_n738_), .A3(new_n731_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n733_), .A2(new_n735_), .A3(new_n737_), .A4(new_n739_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n740_), .A2(KEYINPUT56), .A3(new_n535_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT56), .B1(new_n740_), .B2(new_n535_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(KEYINPUT121), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n535_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT56), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(KEYINPUT121), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n221_), .A2(new_n230_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n238_), .B1(new_n747_), .B2(new_n228_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n221_), .A2(new_n227_), .A3(G229gat), .A4(G233gat), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n232_), .A2(new_n238_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n542_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n746_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT122), .B1(new_n743_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT58), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT122), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n744_), .A2(new_n745_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT121), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n740_), .A2(KEYINPUT56), .A3(new_n535_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n751_), .B1(new_n742_), .B2(KEYINPUT121), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n756_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT58), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n755_), .A2(new_n585_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n241_), .A2(new_n542_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n541_), .A2(new_n542_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n750_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT57), .B1(new_n771_), .B2(new_n582_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT57), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n773_), .B(new_n612_), .C1(new_n768_), .C2(new_n770_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n604_), .B1(new_n765_), .B2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n584_), .A2(new_n544_), .A3(new_n242_), .A4(new_n604_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(KEYINPUT118), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(KEYINPUT118), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT119), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n779_), .A2(new_n783_), .A3(new_n780_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n778_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n786_));
  AOI211_X1 g585(.A(KEYINPUT119), .B(KEYINPUT54), .C1(new_n777_), .C2(KEYINPUT118), .ZN(new_n787_));
  INV_X1    g586(.A(new_n778_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n776_), .A2(new_n785_), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n457_), .A2(new_n630_), .A3(new_n435_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(G113gat), .B1(new_n792_), .B2(new_n241_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT123), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT59), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n766_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n770_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n582_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n773_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n771_), .A2(KEYINPUT57), .A3(new_n582_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n585_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n756_), .B(KEYINPUT58), .C1(new_n760_), .C2(new_n761_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n799_), .B(new_n800_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n786_), .A2(new_n787_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n803_), .A2(new_n605_), .B1(new_n804_), .B2(new_n778_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n788_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n795_), .B(new_n791_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n801_), .A2(new_n802_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n799_), .A2(new_n800_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n605_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n804_), .A2(new_n778_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n806_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n791_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT59), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n794_), .B1(new_n807_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n795_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(KEYINPUT59), .A3(new_n813_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(KEYINPUT123), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n241_), .A2(G113gat), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT124), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n793_), .B1(new_n819_), .B2(new_n821_), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n544_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n792_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n544_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n823_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n792_), .B2(new_n604_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n605_), .A2(new_n297_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n819_), .B2(new_n829_), .ZN(G1342gat));
  AOI21_X1  g629(.A(G134gat), .B1(new_n792_), .B2(new_n612_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n584_), .A2(new_n295_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n819_), .B2(new_n832_), .ZN(G1343gat));
  INV_X1    g632(.A(new_n356_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n630_), .A2(new_n453_), .A3(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n812_), .A2(new_n452_), .A3(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n242_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(new_n321_), .ZN(G1344gat));
  NOR2_X1   g637(.A1(new_n836_), .A2(new_n544_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(new_n322_), .ZN(G1345gat));
  NOR2_X1   g639(.A1(new_n836_), .A2(new_n605_), .ZN(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT61), .B(G155gat), .Z(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1346gat));
  INV_X1    g642(.A(G162gat), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n836_), .A2(new_n844_), .A3(new_n584_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n836_), .B2(new_n582_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT125), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT125), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n848_), .B(new_n844_), .C1(new_n836_), .C2(new_n582_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n845_), .B1(new_n847_), .B2(new_n849_), .ZN(G1347gat));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n456_), .A2(new_n458_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n700_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n241_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n790_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G169gat), .B1(new_n855_), .B2(KEYINPUT126), .ZN(new_n856_));
  INV_X1    g655(.A(new_n854_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n812_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n851_), .B1(new_n856_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n855_), .A2(new_n246_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n244_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n863_), .B(KEYINPUT62), .C1(new_n859_), .C2(new_n858_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n862_), .A3(new_n864_), .ZN(G1348gat));
  AND2_X1   g664(.A1(new_n812_), .A2(new_n853_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G176gat), .B1(new_n866_), .B2(new_n614_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n790_), .A2(new_n356_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n852_), .A2(new_n243_), .A3(new_n544_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(G1349gat));
  NAND4_X1  g669(.A1(new_n868_), .A2(new_n456_), .A3(new_n458_), .A4(new_n604_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n605_), .B1(new_n278_), .B2(new_n276_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n871_), .A2(new_n254_), .B1(new_n866_), .B2(new_n872_), .ZN(G1350gat));
  NAND4_X1  g672(.A1(new_n866_), .A2(new_n283_), .A3(new_n274_), .A4(new_n612_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n866_), .A2(new_n585_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n255_), .ZN(G1351gat));
  NAND4_X1  g675(.A1(new_n456_), .A2(new_n320_), .A3(new_n453_), .A4(new_n356_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n790_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n241_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n614_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g681(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT127), .ZN(new_n884_));
  NAND2_X1  g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n878_), .A2(new_n604_), .A3(new_n884_), .A4(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n883_), .A2(KEYINPUT127), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1354gat));
  INV_X1    g687(.A(G218gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n878_), .A2(new_n889_), .A3(new_n612_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n790_), .A2(new_n584_), .A3(new_n877_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1355gat));
endmodule


