//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_, new_n973_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G43gat), .B(G50gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(G29gat), .B(G36gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT8), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(KEYINPUT67), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT7), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT6), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n213_), .B1(new_n218_), .B2(new_n224_), .ZN(new_n225_));
  AOI211_X1 g024(.A(new_n223_), .B(new_n212_), .C1(new_n215_), .C2(new_n217_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228_));
  OR2_X1    g027(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n228_), .B1(new_n231_), .B2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(G106gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n229_), .A2(KEYINPUT64), .A3(new_n233_), .A4(new_n230_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n234_), .A3(new_n217_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n222_), .A2(KEYINPUT65), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n237_), .A2(KEYINPUT9), .B1(new_n219_), .B2(new_n220_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT9), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n222_), .A2(KEYINPUT65), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n236_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n235_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n210_), .B1(new_n227_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n214_), .B(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT6), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n216_), .B(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n224_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n212_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n218_), .A2(new_n224_), .A3(new_n213_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n217_), .A2(new_n234_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n238_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n232_), .B(new_n254_), .C1(new_n255_), .C2(new_n241_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n208_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G232gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT35), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n245_), .A2(KEYINPUT75), .A3(new_n258_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT73), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n245_), .A2(new_n266_), .A3(new_n258_), .A4(new_n263_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n261_), .A2(new_n262_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n245_), .A2(new_n258_), .A3(new_n263_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT75), .ZN(new_n271_));
  OAI221_X1 g070(.A(KEYINPUT73), .B1(new_n262_), .B2(new_n261_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G190gat), .B(G218gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(G134gat), .B(G162gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT36), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n269_), .A2(new_n272_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n276_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n278_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n281_), .ZN(new_n283_));
  AOI211_X1 g082(.A(new_n279_), .B(new_n283_), .C1(new_n269_), .C2(new_n272_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT37), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n269_), .A2(new_n272_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT74), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n283_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT37), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n280_), .A2(new_n281_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .A4(new_n278_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n285_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  INV_X1    g092(.A(G1gat), .ZN(new_n294_));
  INV_X1    g093(.A(G8gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT14), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT76), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G231gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G57gat), .B(G64gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G71gat), .B(G78gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(KEYINPUT11), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(KEYINPUT11), .ZN(new_n308_));
  INV_X1    g107(.A(new_n306_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n305_), .A2(KEYINPUT11), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n304_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n302_), .A2(new_n303_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n307_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n302_), .A2(new_n303_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G127gat), .B(G155gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G183gat), .B(G211gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT17), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n313_), .A2(new_n317_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n322_), .A2(KEYINPUT17), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n313_), .A2(new_n317_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n313_), .A2(KEYINPUT68), .A3(new_n317_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT78), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n332_), .A2(new_n336_), .A3(new_n333_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n326_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n292_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT79), .ZN(new_n340_));
  OR2_X1    g139(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n341_));
  NAND2_X1  g140(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n315_), .B(new_n331_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n253_), .A2(new_n256_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT12), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n343_), .A2(new_n344_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G230gat), .A2(G233gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n312_), .A2(KEYINPUT12), .A3(new_n307_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT69), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n352_), .A2(new_n344_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n352_), .B2(new_n344_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n349_), .A2(new_n350_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n348_), .A2(new_n345_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n350_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G120gat), .B(G148gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(G176gat), .B(G204gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n357_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n341_), .B(new_n342_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n369_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n371_), .A2(KEYINPUT71), .A3(KEYINPUT13), .A4(new_n367_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n210_), .A2(new_n301_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n257_), .A2(new_n300_), .A3(new_n299_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G229gat), .A2(G233gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT80), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n381_), .A3(new_n378_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n301_), .A2(new_n208_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n376_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(G229gat), .A3(G233gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G113gat), .B(G141gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT81), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G169gat), .B(G197gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n380_), .A2(new_n382_), .A3(new_n385_), .A4(new_n390_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n374_), .A2(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(G1gat), .B(G29gat), .Z(new_n396_));
  XNOR2_X1  g195(.A(G57gat), .B(G85gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(G141gat), .B(G148gat), .Z(new_n403_));
  NAND2_X1  g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT1), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT89), .ZN(new_n406_));
  INV_X1    g205(.A(G155gat), .ZN(new_n407_));
  INV_X1    g206(.A(G162gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT89), .B1(G155gat), .B2(G162gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n403_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n409_), .A2(new_n404_), .A3(new_n410_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n415_));
  INV_X1    g214(.A(G141gat), .ZN(new_n416_));
  INV_X1    g215(.A(G148gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G141gat), .A2(G148gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT2), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n418_), .A2(new_n421_), .A3(new_n422_), .A4(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n413_), .A2(new_n414_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n414_), .B1(new_n413_), .B2(new_n424_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n412_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT96), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G127gat), .B(G134gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G113gat), .B(G120gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT87), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n429_), .A2(new_n430_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n429_), .A2(new_n430_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n432_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n427_), .A2(new_n428_), .A3(new_n437_), .ZN(new_n438_));
  AND4_X1   g237(.A1(new_n421_), .A2(new_n418_), .A3(new_n422_), .A4(new_n423_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n409_), .A2(new_n404_), .A3(new_n410_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT90), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n413_), .A2(new_n414_), .A3(new_n424_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n405_), .A2(new_n411_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n441_), .A2(new_n442_), .B1(new_n443_), .B2(new_n403_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n433_), .A2(new_n431_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n438_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n428_), .B1(new_n427_), .B2(new_n437_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT4), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT4), .B1(new_n427_), .B2(new_n437_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n402_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT96), .B1(new_n444_), .B2(new_n436_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n438_), .A3(new_n446_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n402_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n401_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n454_), .A2(new_n455_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n450_), .B1(new_n454_), .B2(KEYINPUT4), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n458_), .B(new_n400_), .C1(new_n459_), .C2(new_n402_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G218gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G211gat), .ZN(new_n463_));
  INV_X1    g262(.A(G211gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(G218gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT21), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G197gat), .B(G204gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n463_), .A2(new_n465_), .A3(KEYINPUT21), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n469_), .A2(KEYINPUT21), .A3(new_n463_), .A4(new_n465_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G183gat), .A2(G190gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(KEYINPUT84), .A2(G183gat), .A3(G190gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT23), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT23), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(G183gat), .A3(G190gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G183gat), .ZN(new_n483_));
  INV_X1    g282(.A(G190gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n487_));
  INV_X1    g286(.A(G176gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n488_), .B1(new_n489_), .B2(G169gat), .ZN(new_n490_));
  INV_X1    g289(.A(G169gat), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(KEYINPUT85), .B2(KEYINPUT22), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n487_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(G169gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(KEYINPUT85), .A3(KEYINPUT22), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT86), .A4(new_n488_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G169gat), .A2(G176gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n486_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n500_));
  AND2_X1   g299(.A1(G169gat), .A2(G176gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT83), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n491_), .A2(new_n488_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n503_), .A2(new_n504_), .A3(KEYINPUT24), .A4(new_n498_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n475_), .A2(new_n480_), .ZN(new_n507_));
  AND3_X1   g306(.A1(KEYINPUT84), .A2(G183gat), .A3(G190gat), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT84), .B1(G183gat), .B2(G190gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n507_), .B1(new_n510_), .B2(new_n480_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n503_), .A2(KEYINPUT24), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n483_), .A2(KEYINPUT25), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT82), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT26), .B(G190gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT25), .B(G183gat), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n516_), .B(new_n517_), .C1(new_n518_), .C2(new_n515_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n506_), .A2(new_n511_), .A3(new_n513_), .A4(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n474_), .A2(new_n499_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n491_), .A2(KEYINPUT22), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT22), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(G169gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n524_), .A3(new_n488_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n498_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(new_n511_), .B2(new_n485_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT25), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(G183gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n484_), .A2(KEYINPUT26), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT26), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(G190gat), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n514_), .A2(new_n529_), .A3(new_n530_), .A4(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n503_), .A2(KEYINPUT24), .A3(new_n498_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT93), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(KEYINPUT93), .A3(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n512_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n527_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(KEYINPUT20), .B(new_n521_), .C1(new_n541_), .C2(new_n474_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G226gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n542_), .A2(KEYINPUT94), .A3(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n499_), .A2(new_n520_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n474_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n538_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT93), .B1(new_n533_), .B2(new_n534_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n540_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n527_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n474_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n545_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n559_), .A2(KEYINPUT20), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n548_), .A2(new_n549_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G8gat), .B(G36gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G64gat), .B(G92gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT32), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n552_), .A2(new_n557_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n545_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n555_), .A2(new_n556_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n551_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n572_), .A2(KEYINPUT20), .A3(new_n559_), .A4(new_n521_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n567_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n561_), .A2(new_n567_), .B1(new_n576_), .B2(KEYINPUT99), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n576_), .A2(KEYINPUT99), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n461_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n460_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AOI211_X1 g381(.A(new_n455_), .B(new_n450_), .C1(new_n454_), .C2(KEYINPUT4), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n454_), .A2(new_n455_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT33), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n401_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n580_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n558_), .A2(new_n560_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n542_), .A2(KEYINPUT94), .A3(new_n545_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT94), .B1(new_n542_), .B2(new_n545_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n566_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n588_), .B(new_n566_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n586_), .A2(new_n587_), .A3(new_n593_), .A4(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n579_), .B1(new_n582_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n436_), .B(KEYINPUT88), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G71gat), .B(G99gat), .ZN(new_n598_));
  INV_X1    g397(.A(G43gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G227gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(G15gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n600_), .B(new_n602_), .Z(new_n603_));
  NAND3_X1  g402(.A1(new_n499_), .A2(new_n520_), .A3(KEYINPUT30), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT30), .B1(new_n499_), .B2(new_n520_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n603_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n600_), .B(new_n602_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n604_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT31), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n607_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n607_), .B2(new_n610_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n597_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n605_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n609_), .B1(new_n608_), .B2(new_n604_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT31), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n607_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n597_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G228gat), .A2(G233gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT29), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n444_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n474_), .B1(new_n427_), .B2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n626_), .B1(new_n629_), .B2(new_n622_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G78gat), .B(G106gat), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n631_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n626_), .B(new_n633_), .C1(new_n629_), .C2(new_n622_), .ZN(new_n634_));
  XOR2_X1   g433(.A(G22gat), .B(G50gat), .Z(new_n635_));
  AND3_X1   g434(.A1(new_n632_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n444_), .A2(new_n625_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT28), .Z(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n636_), .A2(new_n637_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n635_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n551_), .B1(new_n444_), .B2(new_n627_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n623_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n633_), .B1(new_n644_), .B2(new_n626_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n634_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n632_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n639_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n621_), .B1(new_n641_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n612_), .A2(new_n613_), .A3(new_n597_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n619_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n654_), .B1(new_n641_), .B2(new_n649_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n640_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n647_), .A2(new_n639_), .A3(new_n648_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n621_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT27), .B1(new_n593_), .B2(new_n594_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT27), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n574_), .B2(new_n592_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(new_n594_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n660_), .A2(new_n461_), .A3(new_n663_), .ZN(new_n664_));
  AOI22_X1  g463(.A1(new_n596_), .A2(new_n651_), .B1(new_n659_), .B2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n395_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n340_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT100), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n340_), .A2(new_n669_), .A3(new_n666_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n294_), .A3(new_n461_), .ZN(new_n672_));
  XOR2_X1   g471(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n282_), .A2(new_n284_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n665_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n677_), .A2(new_n394_), .A3(new_n374_), .A4(new_n338_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT103), .Z(new_n679_));
  AND2_X1   g478(.A1(new_n457_), .A2(new_n460_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G1gat), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n673_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n671_), .A2(new_n294_), .A3(new_n461_), .A4(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT102), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(KEYINPUT102), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n674_), .B(new_n681_), .C1(new_n684_), .C2(new_n685_), .ZN(G1324gat));
  NOR2_X1   g485(.A1(new_n660_), .A2(new_n663_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G8gat), .B1(new_n678_), .B2(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT39), .Z(new_n689_));
  NOR2_X1   g488(.A1(new_n687_), .A2(G8gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n668_), .A2(new_n670_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT104), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n668_), .A2(new_n693_), .A3(new_n670_), .A4(new_n690_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n689_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(G1325gat));
  OAI21_X1  g496(.A(G15gat), .B1(new_n679_), .B2(new_n621_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n699_), .ZN(new_n701_));
  OAI211_X1 g500(.A(G15gat), .B(new_n701_), .C1(new_n679_), .C2(new_n621_), .ZN(new_n702_));
  OR3_X1    g501(.A1(new_n667_), .A2(G15gat), .A3(new_n621_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n700_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT107), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n700_), .A2(new_n706_), .A3(new_n702_), .A4(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1326gat));
  NOR2_X1   g507(.A1(new_n641_), .A2(new_n649_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G22gat), .B1(new_n679_), .B2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n712_));
  OR2_X1    g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n712_), .ZN(new_n714_));
  OR3_X1    g513(.A1(new_n667_), .A2(G22gat), .A3(new_n710_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(new_n714_), .A3(new_n715_), .ZN(G1327gat));
  NOR2_X1   g515(.A1(new_n338_), .A2(new_n675_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n666_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G29gat), .B1(new_n718_), .B2(new_n461_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n665_), .B2(new_n292_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n285_), .A2(new_n291_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n659_), .A2(new_n664_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n548_), .A2(new_n549_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n566_), .B1(new_n724_), .B2(new_n588_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n594_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n727_), .A2(new_n581_), .A3(new_n586_), .A4(new_n587_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n650_), .B1(new_n728_), .B2(new_n579_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n721_), .B(new_n722_), .C1(new_n723_), .C2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n720_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n395_), .A2(new_n338_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(G29gat), .A3(new_n461_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n733_), .A2(new_n734_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n733_), .A2(KEYINPUT109), .A3(new_n734_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n719_), .B1(new_n737_), .B2(new_n742_), .ZN(G1328gat));
  NAND2_X1  g542(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(G36gat), .ZN(new_n748_));
  INV_X1    g547(.A(new_n687_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n718_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT45), .Z(new_n751_));
  NOR2_X1   g550(.A1(new_n735_), .A2(new_n687_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n748_), .B1(new_n742_), .B2(new_n752_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n744_), .B(new_n747_), .C1(new_n751_), .C2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n742_), .A2(new_n752_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(G36gat), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n750_), .B(KEYINPUT45), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n756_), .A2(new_n745_), .A3(new_n746_), .A4(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n754_), .A2(new_n758_), .ZN(G1329gat));
  NOR2_X1   g558(.A1(new_n621_), .A2(new_n599_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n742_), .A2(new_n736_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n718_), .A2(new_n654_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n599_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OR3_X1    g563(.A1(new_n761_), .A2(KEYINPUT47), .A3(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT47), .B1(new_n761_), .B2(new_n764_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1330gat));
  INV_X1    g566(.A(G50gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n709_), .A2(new_n768_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT111), .Z(new_n770_));
  NAND2_X1  g569(.A1(new_n718_), .A2(new_n770_), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n710_), .B(new_n735_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n768_), .ZN(G1331gat));
  INV_X1    g572(.A(new_n394_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n373_), .A2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(new_n665_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n340_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(G57gat), .B1(new_n778_), .B2(new_n461_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n337_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n336_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n325_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n775_), .A2(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n783_), .A2(new_n677_), .A3(G57gat), .A4(new_n461_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT112), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n784_), .A2(KEYINPUT112), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n779_), .B1(new_n785_), .B2(new_n786_), .ZN(G1332gat));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n677_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G64gat), .B1(new_n788_), .B2(new_n687_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT48), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n687_), .A2(G64gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n777_), .B2(new_n791_), .ZN(G1333gat));
  OAI21_X1  g591(.A(G71gat), .B1(new_n788_), .B2(new_n621_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT49), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n621_), .A2(G71gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n777_), .B2(new_n795_), .ZN(G1334gat));
  OAI21_X1  g595(.A(G78gat), .B1(new_n788_), .B2(new_n710_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT50), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n710_), .A2(G78gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n777_), .B2(new_n799_), .ZN(G1335gat));
  NAND3_X1  g599(.A1(new_n782_), .A2(new_n373_), .A3(new_n774_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT113), .B1(new_n731_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n804_), .B(new_n801_), .C1(new_n720_), .C2(new_n730_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(G85gat), .B1(new_n806_), .B2(new_n680_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n776_), .A2(new_n717_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(new_n219_), .A3(new_n461_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(G1336gat));
  OAI21_X1  g610(.A(G92gat), .B1(new_n806_), .B2(new_n687_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n220_), .A3(new_n749_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1337gat));
  OR3_X1    g613(.A1(new_n808_), .A2(new_n231_), .A3(new_n621_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n654_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(G99gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n816_), .B2(G99gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n815_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OR2_X1    g619(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n821_));
  NAND2_X1  g620(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n816_), .A2(G99gat), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT114), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n816_), .A2(new_n817_), .A3(G99gat), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n827_), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n815_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n823_), .A2(new_n828_), .ZN(G1338gat));
  NAND3_X1  g628(.A1(new_n731_), .A2(new_n709_), .A3(new_n802_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G106gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT52), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n809_), .A2(new_n233_), .A3(new_n709_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(G1339gat));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n347_), .B(new_n348_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n359_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n349_), .A2(new_n356_), .A3(KEYINPUT55), .A4(new_n350_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n359_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n365_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n842_), .A2(KEYINPUT56), .A3(new_n365_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n390_), .B1(new_n384_), .B2(new_n378_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n377_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n378_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n393_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n368_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT118), .B1(new_n847_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n292_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n842_), .A2(KEYINPUT56), .A3(new_n365_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT56), .B1(new_n842_), .B2(new_n365_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n852_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT58), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n394_), .A2(new_n367_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n851_), .B1(new_n371_), .B2(new_n367_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n676_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n855_), .A2(new_n861_), .B1(KEYINPUT57), .B2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT117), .B1(new_n866_), .B2(KEYINPUT57), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n394_), .A2(new_n367_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n675_), .B1(new_n870_), .B2(new_n864_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n868_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n338_), .B1(new_n867_), .B2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n374_), .A2(new_n292_), .A3(new_n774_), .A4(new_n338_), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT54), .Z(new_n878_));
  OR2_X1    g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n687_), .A2(new_n461_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n655_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(G113gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n884_), .A3(new_n394_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n853_), .A2(new_n854_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n858_), .A2(new_n859_), .A3(new_n854_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n722_), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n886_), .A2(new_n888_), .B1(new_n873_), .B2(new_n871_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n866_), .A2(KEYINPUT57), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n782_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n877_), .B(KEYINPUT54), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n881_), .B(KEYINPUT119), .Z(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(KEYINPUT59), .ZN(new_n895_));
  AOI221_X4 g694(.A(new_n774_), .B1(new_n893_), .B2(new_n895_), .C1(new_n882_), .C2(KEYINPUT59), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n885_), .B1(new_n896_), .B2(new_n884_), .ZN(G1340gat));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n898_));
  INV_X1    g697(.A(G120gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n373_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n883_), .A2(new_n901_), .ZN(new_n902_));
  AOI221_X4 g701(.A(new_n374_), .B1(new_n893_), .B2(new_n895_), .C1(new_n882_), .C2(KEYINPUT59), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n899_), .ZN(G1341gat));
  INV_X1    g703(.A(G127gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n883_), .A2(new_n905_), .A3(new_n338_), .ZN(new_n906_));
  AOI221_X4 g705(.A(new_n782_), .B1(new_n893_), .B2(new_n895_), .C1(new_n882_), .C2(KEYINPUT59), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n905_), .ZN(G1342gat));
  INV_X1    g707(.A(G134gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n883_), .A2(new_n909_), .A3(new_n676_), .ZN(new_n910_));
  AOI221_X4 g709(.A(new_n292_), .B1(new_n893_), .B2(new_n895_), .C1(new_n882_), .C2(KEYINPUT59), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n909_), .ZN(G1343gat));
  INV_X1    g711(.A(new_n658_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n880_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n879_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n774_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n416_), .ZN(G1344gat));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n374_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT120), .B(G148gat), .Z(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n918_), .B(new_n920_), .ZN(G1345gat));
  NOR2_X1   g720(.A1(new_n915_), .A2(new_n782_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT61), .B(G155gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n922_), .B(new_n924_), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n915_), .B2(new_n292_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n676_), .A2(new_n408_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n915_), .B2(new_n927_), .ZN(G1347gat));
  NOR3_X1   g727(.A1(new_n687_), .A2(new_n655_), .A3(new_n461_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n893_), .A2(new_n394_), .A3(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n930_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n522_), .A2(new_n524_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n933_), .B2(new_n930_), .ZN(new_n934_));
  AOI21_X1  g733(.A(KEYINPUT62), .B1(new_n930_), .B2(G169gat), .ZN(new_n935_));
  OR2_X1    g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1348gat));
  NAND2_X1  g735(.A1(new_n893_), .A2(new_n929_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n488_), .B1(new_n937_), .B2(new_n374_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n374_), .A2(new_n488_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n929_), .B(new_n939_), .C1(new_n876_), .C2(new_n878_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n940_), .A2(KEYINPUT121), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(KEYINPUT121), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n938_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  OAI211_X1 g744(.A(KEYINPUT122), .B(new_n938_), .C1(new_n941_), .C2(new_n942_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1349gat));
  NOR3_X1   g746(.A1(new_n937_), .A2(new_n518_), .A3(new_n782_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n879_), .A2(new_n338_), .A3(new_n929_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(new_n483_), .ZN(G1350gat));
  OAI21_X1  g749(.A(G190gat), .B1(new_n937_), .B2(new_n292_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n676_), .A2(new_n517_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n937_), .B2(new_n952_), .ZN(G1351gat));
  NOR2_X1   g752(.A1(new_n687_), .A2(new_n461_), .ZN(new_n954_));
  OAI211_X1 g753(.A(new_n913_), .B(new_n954_), .C1(new_n876_), .C2(new_n878_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n955_), .A2(new_n774_), .ZN(new_n956_));
  AND3_X1   g755(.A1(new_n956_), .A2(KEYINPUT123), .A3(G197gat), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(G197gat), .ZN(new_n958_));
  OAI21_X1  g757(.A(KEYINPUT123), .B1(new_n956_), .B2(G197gat), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n957_), .B1(new_n958_), .B2(new_n959_), .ZN(G1352gat));
  NOR2_X1   g759(.A1(new_n955_), .A2(new_n374_), .ZN(new_n961_));
  XOR2_X1   g760(.A(KEYINPUT124), .B(G204gat), .Z(new_n962_));
  XNOR2_X1  g761(.A(new_n961_), .B(new_n962_), .ZN(G1353gat));
  INV_X1    g762(.A(new_n955_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n782_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(KEYINPUT125), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(KEYINPUT126), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n966_), .B(new_n969_), .ZN(G1354gat));
  AOI21_X1  g769(.A(G218gat), .B1(new_n964_), .B2(new_n676_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n722_), .A2(G218gat), .ZN(new_n972_));
  XOR2_X1   g771(.A(new_n972_), .B(KEYINPUT127), .Z(new_n973_));
  AOI21_X1  g772(.A(new_n971_), .B1(new_n964_), .B2(new_n973_), .ZN(G1355gat));
endmodule


