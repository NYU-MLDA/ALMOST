//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n204_), .B2(KEYINPUT21), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT90), .A2(KEYINPUT21), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n205_), .B(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G183gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT25), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G183gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n212_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT23), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G183gat), .A3(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT82), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n209_), .A2(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n226_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT92), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT92), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n226_), .A2(new_n232_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n220_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G169gat), .ZN(new_n235_));
  INV_X1    g034(.A(G176gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n211_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n222_), .A2(new_n224_), .ZN(new_n239_));
  OR2_X1    g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n208_), .B1(new_n234_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT20), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT83), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n212_), .A2(new_n228_), .A3(new_n239_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n217_), .A2(KEYINPUT79), .A3(KEYINPUT80), .A4(G183gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n219_), .A2(KEYINPUT79), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT79), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT80), .B1(new_n216_), .B2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n249_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n247_), .B1(new_n253_), .B2(new_n214_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT81), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n237_), .A2(new_n255_), .B1(G169gat), .B2(G176gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n226_), .A2(new_n229_), .A3(new_n240_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n235_), .A2(KEYINPUT81), .A3(new_n236_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n245_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n254_), .A2(new_n259_), .A3(new_n245_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n208_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n244_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G8gat), .B(G36gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT18), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G64gat), .ZN(new_n271_));
  INV_X1    g070(.A(G92gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n208_), .A2(new_n234_), .A3(new_n241_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT20), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n262_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n208_), .B1(new_n277_), .B2(new_n260_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n267_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n276_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n268_), .A2(new_n273_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT27), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT97), .B1(new_n274_), .B2(new_n275_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT97), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n234_), .A2(new_n241_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n284_), .B(KEYINPUT20), .C1(new_n285_), .C2(new_n208_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n286_), .A3(new_n278_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n267_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT98), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(KEYINPUT98), .A3(new_n267_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n265_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n279_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n273_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n282_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n280_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n279_), .B1(new_n244_), .B2(new_n264_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n295_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT27), .B1(new_n299_), .B2(new_n281_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT99), .B1(new_n296_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n300_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT99), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n288_), .A2(new_n289_), .B1(new_n292_), .B2(new_n279_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n273_), .B1(new_n304_), .B2(new_n291_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n302_), .B(new_n303_), .C1(new_n305_), .C2(new_n282_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT87), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT86), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n310_), .A2(new_n312_), .B1(new_n313_), .B2(KEYINPUT85), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT86), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT87), .B1(new_n315_), .B2(KEYINPUT2), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n311_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n318_), .A2(new_n319_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n313_), .A2(KEYINPUT85), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n314_), .A2(new_n317_), .A3(new_n320_), .A4(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G155gat), .B(G162gat), .Z(new_n323_));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n318_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n326_), .A2(new_n311_), .A3(new_n327_), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n322_), .A2(new_n323_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT89), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n331_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n263_), .B1(G228gat), .B2(G233gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n330_), .B2(new_n329_), .ZN(new_n337_));
  XOR2_X1   g136(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n338_));
  OAI21_X1  g137(.A(new_n208_), .B1(new_n329_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G228gat), .A3(G233gat), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n335_), .A2(new_n337_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n335_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G78gat), .B(G106gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G22gat), .B(G50gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  OR3_X1    g145(.A1(new_n341_), .A2(new_n342_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G127gat), .B(G134gat), .Z(new_n351_));
  XOR2_X1   g150(.A(G113gat), .B(G120gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n329_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n322_), .A2(new_n323_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n325_), .A2(new_n328_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n354_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT94), .B1(new_n363_), .B2(KEYINPUT4), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n329_), .A2(new_n353_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT94), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n329_), .A2(new_n353_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT93), .B1(new_n371_), .B2(new_n367_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT93), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n363_), .A2(new_n373_), .A3(KEYINPUT4), .A4(new_n370_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n369_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n359_), .B1(new_n375_), .B2(new_n356_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT0), .ZN(new_n378_));
  INV_X1    g177(.A(G57gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(G85gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n383_), .B(new_n359_), .C1(new_n375_), .C2(new_n356_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G15gat), .B(G43gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT31), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT30), .B1(new_n261_), .B2(new_n262_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT30), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n277_), .A2(new_n390_), .A3(new_n260_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G71gat), .B(G99gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n353_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n353_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n388_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n401_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(new_n387_), .A3(new_n399_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n385_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n307_), .A2(KEYINPUT100), .A3(new_n350_), .A4(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n301_), .A2(new_n405_), .A3(new_n306_), .A4(new_n350_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT100), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n296_), .A2(new_n300_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n385_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n349_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n372_), .A2(new_n374_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n364_), .A2(new_n368_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n356_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(KEYINPUT33), .B(new_n381_), .C1(new_n415_), .C2(new_n358_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT95), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n356_), .A3(new_n414_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n381_), .B1(new_n357_), .B2(new_n355_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n420_), .A2(new_n299_), .A3(new_n281_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT95), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n376_), .A2(new_n422_), .A3(KEYINPUT33), .A4(new_n381_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n417_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n382_), .A2(KEYINPUT96), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n376_), .A2(new_n426_), .A3(new_n381_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n294_), .A2(KEYINPUT32), .A3(new_n273_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n273_), .A2(KEYINPUT32), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n297_), .A2(new_n298_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n382_), .A2(new_n384_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n424_), .A2(new_n429_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n412_), .B1(new_n434_), .B2(new_n349_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n402_), .A2(new_n404_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n406_), .A2(new_n409_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n439_));
  OR2_X1    g238(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n440_));
  INV_X1    g239(.A(G106gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G99gat), .A2(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G85gat), .A2(G92gat), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n449_), .A2(KEYINPUT9), .ZN(new_n450_));
  INV_X1    g249(.A(G85gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n272_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(KEYINPUT9), .A3(new_n449_), .ZN(new_n453_));
  AND4_X1   g252(.A1(new_n443_), .A2(new_n448_), .A3(new_n450_), .A4(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT7), .ZN(new_n455_));
  INV_X1    g254(.A(G99gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n441_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n457_), .A2(new_n446_), .A3(new_n447_), .A4(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n452_), .A2(new_n449_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT8), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n463_), .A3(new_n460_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n454_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G29gat), .B(G36gat), .Z(new_n466_));
  XOR2_X1   g265(.A(G43gat), .B(G50gat), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G232gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT34), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT69), .B(KEYINPUT35), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n465_), .A2(new_n472_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT15), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n468_), .A2(KEYINPUT15), .A3(new_n471_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI221_X1 g280(.A(new_n477_), .B1(new_n475_), .B2(new_n476_), .C1(new_n465_), .C2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT70), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n483_), .B1(new_n465_), .B2(new_n481_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n462_), .A2(new_n464_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n454_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n468_), .A2(KEYINPUT15), .A3(new_n471_), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT15), .B1(new_n468_), .B2(new_n471_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n487_), .A2(KEYINPUT70), .A3(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n477_), .A2(new_n484_), .A3(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n475_), .A2(new_n476_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n492_), .A2(KEYINPUT71), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT71), .B1(new_n492_), .B2(new_n493_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n482_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G190gat), .B(G218gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G134gat), .B(G162gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT36), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(KEYINPUT73), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT74), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n482_), .B(new_n505_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n502_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT73), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n508_), .A2(KEYINPUT74), .ZN(new_n511_));
  INV_X1    g310(.A(new_n496_), .ZN(new_n512_));
  OAI221_X1 g311(.A(new_n506_), .B1(new_n510_), .B2(new_n511_), .C1(new_n512_), .C2(new_n500_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT66), .ZN(new_n516_));
  INV_X1    g315(.A(G78gat), .ZN(new_n517_));
  AND2_X1   g316(.A1(KEYINPUT64), .A2(G71gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(KEYINPUT64), .A2(G71gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT64), .ZN(new_n521_));
  INV_X1    g320(.A(G71gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(KEYINPUT64), .A2(G71gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(G78gat), .A3(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G57gat), .B(G64gat), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n520_), .B(new_n525_), .C1(KEYINPUT11), .C2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT65), .ZN(new_n528_));
  INV_X1    g327(.A(G64gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(G57gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n379_), .A2(G64gat), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT11), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT65), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n520_), .A4(new_n525_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n526_), .A2(KEYINPUT11), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n528_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n537_), .B1(new_n528_), .B2(new_n535_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n487_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n518_), .A2(new_n519_), .A3(new_n517_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(new_n532_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n534_), .B1(new_n542_), .B2(new_n520_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n527_), .A2(KEYINPUT65), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n536_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n528_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n465_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n540_), .A2(new_n547_), .A3(KEYINPUT12), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n546_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n487_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n516_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  AOI211_X1 g354(.A(KEYINPUT66), .B(new_n555_), .C1(new_n548_), .C2(new_n551_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n540_), .B2(new_n547_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G120gat), .B(G148gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(G204gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT5), .B(G176gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT67), .Z(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT68), .B1(new_n558_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n552_), .A2(new_n553_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT66), .ZN(new_n566_));
  INV_X1    g365(.A(new_n557_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n555_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n516_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT68), .ZN(new_n571_));
  INV_X1    g370(.A(new_n563_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n566_), .A2(new_n567_), .A3(new_n569_), .A4(new_n562_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n564_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT13), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n564_), .A2(KEYINPUT13), .A3(new_n573_), .A4(new_n574_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT78), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G15gat), .B(G22gat), .ZN(new_n583_));
  INV_X1    g382(.A(G1gat), .ZN(new_n584_));
  INV_X1    g383(.A(G8gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT14), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT75), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT75), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n583_), .A2(new_n589_), .A3(new_n586_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G1gat), .B(G8gat), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n588_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n472_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n472_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n582_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n594_), .A2(new_n595_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n490_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n596_), .A3(new_n581_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G169gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(G197gat), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n580_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n599_), .A2(new_n602_), .A3(KEYINPUT78), .A4(new_n606_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n603_), .A2(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT17), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT76), .ZN(new_n619_));
  INV_X1    g418(.A(G231gat), .ZN(new_n620_));
  INV_X1    g419(.A(G233gat), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n545_), .A2(new_n546_), .A3(new_n622_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n619_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n625_), .A3(new_n619_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n600_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n628_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n600_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n630_), .A2(new_n626_), .A3(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n618_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n631_), .B1(new_n630_), .B2(new_n626_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n627_), .A2(new_n600_), .A3(new_n628_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT17), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n617_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n579_), .A2(new_n612_), .A3(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n439_), .A2(new_n515_), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n584_), .A3(new_n385_), .ZN(new_n643_));
  XOR2_X1   g442(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT104), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n420_), .A2(new_n299_), .A3(new_n281_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(KEYINPUT95), .B2(new_n416_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n429_), .A2(new_n648_), .A3(new_n423_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n433_), .A2(new_n430_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n349_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n412_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n438_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n409_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n407_), .A2(new_n408_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n653_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n510_), .B1(new_n512_), .B2(new_n500_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT103), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n656_), .A2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n641_), .B(KEYINPUT102), .Z(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G1gat), .B1(new_n662_), .B2(new_n411_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n646_), .B(new_n663_), .C1(new_n644_), .C2(new_n643_), .ZN(G1324gat));
  INV_X1    g463(.A(new_n307_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n642_), .A2(new_n585_), .A3(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n660_), .A2(new_n661_), .A3(new_n665_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G8gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G8gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT105), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n673_), .B(new_n666_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n672_), .A2(KEYINPUT40), .A3(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  OAI21_X1  g478(.A(G15gat), .B1(new_n662_), .B2(new_n438_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT106), .Z(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT41), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT41), .ZN(new_n683_));
  INV_X1    g482(.A(G15gat), .ZN(new_n684_));
  INV_X1    g483(.A(new_n438_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n642_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n682_), .A2(new_n683_), .A3(new_n686_), .ZN(G1326gat));
  OAI21_X1  g486(.A(G22gat), .B1(new_n662_), .B2(new_n350_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT42), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n350_), .A2(G22gat), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT107), .Z(new_n691_));
  NAND2_X1  g490(.A1(new_n642_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(G1327gat));
  NAND3_X1  g492(.A1(new_n579_), .A2(new_n612_), .A3(new_n639_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n439_), .A2(new_n658_), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n385_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n694_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n439_), .A2(KEYINPUT43), .A3(new_n514_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n656_), .B2(new_n515_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(G29gat), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n411_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n701_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n439_), .B2(new_n514_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n656_), .A2(new_n699_), .A3(new_n515_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n694_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT108), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n707_), .A2(new_n711_), .A3(new_n702_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n696_), .B1(new_n705_), .B2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n717_));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n307_), .B1(new_n710_), .B2(KEYINPUT44), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n712_), .B2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n695_), .A2(new_n718_), .A3(new_n665_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT45), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n716_), .B(new_n717_), .C1(new_n720_), .C2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n701_), .A2(new_n706_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n702_), .B1(new_n710_), .B2(KEYINPUT108), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n719_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G36gat), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n728_), .A2(new_n714_), .A3(new_n722_), .A4(new_n715_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n724_), .A2(new_n729_), .ZN(G1329gat));
  AOI21_X1  g529(.A(G43gat), .B1(new_n695_), .B2(new_n685_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n436_), .A2(G43gat), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n703_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n733_), .B2(new_n712_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g534(.A(G50gat), .B1(new_n695_), .B2(new_n349_), .ZN(new_n736_));
  INV_X1    g535(.A(G50gat), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n703_), .A2(new_n737_), .A3(new_n350_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n738_), .B2(new_n712_), .ZN(G1331gat));
  INV_X1    g538(.A(new_n579_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n612_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n660_), .A2(new_n740_), .A3(new_n741_), .A4(new_n640_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n411_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n741_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n744_), .A2(new_n515_), .A3(new_n639_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n656_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n379_), .A3(new_n385_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n743_), .A2(new_n748_), .ZN(G1332gat));
  OAI21_X1  g548(.A(G64gat), .B1(new_n742_), .B2(new_n307_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT48), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n747_), .A2(new_n529_), .A3(new_n665_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1333gat));
  OAI21_X1  g552(.A(G71gat), .B1(new_n742_), .B2(new_n438_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT49), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n685_), .A2(new_n522_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT110), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n746_), .B2(new_n757_), .ZN(G1334gat));
  OAI21_X1  g557(.A(G78gat), .B1(new_n742_), .B2(new_n350_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT50), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n747_), .A2(new_n517_), .A3(new_n349_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1335gat));
  NAND3_X1  g561(.A1(new_n740_), .A2(new_n741_), .A3(new_n639_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n439_), .A2(new_n658_), .A3(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n451_), .A3(new_n385_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(new_n385_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n765_), .B1(new_n767_), .B2(new_n451_), .ZN(G1336gat));
  NAND3_X1  g567(.A1(new_n764_), .A2(new_n272_), .A3(new_n665_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n766_), .A2(new_n665_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n272_), .ZN(G1337gat));
  NAND4_X1  g570(.A1(new_n764_), .A2(new_n436_), .A3(new_n440_), .A4(new_n442_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(KEYINPUT111), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n456_), .B1(new_n766_), .B2(new_n685_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(KEYINPUT111), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n776_), .B(new_n777_), .Z(G1338gat));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n350_), .B(new_n763_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT52), .B1(new_n781_), .B2(new_n441_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n763_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n349_), .B(new_n783_), .C1(new_n698_), .C2(new_n700_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n782_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n764_), .A2(new_n441_), .A3(new_n349_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n780_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n788_), .ZN(new_n790_));
  AOI211_X1 g589(.A(KEYINPUT112), .B(new_n790_), .C1(new_n782_), .C2(new_n786_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n779_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n786_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n788_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT112), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n787_), .A2(new_n780_), .A3(new_n788_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(KEYINPUT53), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n792_), .A2(new_n798_), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n548_), .A2(new_n555_), .A3(new_n551_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n565_), .B2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n554_), .A2(new_n556_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n801_), .B1(new_n807_), .B2(new_n563_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n566_), .A2(new_n569_), .A3(new_n806_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n802_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(KEYINPUT55), .B2(new_n568_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n572_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n808_), .A2(new_n813_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n574_), .A2(KEYINPUT114), .A3(new_n612_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT114), .B1(new_n574_), .B2(new_n612_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n581_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n601_), .A2(new_n596_), .A3(new_n582_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n607_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n610_), .A2(new_n820_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n814_), .A2(new_n817_), .B1(new_n575_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n658_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n800_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n575_), .A2(new_n821_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n572_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n801_), .B(new_n563_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n816_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n574_), .A2(new_n612_), .A3(KEYINPUT114), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n825_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT57), .A3(new_n658_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n824_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n821_), .A2(new_n574_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n827_), .B2(KEYINPUT116), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n808_), .A2(new_n837_), .A3(new_n813_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n836_), .A2(new_n838_), .A3(KEYINPUT58), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n836_), .B2(new_n838_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n514_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n639_), .B1(new_n834_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n509_), .A2(new_n640_), .A3(new_n513_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n844_), .A2(new_n577_), .A3(new_n578_), .A4(new_n741_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n845_), .A2(KEYINPUT113), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(KEYINPUT113), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n843_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n845_), .A2(KEYINPUT113), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n845_), .A2(KEYINPUT113), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(KEYINPUT54), .A3(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n842_), .A2(new_n848_), .A3(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n307_), .A2(new_n350_), .A3(new_n385_), .A4(new_n436_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT117), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n612_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n852_), .A2(new_n859_), .A3(new_n854_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n855_), .A2(KEYINPUT59), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n852_), .A2(new_n859_), .A3(new_n854_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(KEYINPUT118), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT119), .B(G113gat), .Z(new_n867_));
  NAND2_X1  g666(.A1(new_n612_), .A2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT120), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n857_), .B1(new_n866_), .B2(new_n869_), .ZN(G1340gat));
  NOR2_X1   g669(.A1(new_n579_), .A2(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n856_), .B1(KEYINPUT60), .B2(new_n871_), .ZN(new_n872_));
  AND4_X1   g671(.A1(new_n740_), .A2(new_n872_), .A3(new_n863_), .A4(new_n864_), .ZN(new_n873_));
  INV_X1    g672(.A(G120gat), .ZN(new_n874_));
  OAI22_X1  g673(.A1(new_n873_), .A2(new_n874_), .B1(KEYINPUT60), .B2(new_n872_), .ZN(G1341gat));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876_));
  INV_X1    g675(.A(G127gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n866_), .B2(new_n640_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n855_), .A2(G127gat), .A3(new_n639_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n876_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n879_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n639_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT121), .B(new_n881_), .C1(new_n882_), .C2(new_n877_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(G1342gat));
  OR3_X1    g683(.A1(new_n855_), .A2(G134gat), .A3(new_n659_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n514_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n886_));
  INV_X1    g685(.A(G134gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1343gat));
  NOR3_X1   g687(.A1(new_n685_), .A2(new_n350_), .A3(new_n411_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n852_), .A2(new_n307_), .A3(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n741_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT122), .B(G141gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1344gat));
  NOR2_X1   g692(.A1(new_n890_), .A2(new_n579_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g694(.A1(new_n890_), .A2(new_n639_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT61), .B(G155gat), .Z(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n890_), .B2(new_n514_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n659_), .A2(G162gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n890_), .B2(new_n900_), .ZN(G1347gat));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n852_), .A2(new_n350_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n438_), .A2(new_n307_), .A3(new_n385_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n612_), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(KEYINPUT123), .Z(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n902_), .B1(new_n907_), .B2(G169gat), .ZN(new_n908_));
  INV_X1    g707(.A(G169gat), .ZN(new_n909_));
  AOI211_X1 g708(.A(KEYINPUT62), .B(new_n909_), .C1(new_n903_), .C2(new_n906_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n903_), .A2(new_n904_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n612_), .A2(new_n235_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT124), .ZN(new_n913_));
  OAI22_X1  g712(.A1(new_n908_), .A2(new_n910_), .B1(new_n911_), .B2(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT125), .ZN(G1348gat));
  NOR2_X1   g714(.A1(new_n911_), .A2(new_n579_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT126), .B(G176gat), .Z(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1349gat));
  NOR2_X1   g717(.A1(new_n911_), .A2(new_n639_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(G183gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n920_), .B1(new_n219_), .B2(new_n919_), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n911_), .B2(new_n514_), .ZN(new_n922_));
  OR2_X1    g721(.A1(new_n659_), .A2(new_n214_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n911_), .B2(new_n923_), .ZN(G1351gat));
  NOR4_X1   g723(.A1(new_n685_), .A2(new_n350_), .A3(new_n385_), .A4(new_n307_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n852_), .A2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n612_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n740_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g729(.A1(new_n926_), .A2(new_n640_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  AND2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n931_), .B2(new_n932_), .ZN(G1354gat));
  NAND2_X1  g734(.A1(new_n926_), .A2(new_n515_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(G218gat), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n659_), .A2(G218gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n926_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


