//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(KEYINPUT74), .B(G15gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G22gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G1gat), .B(G8gat), .Z(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G57gat), .B(G64gat), .Z(new_n210_));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(KEYINPUT66), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT11), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G71gat), .B(G78gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n210_), .A2(new_n211_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n213_), .A2(KEYINPUT66), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n215_), .A2(new_n217_), .A3(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(KEYINPUT11), .B(new_n216_), .C1(new_n212_), .C2(new_n214_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n209_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G231gat), .A2(G233gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT75), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G127gat), .B(G155gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT16), .ZN(new_n230_));
  XOR2_X1   g029(.A(G183gat), .B(G211gat), .Z(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n233_), .A2(KEYINPUT17), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n227_), .A2(new_n228_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n227_), .A2(KEYINPUT17), .A3(new_n233_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT15), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n246_));
  INV_X1    g045(.A(G85gat), .ZN(new_n247_));
  INV_X1    g046(.A(G92gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G85gat), .A2(G92gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n246_), .B1(new_n251_), .B2(KEYINPUT9), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT6), .ZN(new_n255_));
  INV_X1    g054(.A(G99gat), .ZN(new_n256_));
  INV_X1    g055(.A(G106gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT10), .B(G99gat), .Z(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(new_n257_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT9), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT64), .B1(new_n264_), .B2(new_n246_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n254_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n266_));
  OR3_X1    g065(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n267_), .A2(new_n258_), .A3(new_n259_), .A4(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n251_), .A2(KEYINPUT65), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(KEYINPUT8), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n270_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT8), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n266_), .A2(new_n271_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n245_), .A2(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n274_), .A2(new_n271_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(new_n244_), .A3(new_n266_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G232gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT34), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n280_), .A2(KEYINPUT35), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n276_), .A2(new_n278_), .A3(KEYINPUT71), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(KEYINPUT35), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT70), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n282_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G190gat), .B(G218gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G134gat), .B(G162gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n288_), .A2(KEYINPUT36), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(KEYINPUT36), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n285_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  OR3_X1    g094(.A1(new_n293_), .A2(KEYINPUT72), .A3(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n295_), .B1(new_n293_), .B2(KEYINPUT72), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n241_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G230gat), .A2(G233gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n224_), .A2(new_n266_), .A3(new_n277_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n275_), .A2(new_n223_), .A3(new_n222_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(KEYINPUT12), .A3(new_n302_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT12), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n275_), .A2(new_n305_), .A3(new_n223_), .A4(new_n222_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n303_), .B1(new_n307_), .B2(new_n300_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G120gat), .B(G148gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(G176gat), .B(G204gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT68), .Z(new_n316_));
  OR2_X1    g115(.A1(new_n308_), .A2(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n318_), .B1(new_n319_), .B2(KEYINPUT13), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n321_));
  NAND3_X1  g120(.A1(new_n316_), .A2(new_n317_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n299_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT23), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(G183gat), .B2(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT22), .B(G169gat), .ZN(new_n330_));
  INV_X1    g129(.A(G176gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G183gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT77), .B1(new_n334_), .B2(KEYINPUT25), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT26), .B(G190gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT25), .B(G183gat), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n335_), .B(new_n336_), .C1(new_n337_), .C2(KEYINPUT77), .ZN(new_n338_));
  INV_X1    g137(.A(G169gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(new_n331_), .A3(KEYINPUT78), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n341_), .B1(G169gat), .B2(G176gat), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n340_), .A2(new_n342_), .A3(KEYINPUT24), .A4(new_n328_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT24), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n341_), .A2(G169gat), .A3(G176gat), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT78), .B1(new_n339_), .B2(new_n331_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n344_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n338_), .A2(new_n326_), .A3(new_n343_), .A4(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n333_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350_));
  INV_X1    g149(.A(G43gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT30), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G227gat), .A2(G233gat), .ZN(new_n354_));
  INV_X1    g153(.A(G15gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n353_), .A2(new_n356_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n349_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n359_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n333_), .A2(new_n348_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n357_), .A3(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n363_), .A3(KEYINPUT79), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT31), .ZN(new_n365_));
  XOR2_X1   g164(.A(G127gat), .B(G134gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(G113gat), .B(G120gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT31), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n360_), .A2(new_n363_), .A3(KEYINPUT79), .A4(new_n369_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n365_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G141gat), .A2(G148gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G141gat), .A2(G148gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT80), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(G155gat), .A3(G162gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(KEYINPUT1), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G155gat), .A2(G162gat), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n383_), .B2(KEYINPUT1), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n384_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT81), .B1(new_n390_), .B2(new_n385_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n378_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n376_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT2), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n374_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n394_), .A2(new_n396_), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n385_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n383_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n368_), .B1(new_n392_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n381_), .B1(G155gat), .B2(G162gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n379_), .A2(KEYINPUT80), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT1), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n387_), .A3(new_n400_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n384_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n391_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n377_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n368_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n401_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n403_), .A2(KEYINPUT4), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n403_), .A2(new_n412_), .A3(KEYINPUT90), .A4(KEYINPUT4), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G225gat), .A2(G233gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n418_), .B(KEYINPUT91), .Z(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(new_n403_), .B2(KEYINPUT4), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n403_), .A2(new_n412_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(new_n419_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT93), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(new_n204_), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT92), .B(KEYINPUT0), .Z(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G29gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n428_), .B(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n422_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n431_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n420_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n424_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n373_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G228gat), .A2(G233gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n438_), .B(KEYINPUT82), .Z(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT29), .B1(new_n392_), .B2(new_n402_), .ZN(new_n440_));
  OR2_X1    g239(.A1(G197gat), .A2(G204gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G197gat), .A2(G204gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT21), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n441_), .A2(KEYINPUT21), .A3(new_n442_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G211gat), .B(G218gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT83), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n445_), .A2(new_n450_), .A3(new_n446_), .A4(new_n447_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n446_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n447_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n449_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n439_), .B1(new_n440_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n402_), .B1(new_n409_), .B2(new_n377_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n455_), .B(new_n439_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT84), .B1(new_n456_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G78gat), .B(G106gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n455_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n439_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n459_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n462_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n462_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G22gat), .B(G50gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT28), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n457_), .A2(new_n475_), .A3(new_n458_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n474_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(new_n476_), .A3(new_n473_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n465_), .A2(new_n459_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(KEYINPUT85), .A3(new_n469_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n468_), .A2(new_n472_), .A3(new_n482_), .A4(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n465_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n470_), .A2(new_n486_), .B1(new_n481_), .B2(new_n479_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT27), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT20), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n332_), .A2(KEYINPUT87), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n339_), .A2(KEYINPUT22), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT22), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G169gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n495_), .A3(new_n331_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n328_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n492_), .A2(new_n499_), .A3(new_n327_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n502_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n501_), .A2(new_n328_), .A3(new_n340_), .A4(new_n342_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n337_), .A2(new_n336_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n503_), .A2(new_n326_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n500_), .A2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n449_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n491_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT88), .B1(new_n508_), .B2(new_n362_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G226gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT19), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n455_), .A2(new_n349_), .A3(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .A4(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G8gat), .B(G36gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G64gat), .B(G92gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n500_), .A2(new_n506_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n455_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n448_), .A2(KEYINPUT83), .B1(new_n452_), .B2(new_n453_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n524_), .A2(new_n333_), .A3(new_n348_), .A4(new_n451_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(KEYINPUT20), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n512_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n516_), .A2(new_n521_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n521_), .B1(new_n516_), .B2(new_n527_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n490_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n516_), .A2(new_n521_), .A3(new_n527_), .ZN(new_n531_));
  AND4_X1   g330(.A1(KEYINPUT20), .A2(new_n523_), .A3(new_n513_), .A4(new_n525_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n509_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n533_), .B2(new_n512_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n521_), .B(KEYINPUT97), .Z(new_n535_));
  OAI211_X1 g334(.A(KEYINPUT27), .B(new_n531_), .C1(new_n534_), .C2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n437_), .A2(new_n489_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT85), .B1(new_n483_), .B2(new_n469_), .ZN(new_n540_));
  AOI211_X1 g339(.A(new_n471_), .B(new_n462_), .C1(new_n465_), .C2(new_n459_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n479_), .A2(new_n481_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n487_), .B1(new_n543_), .B2(new_n468_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n432_), .A2(new_n530_), .A3(new_n435_), .A4(new_n536_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT98), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT98), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n436_), .A2(new_n489_), .A3(new_n537_), .A4(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n516_), .A2(new_n527_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n521_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT95), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n457_), .A2(new_n411_), .ZN(new_n553_));
  AOI211_X1 g352(.A(new_n368_), .B(new_n402_), .C1(new_n409_), .C2(new_n377_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n552_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n403_), .A2(KEYINPUT95), .A3(new_n412_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n419_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n433_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n419_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n403_), .B2(KEYINPUT4), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n531_), .B(new_n551_), .C1(new_n558_), .C2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n431_), .A2(KEYINPUT33), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n434_), .A2(new_n424_), .A3(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT94), .B(KEYINPUT33), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n432_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n432_), .A2(new_n435_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n521_), .A2(KEYINPUT32), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n549_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT96), .B1(new_n534_), .B2(new_n569_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT96), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT20), .B1(new_n522_), .B2(new_n455_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n514_), .B1(new_n455_), .B2(new_n349_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n513_), .B1(new_n576_), .B2(new_n515_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n573_), .B(new_n570_), .C1(new_n577_), .C2(new_n532_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n571_), .B1(new_n572_), .B2(new_n578_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n565_), .A2(new_n567_), .B1(new_n568_), .B2(new_n579_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n546_), .B(new_n548_), .C1(new_n580_), .C2(new_n489_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n373_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n539_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n209_), .B(new_n244_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n209_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n245_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n586_), .B1(new_n209_), .B2(new_n244_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n584_), .A2(new_n586_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G113gat), .B(G141gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT76), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G169gat), .B(G197gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n590_), .A2(new_n595_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n324_), .A2(new_n583_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n204_), .A3(new_n568_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT99), .Z(new_n603_));
  OR2_X1    g402(.A1(new_n603_), .A2(KEYINPUT38), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(KEYINPUT38), .ZN(new_n605_));
  INV_X1    g404(.A(new_n293_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n583_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n607_), .A2(new_n599_), .A3(new_n323_), .A4(new_n240_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n608_), .B2(new_n436_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n604_), .A2(new_n605_), .A3(new_n609_), .ZN(G1324gat));
  OR3_X1    g409(.A1(new_n608_), .A2(KEYINPUT101), .A3(new_n537_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT101), .B1(new_n608_), .B2(new_n537_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(G8gat), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n611_), .A2(KEYINPUT39), .A3(new_n612_), .A4(G8gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n601_), .A2(new_n205_), .A3(new_n538_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT100), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT40), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n615_), .A2(KEYINPUT40), .A3(new_n616_), .A4(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1325gat));
  OAI21_X1  g422(.A(G15gat), .B1(new_n608_), .B2(new_n582_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT41), .Z(new_n625_));
  NAND3_X1  g424(.A1(new_n601_), .A2(new_n355_), .A3(new_n373_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1326gat));
  OAI21_X1  g426(.A(G22gat), .B1(new_n608_), .B2(new_n544_), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n544_), .A2(G22gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT103), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n601_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n633_), .ZN(G1327gat));
  AND2_X1   g433(.A1(new_n320_), .A2(new_n322_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n241_), .A2(new_n636_), .A3(new_n606_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT104), .B1(new_n240_), .B2(new_n293_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n635_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n583_), .A2(new_n600_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n568_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n323_), .A2(new_n599_), .A3(new_n241_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n572_), .A2(new_n578_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n571_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n563_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n422_), .A2(new_n425_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n559_), .B1(new_n423_), .B2(new_n552_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n431_), .B1(new_n651_), .B2(new_n556_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n417_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(new_n560_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n528_), .A2(new_n529_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n650_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n566_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n434_), .A2(new_n424_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(new_n431_), .ZN(new_n659_));
  OAI22_X1  g458(.A1(new_n436_), .A2(new_n648_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n436_), .A2(new_n489_), .A3(new_n537_), .ZN(new_n661_));
  AOI22_X1  g460(.A1(new_n660_), .A2(new_n544_), .B1(new_n661_), .B2(KEYINPUT98), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n373_), .B1(new_n662_), .B2(new_n548_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n645_), .B(new_n298_), .C1(new_n663_), .C2(new_n539_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n298_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n583_), .B2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n644_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT44), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n668_), .A2(G29gat), .A3(new_n568_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n644_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n581_), .A2(new_n582_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n539_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n645_), .B1(new_n673_), .B2(new_n298_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n583_), .A2(KEYINPUT43), .A3(new_n665_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n670_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n643_), .B1(new_n669_), .B2(new_n678_), .ZN(G1328gat));
  NOR2_X1   g478(.A1(new_n537_), .A2(G36gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n639_), .A2(new_n640_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT106), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n639_), .A2(new_n683_), .A3(new_n640_), .A4(new_n680_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n682_), .A2(KEYINPUT45), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT45), .B1(new_n682_), .B2(new_n684_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n537_), .B1(new_n667_), .B2(KEYINPUT44), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n678_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n690_), .B2(G36gat), .ZN(new_n691_));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT105), .B(new_n692_), .C1(new_n689_), .C2(new_n678_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n687_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT46), .B(new_n687_), .C1(new_n691_), .C2(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1329gat));
  OAI21_X1  g497(.A(new_n351_), .B1(new_n641_), .B2(new_n582_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n668_), .A2(G43gat), .A3(new_n373_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n678_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g502(.A(G50gat), .B1(new_n642_), .B2(new_n489_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n668_), .A2(G50gat), .A3(new_n489_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n678_), .ZN(G1331gat));
  NAND4_X1  g505(.A1(new_n607_), .A2(new_n600_), .A3(new_n635_), .A4(new_n240_), .ZN(new_n707_));
  XOR2_X1   g506(.A(KEYINPUT109), .B(G57gat), .Z(new_n708_));
  NOR3_X1   g507(.A1(new_n707_), .A2(new_n436_), .A3(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n583_), .A2(new_n599_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n635_), .A3(new_n299_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT107), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n568_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n714_), .A2(KEYINPUT108), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(KEYINPUT108), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n709_), .B1(new_n715_), .B2(new_n716_), .ZN(G1332gat));
  OR3_X1    g516(.A1(new_n712_), .A2(G64gat), .A3(new_n537_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G64gat), .B1(new_n707_), .B2(new_n537_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(KEYINPUT48), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(KEYINPUT48), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT110), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n718_), .B(new_n724_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n707_), .B2(new_n582_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT49), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n582_), .A2(G71gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n712_), .B2(new_n729_), .ZN(G1334gat));
  OAI21_X1  g529(.A(G78gat), .B1(new_n707_), .B2(new_n544_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n544_), .A2(G78gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n712_), .B2(new_n733_), .ZN(G1335gat));
  NOR2_X1   g533(.A1(new_n674_), .A2(new_n675_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n635_), .A2(new_n600_), .A3(new_n241_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT111), .Z(new_n738_));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n436_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n323_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n710_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n247_), .A3(new_n568_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1336gat));
  OAI21_X1  g542(.A(G92gat), .B1(new_n738_), .B2(new_n537_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n741_), .A2(new_n248_), .A3(new_n538_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1337gat));
  AOI21_X1  g545(.A(new_n256_), .B1(new_n737_), .B2(new_n373_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n741_), .A2(new_n373_), .A3(new_n261_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(KEYINPUT112), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n749_), .B(new_n751_), .Z(G1338gat));
  NAND3_X1  g551(.A1(new_n741_), .A2(new_n257_), .A3(new_n489_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n257_), .B1(new_n737_), .B2(new_n489_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(KEYINPUT52), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(KEYINPUT52), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT53), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n756_), .A2(KEYINPUT52), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n758_), .A3(new_n762_), .A4(new_n755_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765_));
  INV_X1    g564(.A(new_n300_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT55), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n766_), .B(new_n768_), .C1(new_n304_), .C2(new_n306_), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n767_), .A2(KEYINPUT55), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n307_), .A2(new_n300_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(new_n768_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n304_), .A2(new_n766_), .A3(new_n306_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT114), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n304_), .A2(new_n775_), .A3(new_n766_), .A4(new_n306_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n765_), .B1(new_n772_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n771_), .A2(new_n768_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n769_), .ZN(new_n780_));
  AND4_X1   g579(.A1(new_n765_), .A2(new_n777_), .A3(new_n779_), .A4(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n313_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n584_), .A2(new_n585_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n585_), .B1(new_n209_), .B2(new_n244_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n588_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n784_), .A2(new_n594_), .A3(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n596_), .A2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT117), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n313_), .C1(new_n778_), .C2(new_n781_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n783_), .A2(new_n316_), .A3(new_n790_), .A4(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n665_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n793_), .A2(KEYINPUT119), .A3(new_n794_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT119), .B1(new_n793_), .B2(new_n794_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n783_), .A2(new_n599_), .A3(new_n316_), .A4(new_n792_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n790_), .A2(new_n318_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n606_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT57), .ZN(new_n804_));
  XNOR2_X1  g603(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n241_), .B1(new_n800_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808_));
  INV_X1    g607(.A(new_n324_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n600_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n324_), .A2(KEYINPUT54), .A3(new_n599_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n807_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n537_), .A2(new_n568_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n582_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n814_), .A2(KEYINPUT59), .A3(new_n544_), .A4(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n801_), .A2(new_n802_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n805_), .B1(new_n818_), .B2(new_n293_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n820_), .B(new_n606_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n779_), .A2(new_n780_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n777_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT116), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n772_), .A2(new_n765_), .A3(new_n777_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n314_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n316_), .B1(new_n828_), .B2(new_n791_), .ZN(new_n829_));
  AOI211_X1 g628(.A(KEYINPUT56), .B(new_n314_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n829_), .A2(new_n789_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n823_), .B1(new_n831_), .B2(KEYINPUT58), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n795_), .B1(new_n832_), .B2(new_n797_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n240_), .B1(new_n822_), .B2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n544_), .B(new_n816_), .C1(new_n834_), .C2(new_n812_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n817_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(G113gat), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n599_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n840_), .B2(new_n839_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n835_), .A2(new_n600_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n838_), .A2(new_n842_), .B1(new_n843_), .B2(new_n839_), .ZN(G1340gat));
  NOR2_X1   g643(.A1(new_n834_), .A2(new_n812_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n489_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n847_));
  AOI21_X1  g646(.A(G120gat), .B1(new_n635_), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n847_), .B2(G120gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n846_), .A2(new_n816_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n323_), .B1(new_n817_), .B2(new_n837_), .ZN(new_n851_));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(G1341gat));
  AOI21_X1  g652(.A(new_n241_), .B1(new_n817_), .B2(new_n837_), .ZN(new_n854_));
  INV_X1    g653(.A(G127gat), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n240_), .A2(new_n855_), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n854_), .A2(new_n855_), .B1(new_n835_), .B2(new_n856_), .ZN(G1342gat));
  XNOR2_X1  g656(.A(KEYINPUT121), .B(G134gat), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n665_), .A2(new_n858_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n835_), .A2(new_n293_), .ZN(new_n860_));
  INV_X1    g659(.A(G134gat), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n838_), .A2(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(G1343gat));
  NAND2_X1  g661(.A1(new_n582_), .A2(new_n489_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n815_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n814_), .A2(new_n599_), .A3(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT122), .B(G141gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1344gat));
  NAND3_X1  g666(.A1(new_n814_), .A2(new_n635_), .A3(new_n864_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g668(.A1(new_n814_), .A2(new_n240_), .A3(new_n864_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT61), .B(G155gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1346gat));
  NAND2_X1  g671(.A1(new_n814_), .A2(new_n864_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G162gat), .B1(new_n873_), .B2(new_n665_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n293_), .A2(G162gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n873_), .B2(new_n875_), .ZN(G1347gat));
  NOR3_X1   g675(.A1(new_n437_), .A2(new_n600_), .A3(new_n537_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n544_), .B(new_n877_), .C1(new_n834_), .C2(new_n812_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G169gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT123), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n881_), .A3(G169gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(KEYINPUT62), .A3(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n437_), .A2(new_n537_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n544_), .B(new_n884_), .C1(new_n834_), .C2(new_n812_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n599_), .A2(new_n330_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT124), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n881_), .B1(new_n878_), .B2(G169gat), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n883_), .A2(new_n891_), .ZN(G1348gat));
  NOR2_X1   g691(.A1(new_n885_), .A2(new_n323_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n331_), .ZN(G1349gat));
  NOR3_X1   g693(.A1(new_n885_), .A2(new_n337_), .A3(new_n241_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n885_), .A2(new_n241_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n334_), .B2(new_n896_), .ZN(G1350gat));
  NAND4_X1  g696(.A1(new_n846_), .A2(new_n336_), .A3(new_n606_), .A4(new_n884_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n814_), .A2(new_n544_), .A3(new_n298_), .A4(new_n884_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT125), .B1(new_n899_), .B2(G190gat), .ZN(new_n900_));
  OAI211_X1 g699(.A(KEYINPUT125), .B(G190gat), .C1(new_n885_), .C2(new_n665_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n898_), .B1(new_n900_), .B2(new_n902_), .ZN(G1351gat));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n863_), .A2(new_n568_), .A3(new_n537_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n814_), .A2(new_n599_), .A3(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(G197gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n904_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n905_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n845_), .A2(new_n909_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n910_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n599_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n906_), .A2(new_n907_), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n908_), .A2(new_n911_), .A3(new_n912_), .ZN(G1352gat));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n635_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g714(.A(KEYINPUT63), .B(G211gat), .C1(new_n910_), .C2(new_n240_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT63), .B(G211gat), .Z(new_n917_));
  AND3_X1   g716(.A1(new_n910_), .A2(new_n240_), .A3(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1354gat));
  AOI21_X1  g718(.A(G218gat), .B1(new_n910_), .B2(new_n606_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n298_), .A2(G218gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n910_), .B2(new_n922_), .ZN(G1355gat));
endmodule


