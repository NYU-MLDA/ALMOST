//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n966_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_,
    new_n983_, new_n985_, new_n986_, new_n987_, new_n988_, new_n990_,
    new_n991_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1022_, new_n1023_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G71gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT30), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT22), .B(G169gat), .ZN(new_n209_));
  INV_X1    g008(.A(G176gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT83), .ZN(new_n212_));
  INV_X1    g011(.A(G169gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT22), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT22), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G169gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n216_), .A3(new_n210_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(new_n207_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT83), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(new_n224_), .A3(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n212_), .A2(new_n220_), .A3(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n223_), .A2(new_n224_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n213_), .A2(new_n210_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n230_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT81), .B1(new_n225_), .B2(KEYINPUT25), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT81), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(G183gat), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n226_), .A2(KEYINPUT26), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT26), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G190gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n225_), .A2(KEYINPUT25), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n240_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT82), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n239_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n235_), .A2(new_n238_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n240_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT82), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n234_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n206_), .B1(new_n229_), .B2(new_n250_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n230_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n245_), .B1(new_n239_), .B2(new_n244_), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT82), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n218_), .A2(new_n219_), .B1(new_n230_), .B2(new_n227_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n212_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n257_), .A3(KEYINPUT30), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT84), .B(G43gat), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n251_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n259_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n205_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G134gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(G127gat), .ZN(new_n264_));
  INV_X1    g063(.A(G127gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G134gat), .ZN(new_n266_));
  INV_X1    g065(.A(G120gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G113gat), .ZN(new_n268_));
  INV_X1    g067(.A(G113gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G120gat), .ZN(new_n270_));
  AND4_X1   g069(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .A4(new_n270_), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n264_), .A2(new_n266_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT85), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT85), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n264_), .A2(new_n266_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n268_), .A2(new_n270_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT31), .ZN(new_n279_));
  INV_X1    g078(.A(G99gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n251_), .A2(new_n258_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n259_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n251_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n205_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n262_), .A2(new_n281_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n281_), .B1(new_n287_), .B2(new_n262_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G8gat), .B(G36gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT18), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G64gat), .B(G92gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  INV_X1    g095(.A(G218gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G211gat), .ZN(new_n298_));
  INV_X1    g097(.A(G211gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G218gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G197gat), .ZN(new_n302_));
  INV_X1    g101(.A(G204gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G197gat), .A2(G204gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n301_), .B1(KEYINPUT91), .B2(new_n306_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n298_), .A2(new_n300_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT21), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n298_), .A2(new_n300_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n305_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G197gat), .A2(G204gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT91), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT21), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT25), .B(G183gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT26), .B(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n320_), .A2(new_n230_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT94), .B1(new_n211_), .B2(new_n228_), .ZN(new_n322_));
  AND4_X1   g121(.A1(KEYINPUT94), .A2(new_n228_), .A3(new_n207_), .A4(new_n217_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n310_), .A2(new_n313_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n301_), .A2(new_n306_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n314_), .B1(new_n327_), .B2(KEYINPUT21), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n317_), .A2(new_n329_), .A3(KEYINPUT20), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT19), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n330_), .A2(KEYINPUT95), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT95), .B1(new_n330_), .B2(new_n332_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n246_), .A2(new_n249_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n336_), .A2(new_n252_), .B1(new_n256_), .B2(new_n212_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT20), .B1(new_n337_), .B2(new_n316_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n332_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT96), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n228_), .A2(new_n217_), .A3(new_n207_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT94), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n211_), .A2(KEYINPUT94), .A3(new_n228_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n344_), .A2(new_n345_), .B1(new_n252_), .B2(new_n320_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n332_), .B1(new_n346_), .B2(new_n316_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n255_), .A2(new_n257_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n328_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT96), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .A4(KEYINPUT20), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n341_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n296_), .B1(new_n335_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n330_), .A2(new_n332_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT95), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n330_), .A2(KEYINPUT95), .A3(new_n332_), .ZN(new_n357_));
  AND4_X1   g156(.A1(new_n296_), .A2(new_n352_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n292_), .B1(new_n353_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT27), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n316_), .A2(new_n321_), .A3(new_n342_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n332_), .B1(new_n338_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n332_), .B2(new_n330_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n296_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n360_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n352_), .A2(new_n356_), .A3(new_n296_), .A4(new_n357_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n370_), .A2(KEYINPUT86), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(KEYINPUT86), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n371_), .A2(new_n372_), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  OR2_X1    g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT87), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT87), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(G155gat), .A3(G162gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT1), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n374_), .B(new_n380_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n383_));
  AOI211_X1 g182(.A(KEYINPUT88), .B(new_n379_), .C1(new_n376_), .C2(new_n378_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n373_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n370_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT2), .ZN(new_n388_));
  INV_X1    g187(.A(G141gat), .ZN(new_n389_));
  INV_X1    g188(.A(G148gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI22_X1  g190(.A1(KEYINPUT89), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n387_), .A2(new_n391_), .A3(new_n392_), .A4(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n376_), .A2(new_n378_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n374_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n385_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n278_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n271_), .A2(new_n272_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n385_), .A2(new_n396_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(KEYINPUT4), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n396_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n395_), .A2(KEYINPUT1), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT88), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n380_), .A2(new_n374_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n381_), .A2(new_n382_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n403_), .B1(new_n408_), .B2(new_n373_), .ZN(new_n409_));
  NOR4_X1   g208(.A1(new_n409_), .A2(KEYINPUT97), .A3(KEYINPUT4), .A4(new_n278_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT97), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n278_), .B1(new_n385_), .B2(new_n396_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n369_), .B(new_n402_), .C1(new_n410_), .C2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT98), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n397_), .A2(new_n413_), .A3(new_n398_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT97), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n412_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT98), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n369_), .A4(new_n402_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G1gat), .B(G29gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G85gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT0), .B(G57gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n401_), .B(new_n368_), .C1(new_n409_), .C2(new_n278_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT99), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT99), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n399_), .A2(new_n430_), .A3(new_n368_), .A4(new_n401_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n416_), .A2(new_n422_), .A3(new_n427_), .A4(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n432_), .B1(new_n415_), .B2(KEYINPUT98), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n402_), .A2(new_n369_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n421_), .B1(new_n435_), .B2(new_n420_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n426_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n359_), .A2(new_n367_), .A3(new_n433_), .A4(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G22gat), .B(G50gat), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT29), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n409_), .B2(new_n443_), .ZN(new_n444_));
  AND4_X1   g243(.A1(new_n443_), .A2(new_n385_), .A3(new_n396_), .A4(new_n442_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n440_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n441_), .B1(new_n397_), .B2(KEYINPUT29), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n409_), .A2(new_n443_), .A3(new_n442_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n439_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT93), .B1(new_n450_), .B2(KEYINPUT92), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n328_), .B1(new_n409_), .B2(new_n443_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(G78gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G106gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n328_), .B(new_n457_), .C1(new_n409_), .C2(new_n443_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n450_), .B2(KEYINPUT92), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT93), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n446_), .A2(new_n449_), .A3(new_n463_), .A4(new_n464_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n451_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n462_), .B1(new_n451_), .B2(new_n465_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n290_), .B1(new_n438_), .B2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n353_), .A2(new_n358_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n433_), .A2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n426_), .A2(new_n471_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n416_), .A2(new_n422_), .A3(new_n432_), .A4(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n420_), .A2(new_n368_), .A3(new_n402_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n399_), .A2(new_n369_), .A3(new_n401_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n426_), .A3(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n470_), .A2(new_n472_), .A3(new_n474_), .A4(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n437_), .A2(new_n433_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n363_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n352_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n296_), .A2(KEYINPUT32), .ZN(new_n482_));
  MUX2_X1   g281(.A(new_n480_), .B(new_n481_), .S(new_n482_), .Z(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n467_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n451_), .A2(new_n462_), .A3(new_n465_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n478_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n359_), .A2(new_n367_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(new_n468_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n290_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n479_), .A2(new_n491_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n469_), .A2(new_n488_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G120gat), .B(G148gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT5), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G176gat), .B(G204gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  XOR2_X1   g296(.A(G85gat), .B(G92gat), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT9), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT10), .B(G99gat), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n456_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT6), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(G99gat), .A3(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT64), .B(G85gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT9), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(G92gat), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n499_), .A2(new_n501_), .A3(new_n506_), .A4(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT8), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n503_), .A2(new_n505_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT65), .ZN(new_n513_));
  NOR2_X1   g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT7), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n506_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n511_), .B1(new_n518_), .B2(new_n498_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n515_), .A2(new_n506_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n520_), .A2(new_n511_), .A3(new_n498_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n510_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n524_));
  XOR2_X1   g323(.A(G71gat), .B(G78gat), .Z(new_n525_));
  OR2_X1    g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT68), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n525_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n526_), .B(new_n527_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n526_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n532_), .A2(KEYINPUT68), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n522_), .B(KEYINPUT12), .C1(new_n531_), .C2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n518_), .A2(new_n498_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT8), .ZN(new_n536_));
  INV_X1    g335(.A(new_n521_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(new_n532_), .A3(new_n510_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n532_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n522_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(KEYINPUT69), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n544_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT69), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n541_), .A2(new_n545_), .A3(new_n548_), .A4(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n539_), .A2(KEYINPUT66), .ZN(new_n551_));
  INV_X1    g350(.A(new_n522_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT66), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n532_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n543_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n549_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(KEYINPUT67), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT67), .B1(new_n555_), .B2(new_n556_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n497_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n497_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n561_), .A2(new_n550_), .A3(new_n557_), .A4(new_n562_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n560_), .A2(new_n563_), .A3(KEYINPUT13), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT13), .B1(new_n560_), .B2(new_n563_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT80), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G113gat), .B(G141gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G169gat), .B(G197gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  XNOR2_X1  g369(.A(G1gat), .B(G8gat), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT75), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G15gat), .B(G22gat), .ZN(new_n574_));
  INV_X1    g373(.A(G1gat), .ZN(new_n575_));
  INV_X1    g374(.A(G8gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT14), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n573_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n571_), .B(KEYINPUT75), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G29gat), .B(G36gat), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT70), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT70), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G43gat), .B(G50gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n591_), .A2(KEYINPUT15), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT15), .B1(new_n591_), .B2(new_n592_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n584_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT79), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n581_), .A2(new_n578_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n573_), .A2(new_n579_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n592_), .B(new_n591_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .A4(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n591_), .A2(new_n592_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n600_), .A3(KEYINPUT78), .ZN(new_n604_));
  INV_X1    g403(.A(new_n597_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT78), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n584_), .A2(new_n606_), .A3(new_n602_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n601_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n595_), .A2(new_n597_), .A3(new_n600_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT79), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n570_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  AND4_X1   g411(.A1(new_n611_), .A2(new_n608_), .A3(new_n601_), .A4(new_n570_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n567_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n570_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n611_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n601_), .A2(new_n608_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n609_), .A2(new_n611_), .A3(new_n570_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(KEYINPUT80), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n566_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n493_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n602_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n629_), .B(new_n510_), .C1(new_n519_), .C2(new_n521_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT34), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT35), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n593_), .A2(new_n594_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n630_), .B(new_n635_), .C1(new_n552_), .C2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n594_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n591_), .A2(KEYINPUT15), .A3(new_n592_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT71), .B1(new_n640_), .B2(new_n522_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n633_), .A2(new_n634_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n637_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(new_n522_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n645_), .A2(KEYINPUT71), .A3(new_n642_), .A4(new_n630_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n628_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT72), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n626_), .B(KEYINPUT36), .Z(new_n649_));
  NAND3_X1  g448(.A1(new_n644_), .A2(new_n646_), .A3(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n644_), .A2(new_n646_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT72), .B1(new_n653_), .B2(new_n627_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT72), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n655_), .B(new_n628_), .C1(new_n644_), .C2(new_n646_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n650_), .A2(KEYINPUT73), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT73), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n644_), .A2(new_n659_), .A3(new_n646_), .A4(new_n649_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT37), .B1(new_n657_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n652_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(G127gat), .B(G155gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT16), .ZN(new_n666_));
  XNOR2_X1  g465(.A(G183gat), .B(G211gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT17), .ZN(new_n669_));
  NAND2_X1  g468(.A1(G231gat), .A2(G233gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n580_), .A2(new_n582_), .A3(G231gat), .A4(G233gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n532_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n542_), .A3(new_n672_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n668_), .A2(KEYINPUT17), .ZN(new_n676_));
  AND4_X1   g475(.A1(new_n669_), .A2(new_n674_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n673_), .A2(KEYINPUT76), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT76), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n671_), .A2(new_n679_), .A3(new_n672_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n681_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n669_), .B(KEYINPUT77), .Z(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n677_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n664_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n623_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT101), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(new_n575_), .A3(new_n479_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT38), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT102), .B1(new_n648_), .B2(new_n650_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT102), .B(new_n650_), .C1(new_n654_), .C2(new_n656_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  NOR4_X1   g496(.A1(new_n493_), .A2(new_n622_), .A3(new_n697_), .A4(new_n687_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n575_), .B1(new_n698_), .B2(new_n479_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n693_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n691_), .A2(new_n692_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT103), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT103), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n702_), .B2(new_n703_), .ZN(G1324gat));
  AOI21_X1  g503(.A(new_n576_), .B1(new_n698_), .B2(new_n489_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT39), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n690_), .A2(new_n576_), .A3(new_n489_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1325gat));
  NAND3_X1  g511(.A1(new_n690_), .A2(new_n203_), .A3(new_n290_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n714_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n203_), .B1(new_n698_), .B2(new_n290_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT41), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n715_), .A2(new_n716_), .A3(new_n718_), .ZN(G1326gat));
  INV_X1    g518(.A(G22gat), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n487_), .B(KEYINPUT106), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n698_), .B2(new_n721_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT107), .Z(new_n723_));
  INV_X1    g522(.A(KEYINPUT42), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n724_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n690_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(G1327gat));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n694_), .A2(new_n696_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(new_n686_), .ZN(new_n731_));
  OAI211_X1 g530(.A(KEYINPUT110), .B(new_n687_), .C1(new_n694_), .C2(new_n696_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(new_n623_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G29gat), .B1(new_n734_), .B2(new_n479_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n438_), .A2(new_n468_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n488_), .A2(new_n738_), .A3(new_n491_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n489_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n479_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n740_), .A2(new_n487_), .A3(new_n741_), .A4(new_n290_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n663_), .B1(new_n739_), .B2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n737_), .B1(new_n743_), .B2(KEYINPUT108), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n745_), .B(KEYINPUT43), .C1(new_n493_), .C2(new_n663_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n622_), .A2(new_n686_), .ZN(new_n748_));
  AND4_X1   g547(.A1(new_n736_), .A2(new_n747_), .A3(KEYINPUT44), .A4(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n748_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n736_), .B1(new_n751_), .B2(KEYINPUT44), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n749_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n481_), .A2(new_n364_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n291_), .B1(new_n755_), .B2(new_n366_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n367_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n479_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n491_), .B1(new_n758_), .B2(new_n487_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n478_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n742_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n664_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT43), .B1(new_n762_), .B2(new_n745_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n746_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n748_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n753_), .B1(new_n754_), .B2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n479_), .A2(G29gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n735_), .B1(new_n766_), .B2(new_n767_), .ZN(G1328gat));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT112), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n740_), .B1(new_n765_), .B2(new_n754_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n749_), .B2(new_n752_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G36gat), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n740_), .A2(G36gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n733_), .A2(new_n623_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT45), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n733_), .A2(new_n779_), .A3(new_n623_), .A4(new_n776_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n778_), .A2(new_n780_), .B1(KEYINPUT112), .B2(new_n770_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n772_), .B1(new_n775_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n781_), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n771_), .B(new_n783_), .C1(new_n774_), .C2(G36gat), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1329gat));
  AND2_X1   g584(.A1(new_n290_), .A2(G43gat), .ZN(new_n786_));
  OAI221_X1 g585(.A(new_n786_), .B1(KEYINPUT44), .B2(new_n751_), .C1(new_n749_), .C2(new_n752_), .ZN(new_n787_));
  AOI21_X1  g586(.A(G43gat), .B1(new_n734_), .B2(new_n290_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n787_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT47), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1330gat));
  AOI21_X1  g594(.A(G50gat), .B1(new_n734_), .B2(new_n721_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n468_), .A2(G50gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n766_), .B2(new_n797_), .ZN(G1331gat));
  NOR2_X1   g597(.A1(new_n493_), .A2(new_n621_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n566_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(new_n688_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(G57gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n479_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n614_), .A2(new_n686_), .A3(new_n620_), .ZN(new_n804_));
  NOR4_X1   g603(.A1(new_n493_), .A2(new_n697_), .A3(new_n566_), .A4(new_n804_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT114), .Z(new_n806_));
  AND2_X1   g605(.A1(new_n806_), .A2(new_n479_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n807_), .B2(new_n802_), .ZN(G1332gat));
  INV_X1    g607(.A(G64gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n801_), .A2(new_n809_), .A3(new_n489_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT48), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n806_), .A2(new_n489_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(G64gat), .ZN(new_n813_));
  AOI211_X1 g612(.A(KEYINPUT48), .B(new_n809_), .C1(new_n806_), .C2(new_n489_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(G1333gat));
  INV_X1    g614(.A(G71gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n801_), .A2(new_n816_), .A3(new_n290_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n806_), .A2(new_n290_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(G71gat), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT49), .B(new_n816_), .C1(new_n806_), .C2(new_n290_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n817_), .B1(new_n820_), .B2(new_n821_), .ZN(G1334gat));
  NAND3_X1  g621(.A1(new_n801_), .A2(new_n454_), .A3(new_n721_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n806_), .A2(new_n721_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(G78gat), .ZN(new_n826_));
  AOI211_X1 g625(.A(KEYINPUT50), .B(new_n454_), .C1(new_n806_), .C2(new_n721_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n823_), .B1(new_n826_), .B2(new_n827_), .ZN(G1335gat));
  AOI21_X1  g627(.A(new_n566_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n799_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G85gat), .B1(new_n831_), .B2(new_n479_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n566_), .A2(new_n686_), .A3(new_n621_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n747_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT115), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n747_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n834_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n479_), .A2(new_n507_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n832_), .B1(new_n839_), .B2(new_n840_), .ZN(G1336gat));
  INV_X1    g640(.A(G92gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n839_), .B2(new_n489_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n830_), .A2(G92gat), .A3(new_n740_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1337gat));
  NAND2_X1  g644(.A1(new_n839_), .A2(new_n290_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G99gat), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n290_), .A2(new_n500_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n830_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n848_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n280_), .B1(new_n839_), .B2(new_n290_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT51), .B1(new_n853_), .B2(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1338gat));
  NAND2_X1  g654(.A1(new_n833_), .A2(new_n468_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G106gat), .B1(new_n835_), .B2(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n857_), .A2(KEYINPUT52), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(KEYINPUT52), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n468_), .A2(new_n456_), .ZN(new_n860_));
  OAI22_X1  g659(.A1(new_n858_), .A2(new_n859_), .B1(new_n830_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT53), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n863_));
  OAI221_X1 g662(.A(new_n863_), .B1(new_n830_), .B2(new_n860_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1339gat));
  NOR4_X1   g664(.A1(new_n489_), .A2(new_n741_), .A3(new_n468_), .A4(new_n491_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n621_), .A2(new_n563_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n550_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n541_), .A2(new_n548_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n545_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n556_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n868_), .B1(new_n871_), .B2(KEYINPUT55), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n869_), .A2(new_n870_), .A3(new_n873_), .A4(new_n556_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n497_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n540_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n549_), .B1(new_n878_), .B2(new_n545_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n550_), .B1(new_n879_), .B2(new_n873_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n871_), .A2(new_n868_), .A3(KEYINPUT55), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(KEYINPUT56), .A3(new_n497_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n867_), .B1(new_n877_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n560_), .A2(new_n563_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n604_), .A2(new_n597_), .A3(new_n607_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n595_), .A2(new_n605_), .A3(new_n600_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n615_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n885_), .A2(new_n619_), .A3(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n730_), .B1(new_n884_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n563_), .A2(new_n619_), .A3(new_n888_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT56), .B1(new_n882_), .B2(new_n497_), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n876_), .B(new_n562_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  OAI221_X1 g697(.A(new_n893_), .B1(KEYINPUT119), .B2(KEYINPUT58), .C1(new_n894_), .C2(new_n895_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n898_), .A2(new_n899_), .A3(new_n664_), .ZN(new_n900_));
  OAI211_X1 g699(.A(KEYINPUT57), .B(new_n730_), .C1(new_n884_), .C2(new_n889_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n892_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n902_), .A2(new_n687_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT117), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n804_), .A2(new_n905_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n614_), .A2(new_n686_), .A3(new_n620_), .A4(KEYINPUT116), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n904_), .B1(new_n908_), .B2(new_n566_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT13), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n885_), .A2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n560_), .A2(new_n563_), .A3(KEYINPUT13), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n911_), .A2(new_n906_), .A3(new_n912_), .A4(new_n907_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(KEYINPUT117), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n663_), .B1(new_n909_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n908_), .A2(new_n904_), .A3(new_n566_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n913_), .A2(KEYINPUT117), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n664_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(KEYINPUT54), .B1(new_n921_), .B2(KEYINPUT118), .ZN(new_n922_));
  AOI211_X1 g721(.A(new_n916_), .B(new_n664_), .C1(new_n919_), .C2(new_n920_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n918_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n866_), .B1(new_n903_), .B2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(new_n269_), .A3(new_n621_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n621_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n917_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n923_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n902_), .A2(new_n687_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(new_n934_), .A3(new_n918_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n935_), .A2(KEYINPUT59), .A3(new_n866_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n928_), .B1(new_n930_), .B2(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n927_), .B1(new_n937_), .B2(new_n269_), .ZN(G1340gat));
  XNOR2_X1  g737(.A(KEYINPUT120), .B(G120gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n939_), .B1(new_n566_), .B2(KEYINPUT60), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n926_), .B(new_n940_), .C1(KEYINPUT60), .C2(new_n939_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n566_), .B1(new_n930_), .B2(new_n936_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n939_), .ZN(G1341gat));
  AOI21_X1  g742(.A(G127gat), .B1(new_n926_), .B2(new_n686_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n930_), .A2(new_n936_), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT121), .B(G127gat), .Z(new_n946_));
  NAND2_X1  g745(.A1(new_n686_), .A2(new_n946_), .ZN(new_n947_));
  XOR2_X1   g746(.A(new_n947_), .B(KEYINPUT122), .Z(new_n948_));
  AOI21_X1  g747(.A(new_n944_), .B1(new_n945_), .B2(new_n948_), .ZN(G1342gat));
  AOI21_X1  g748(.A(G134gat), .B1(new_n926_), .B2(new_n697_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n664_), .A2(G134gat), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(KEYINPUT123), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n950_), .B1(new_n945_), .B2(new_n952_), .ZN(G1343gat));
  NOR2_X1   g752(.A1(new_n903_), .A2(new_n924_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n487_), .A2(new_n290_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n955_), .A2(new_n740_), .A3(new_n479_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n954_), .A2(new_n928_), .A3(new_n956_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(new_n389_), .ZN(G1344gat));
  NOR3_X1   g757(.A1(new_n954_), .A2(new_n566_), .A3(new_n956_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(new_n390_), .ZN(G1345gat));
  NOR3_X1   g759(.A1(new_n954_), .A2(new_n687_), .A3(new_n956_), .ZN(new_n961_));
  XOR2_X1   g760(.A(KEYINPUT61), .B(G155gat), .Z(new_n962_));
  XNOR2_X1  g761(.A(new_n961_), .B(new_n962_), .ZN(G1346gat));
  NOR2_X1   g762(.A1(new_n954_), .A2(new_n956_), .ZN(new_n964_));
  INV_X1    g763(.A(G162gat), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n964_), .A2(new_n965_), .A3(new_n697_), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n954_), .A2(new_n663_), .A3(new_n956_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n966_), .B1(new_n965_), .B2(new_n967_), .ZN(G1347gat));
  NOR2_X1   g767(.A1(new_n740_), .A2(new_n479_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(new_n290_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n970_), .A2(new_n721_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n935_), .A2(new_n621_), .A3(new_n971_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(G169gat), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n973_), .A2(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n971_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n954_), .A2(new_n976_), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n977_), .A2(new_n209_), .A3(new_n621_), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n972_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n975_), .A2(new_n978_), .A3(new_n979_), .ZN(G1348gat));
  NAND2_X1  g779(.A1(new_n977_), .A2(new_n800_), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n954_), .A2(new_n468_), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n970_), .A2(new_n566_), .A3(new_n210_), .ZN(new_n983_));
  AOI22_X1  g782(.A1(new_n981_), .A2(new_n210_), .B1(new_n982_), .B2(new_n983_), .ZN(G1349gat));
  NOR2_X1   g783(.A1(new_n970_), .A2(new_n687_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n982_), .A2(new_n985_), .ZN(new_n986_));
  OR2_X1    g785(.A1(new_n687_), .A2(new_n318_), .ZN(new_n987_));
  INV_X1    g786(.A(new_n987_), .ZN(new_n988_));
  AOI22_X1  g787(.A1(new_n986_), .A2(new_n225_), .B1(new_n977_), .B2(new_n988_), .ZN(G1350gat));
  NAND3_X1  g788(.A1(new_n977_), .A2(new_n319_), .A3(new_n697_), .ZN(new_n990_));
  NOR3_X1   g789(.A1(new_n954_), .A2(new_n663_), .A3(new_n976_), .ZN(new_n991_));
  OAI21_X1  g790(.A(new_n990_), .B1(new_n226_), .B2(new_n991_), .ZN(G1351gat));
  INV_X1    g791(.A(new_n969_), .ZN(new_n993_));
  INV_X1    g792(.A(new_n955_), .ZN(new_n994_));
  NOR2_X1   g793(.A1(new_n993_), .A2(new_n994_), .ZN(new_n995_));
  INV_X1    g794(.A(new_n995_), .ZN(new_n996_));
  NOR3_X1   g795(.A1(new_n921_), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n997_));
  AOI21_X1  g796(.A(new_n997_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n996_), .B1(new_n998_), .B2(new_n934_), .ZN(new_n999_));
  NAND2_X1  g798(.A1(new_n999_), .A2(new_n621_), .ZN(new_n1000_));
  XNOR2_X1  g799(.A(new_n1000_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g800(.A1(new_n999_), .A2(new_n800_), .ZN(new_n1002_));
  AND2_X1   g801(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n1003_));
  NOR2_X1   g802(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n1004_));
  OAI21_X1  g803(.A(new_n1002_), .B1(new_n1003_), .B2(new_n1004_), .ZN(new_n1005_));
  OAI21_X1  g804(.A(new_n1005_), .B1(new_n1002_), .B2(new_n1003_), .ZN(G1353gat));
  INV_X1    g805(.A(KEYINPUT63), .ZN(new_n1007_));
  OAI21_X1  g806(.A(new_n686_), .B1(new_n1007_), .B2(new_n299_), .ZN(new_n1008_));
  INV_X1    g807(.A(new_n1008_), .ZN(new_n1009_));
  OAI211_X1 g808(.A(new_n995_), .B(new_n1009_), .C1(new_n903_), .C2(new_n924_), .ZN(new_n1010_));
  NOR2_X1   g809(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1011_));
  XNOR2_X1  g810(.A(new_n1011_), .B(KEYINPUT125), .ZN(new_n1012_));
  NAND2_X1  g811(.A1(new_n1010_), .A2(new_n1012_), .ZN(new_n1013_));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1014_));
  NAND2_X1  g813(.A1(new_n1013_), .A2(new_n1014_), .ZN(new_n1015_));
  NAND3_X1  g814(.A1(new_n1010_), .A2(KEYINPUT127), .A3(new_n1012_), .ZN(new_n1016_));
  OAI21_X1  g815(.A(KEYINPUT126), .B1(new_n1010_), .B2(new_n1012_), .ZN(new_n1017_));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1018_));
  INV_X1    g817(.A(new_n1012_), .ZN(new_n1019_));
  NAND4_X1  g818(.A1(new_n999_), .A2(new_n1018_), .A3(new_n1019_), .A4(new_n1009_), .ZN(new_n1020_));
  AOI22_X1  g819(.A1(new_n1015_), .A2(new_n1016_), .B1(new_n1017_), .B2(new_n1020_), .ZN(G1354gat));
  NAND3_X1  g820(.A1(new_n999_), .A2(new_n297_), .A3(new_n697_), .ZN(new_n1022_));
  NOR3_X1   g821(.A1(new_n954_), .A2(new_n663_), .A3(new_n996_), .ZN(new_n1023_));
  OAI21_X1  g822(.A(new_n1022_), .B1(new_n1023_), .B2(new_n297_), .ZN(G1355gat));
endmodule


