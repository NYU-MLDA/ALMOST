//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n202_), .A2(new_n203_), .ZN(new_n205_));
  MUX2_X1   g004(.A(new_n204_), .B(new_n205_), .S(KEYINPUT82), .Z(new_n206_));
  XOR2_X1   g005(.A(new_n206_), .B(KEYINPUT31), .Z(new_n207_));
  AND2_X1   g006(.A1(new_n207_), .A2(KEYINPUT83), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(G169gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n212_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(G183gat), .B2(G190gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n210_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  NOR3_X1   g017(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n211_), .B(KEYINPUT23), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n223_), .A2(KEYINPUT81), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT25), .B(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT81), .B1(new_n226_), .B2(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n216_), .B1(new_n222_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(G15gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT30), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n230_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G71gat), .B(G99gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(G43gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n235_), .B(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n208_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n207_), .A2(KEYINPUT83), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n208_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G211gat), .B(G218gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G197gat), .B(G204gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT21), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT87), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n244_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n245_), .A2(new_n246_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n244_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n248_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n252_), .B1(new_n253_), .B2(new_n250_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G141gat), .A2(G148gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G155gat), .A2(G162gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(KEYINPUT1), .B2(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(KEYINPUT1), .ZN(new_n261_));
  AOI211_X1 g060(.A(new_n256_), .B(new_n257_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G155gat), .B(G162gat), .Z(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n264_), .A2(KEYINPUT84), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266_));
  AOI22_X1  g065(.A1(KEYINPUT2), .A2(new_n256_), .B1(new_n257_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(KEYINPUT84), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n263_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT86), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT86), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n275_), .B(new_n263_), .C1(new_n269_), .C2(new_n272_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n262_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n255_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G228gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G78gat), .B(G106gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n277_), .A2(new_n278_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G22gat), .B(G50gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT28), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n285_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n281_), .A2(new_n283_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n284_), .A2(new_n288_), .A3(KEYINPUT88), .A4(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT88), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n293_), .A2(new_n288_), .B1(new_n284_), .B2(new_n289_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n243_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT93), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n277_), .A2(new_n206_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n277_), .B2(new_n204_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G225gat), .A2(G233gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n299_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n277_), .A2(new_n204_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n303_), .B(KEYINPUT4), .C1(new_n277_), .C2(new_n206_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(G85gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G57gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT33), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n296_), .B1(new_n307_), .B2(new_n314_), .ZN(new_n315_));
  NOR4_X1   g114(.A1(new_n306_), .A2(KEYINPUT93), .A3(new_n313_), .A4(new_n312_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT19), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT90), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n223_), .A2(new_n225_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n220_), .A2(new_n221_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n216_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n321_), .B1(new_n255_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n255_), .A2(new_n230_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(KEYINPUT20), .A3(new_n326_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n255_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n320_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n255_), .A2(new_n230_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n251_), .A2(new_n254_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT89), .ZN(new_n334_));
  INV_X1    g133(.A(new_n324_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT89), .B1(new_n255_), .B2(new_n324_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n332_), .B(new_n319_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n329_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G8gat), .B(G36gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n344_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n329_), .A2(new_n338_), .A3(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(KEYINPUT92), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT92), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n339_), .A2(new_n349_), .A3(new_n344_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n299_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n351_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n304_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n311_), .B1(new_n298_), .B2(new_n351_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n348_), .A2(new_n350_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n300_), .A2(new_n305_), .A3(new_n311_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n313_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT94), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n357_), .A2(KEYINPUT94), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n317_), .A2(new_n355_), .A3(new_n358_), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n306_), .A2(new_n312_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n356_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n339_), .A2(KEYINPUT95), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n344_), .A2(KEYINPUT32), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT95), .B1(new_n329_), .B2(new_n338_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n332_), .B(new_n320_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n326_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n367_), .B1(new_n370_), .B2(new_n320_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n366_), .A2(new_n371_), .A3(new_n364_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n362_), .B1(new_n365_), .B2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n295_), .B1(new_n360_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n348_), .A2(new_n375_), .A3(new_n350_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n362_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n346_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n345_), .A3(KEYINPUT27), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n242_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n293_), .A2(new_n288_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n284_), .A2(new_n289_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n290_), .A3(new_n243_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n380_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n374_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G8gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT76), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G1gat), .ZN(new_n392_));
  INV_X1    g191(.A(G8gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT14), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT75), .B(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G22gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n391_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n394_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n390_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G29gat), .B(G36gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G43gat), .B(G50gat), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n402_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n405_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n408_));
  OAI211_X1 g207(.A(G229gat), .B(G233gat), .C1(new_n406_), .C2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n408_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G229gat), .A2(G233gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(KEYINPUT15), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT15), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n405_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n397_), .A2(new_n412_), .A3(new_n399_), .A4(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n410_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G113gat), .B(G141gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT79), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G169gat), .B(G197gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n409_), .A2(new_n416_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n409_), .B2(new_n416_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n388_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(KEYINPUT80), .A3(new_n421_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n387_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G231gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n400_), .B(new_n429_), .ZN(new_n430_));
  AND2_X1   g229(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(G78gat), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT66), .ZN(new_n434_));
  INV_X1    g233(.A(G71gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(G78gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(G57gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(G64gat), .ZN(new_n441_));
  INV_X1    g240(.A(G64gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(G57gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT11), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n441_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(G57gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n440_), .A2(G64gat), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT11), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n433_), .B(new_n439_), .C1(new_n445_), .C2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G57gat), .B(G64gat), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n433_), .A2(new_n439_), .B1(new_n450_), .B2(KEYINPUT11), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n430_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n430_), .A2(new_n453_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G127gat), .B(G155gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G183gat), .B(G211gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT17), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n456_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n461_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n454_), .A2(KEYINPUT17), .A3(new_n464_), .A4(new_n455_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT78), .Z(new_n467_));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468_));
  INV_X1    g267(.A(G85gat), .ZN(new_n469_));
  INV_X1    g268(.A(G92gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G85gat), .A2(G92gat), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT6), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(G99gat), .A3(G106gat), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT7), .ZN(new_n479_));
  INV_X1    g278(.A(G99gat), .ZN(new_n480_));
  INV_X1    g279(.A(G106gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n473_), .B1(new_n478_), .B2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT8), .B1(new_n473_), .B2(KEYINPUT65), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT8), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n471_), .A2(new_n472_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n491_), .B(new_n473_), .C1(new_n478_), .C2(new_n484_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n470_), .A2(KEYINPUT64), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT64), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G92gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n469_), .A2(KEYINPUT9), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n475_), .A2(new_n477_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n471_), .A2(KEYINPUT9), .A3(new_n472_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT10), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n480_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n481_), .A3(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .A4(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n487_), .A2(new_n492_), .A3(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n412_), .A2(new_n506_), .A3(new_n414_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT34), .Z(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n500_), .A2(new_n504_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n496_), .A2(new_n497_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n485_), .A2(new_n486_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(new_n405_), .A3(new_n492_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n507_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n509_), .A2(new_n510_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n517_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n507_), .A2(new_n519_), .A3(new_n511_), .A4(new_n515_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G190gat), .B(G218gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT72), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n525_), .A2(KEYINPUT36), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n521_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n525_), .B(KEYINPUT36), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(KEYINPUT73), .B2(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n529_), .A2(KEYINPUT73), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n468_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n518_), .A2(KEYINPUT74), .A3(new_n520_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT74), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n528_), .B1(new_n521_), .B2(new_n534_), .ZN(new_n535_));
  AOI211_X1 g334(.A(KEYINPUT37), .B(new_n527_), .C1(new_n533_), .C2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n467_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n506_), .A2(new_n453_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n444_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n431_), .A2(new_n432_), .A3(G78gat), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n437_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n451_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n514_), .B2(new_n492_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT12), .B1(new_n540_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT12), .B1(new_n506_), .B2(new_n453_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT68), .ZN(new_n554_));
  INV_X1    g353(.A(new_n483_), .ZN(new_n555_));
  NOR3_X1   g354(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n489_), .B1(new_n557_), .B2(new_n499_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n505_), .B1(new_n558_), .B2(new_n491_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n485_), .A2(new_n486_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n453_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n514_), .A2(new_n547_), .A3(new_n492_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n550_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT67), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n562_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n551_), .B1(new_n565_), .B2(KEYINPUT12), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT68), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n550_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n554_), .A2(new_n564_), .A3(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G120gat), .B(G148gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n554_), .A2(new_n564_), .A3(new_n568_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n575_), .B(new_n577_), .C1(KEYINPUT70), .C2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n539_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n428_), .A2(new_n585_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n586_), .A2(G1gat), .A3(new_n377_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT38), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(KEYINPUT38), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n527_), .B1(new_n535_), .B2(new_n533_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n387_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n427_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n583_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n466_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n377_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n589_), .A3(new_n596_), .ZN(G1324gat));
  INV_X1    g396(.A(new_n586_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n376_), .A2(new_n379_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n393_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G8gat), .B1(new_n595_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT97), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT97), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n605_), .B(G8gat), .C1(new_n595_), .C2(new_n601_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n604_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n600_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT40), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(KEYINPUT40), .B(new_n600_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1325gat));
  OAI21_X1  g412(.A(G15gat), .B1(new_n595_), .B2(new_n243_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT98), .B(KEYINPUT41), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n615_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n598_), .A2(new_n232_), .A3(new_n242_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .ZN(G1326gat));
  NAND2_X1  g418(.A1(new_n384_), .A2(new_n290_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G22gat), .B1(new_n595_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT42), .ZN(new_n622_));
  OR3_X1    g421(.A1(new_n586_), .A2(G22gat), .A3(new_n620_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT99), .Z(G1327gat));
  INV_X1    g424(.A(new_n467_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n428_), .A2(new_n583_), .A3(new_n626_), .A4(new_n590_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G29gat), .B1(new_n628_), .B2(new_n362_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n537_), .B1(new_n374_), .B2(new_n386_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT43), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n632_), .B(new_n537_), .C1(new_n374_), .C2(new_n386_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n467_), .A2(new_n593_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT44), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(KEYINPUT44), .A3(new_n635_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n634_), .A2(KEYINPUT100), .A3(KEYINPUT44), .A4(new_n635_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n362_), .A2(G29gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n629_), .B1(new_n641_), .B2(new_n642_), .ZN(G1328gat));
  INV_X1    g442(.A(KEYINPUT46), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT101), .ZN(new_n645_));
  INV_X1    g444(.A(G36gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n628_), .A2(new_n646_), .A3(new_n599_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT45), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n641_), .A2(new_n599_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n645_), .B(new_n648_), .C1(new_n649_), .C2(new_n646_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n646_), .B1(new_n641_), .B2(new_n599_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT45), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n647_), .B(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT101), .B(new_n644_), .C1(new_n651_), .C2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n650_), .A2(new_n654_), .ZN(G1329gat));
  XNOR2_X1  g454(.A(KEYINPUT102), .B(G43gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n628_), .B2(new_n242_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n242_), .A2(G43gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n641_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT47), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1330gat));
  INV_X1    g460(.A(new_n620_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G50gat), .B1(new_n628_), .B2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n662_), .A2(G50gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n641_), .B2(new_n664_), .ZN(G1331gat));
  NAND4_X1  g464(.A1(new_n591_), .A2(new_n427_), .A3(new_n584_), .A4(new_n467_), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT104), .B(G57gat), .Z(new_n667_));
  NOR3_X1   g466(.A1(new_n666_), .A2(new_n377_), .A3(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT105), .Z(new_n669_));
  NOR2_X1   g468(.A1(new_n387_), .A2(new_n592_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n539_), .A2(new_n583_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n673_), .A2(KEYINPUT103), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(KEYINPUT103), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n362_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n669_), .B1(new_n440_), .B2(new_n676_), .ZN(G1332gat));
  OAI21_X1  g476(.A(G64gat), .B1(new_n666_), .B2(new_n601_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT48), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n599_), .A2(new_n442_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT106), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n679_), .B1(new_n672_), .B2(new_n681_), .ZN(G1333gat));
  OAI21_X1  g481(.A(G71gat), .B1(new_n666_), .B2(new_n243_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT49), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n673_), .A2(new_n435_), .A3(new_n242_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1334gat));
  OAI21_X1  g485(.A(G78gat), .B1(new_n666_), .B2(new_n620_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT50), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n673_), .A2(new_n437_), .A3(new_n662_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT107), .ZN(G1335gat));
  INV_X1    g490(.A(new_n590_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n467_), .A2(new_n583_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n670_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G85gat), .B1(new_n695_), .B2(new_n362_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n467_), .A2(new_n592_), .A3(new_n583_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n362_), .A2(G85gat), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT108), .Z(new_n701_));
  AOI21_X1  g500(.A(new_n696_), .B1(new_n699_), .B2(new_n701_), .ZN(G1336gat));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n599_), .A3(new_n496_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n470_), .B1(new_n694_), .B2(new_n601_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1337gat));
  AND2_X1   g504(.A1(new_n699_), .A2(new_n242_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n242_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n707_));
  OAI22_X1  g506(.A1(new_n706_), .A2(new_n480_), .B1(new_n694_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n634_), .A2(KEYINPUT109), .A3(new_n662_), .A4(new_n697_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G106gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT109), .B1(new_n699_), .B2(new_n662_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n634_), .A2(new_n662_), .A3(new_n697_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n717_), .A2(KEYINPUT110), .A3(G106gat), .A4(new_n711_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n714_), .A2(KEYINPUT52), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n710_), .B(new_n720_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n695_), .A2(new_n481_), .A3(new_n662_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT53), .B1(new_n719_), .B2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n714_), .A2(KEYINPUT52), .A3(new_n718_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n721_), .A4(new_n722_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(G1339gat));
  INV_X1    g527(.A(KEYINPUT114), .ZN(new_n729_));
  INV_X1    g528(.A(new_n466_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n424_), .A2(new_n426_), .A3(new_n577_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n549_), .A2(KEYINPUT55), .A3(new_n550_), .A4(new_n552_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT111), .ZN(new_n733_));
  INV_X1    g532(.A(new_n566_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n550_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n566_), .A2(new_n737_), .A3(KEYINPUT55), .A4(new_n550_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(new_n736_), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n567_), .B1(new_n566_), .B2(new_n550_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT12), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n742_));
  NOR4_X1   g541(.A1(new_n742_), .A2(new_n551_), .A3(KEYINPUT68), .A4(new_n735_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n740_), .A2(new_n743_), .A3(KEYINPUT55), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT56), .B(new_n574_), .C1(new_n739_), .C2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n554_), .A2(new_n747_), .A3(new_n568_), .ZN(new_n748_));
  AOI22_X1  g547(.A1(new_n732_), .A2(KEYINPUT111), .B1(new_n734_), .B2(new_n735_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n738_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT56), .B1(new_n750_), .B2(new_n574_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n731_), .B1(new_n746_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n410_), .A2(new_n415_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n411_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n754_), .B2(new_n753_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n406_), .A2(new_n408_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n420_), .B1(new_n757_), .B2(new_n411_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n422_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n578_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n752_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT57), .B1(new_n761_), .B2(new_n692_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT57), .ZN(new_n763_));
  AOI211_X1 g562(.A(new_n763_), .B(new_n590_), .C1(new_n752_), .C2(new_n760_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n759_), .A2(new_n577_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n574_), .B1(new_n739_), .B2(new_n744_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n766_), .B1(new_n769_), .B2(new_n745_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n537_), .B1(new_n770_), .B2(KEYINPUT58), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(KEYINPUT58), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n537_), .B(KEYINPUT113), .C1(new_n770_), .C2(KEYINPUT58), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n730_), .B1(new_n765_), .B2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n467_), .A2(new_n427_), .A3(new_n583_), .A4(new_n538_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n729_), .B1(new_n777_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n775_), .A2(new_n774_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n759_), .A2(new_n577_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n746_), .B2(new_n751_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT58), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT113), .B1(new_n786_), .B2(new_n537_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n782_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n424_), .A2(new_n426_), .A3(new_n577_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n769_), .B2(new_n745_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n760_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n692_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n763_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n761_), .A2(KEYINPUT57), .A3(new_n692_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n466_), .B1(new_n788_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n778_), .B(KEYINPUT54), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(KEYINPUT114), .A3(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n381_), .A2(new_n377_), .A3(new_n599_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n781_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(G113gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n592_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(KEYINPUT59), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n799_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n626_), .B1(new_n788_), .B2(new_n795_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n797_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT115), .B1(new_n804_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n811_), .B(new_n808_), .C1(new_n800_), .C2(KEYINPUT59), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n810_), .A2(new_n812_), .A3(new_n427_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n803_), .B1(new_n813_), .B2(new_n802_), .ZN(G1340gat));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n583_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n801_), .B(new_n816_), .C1(KEYINPUT60), .C2(new_n815_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n817_), .A2(new_n818_), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n583_), .B(new_n808_), .C1(new_n800_), .C2(KEYINPUT59), .ZN(new_n821_));
  OAI22_X1  g620(.A1(new_n819_), .A2(new_n820_), .B1(new_n815_), .B2(new_n821_), .ZN(G1341gat));
  INV_X1    g621(.A(G127gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n800_), .B2(new_n626_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT117), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n810_), .A2(new_n812_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n466_), .A2(new_n823_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(G1342gat));
  INV_X1    g627(.A(G134gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n801_), .A2(new_n829_), .A3(new_n590_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n810_), .A2(new_n812_), .A3(new_n538_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n829_), .ZN(G1343gat));
  INV_X1    g631(.A(new_n385_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n599_), .A2(new_n377_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n781_), .A2(new_n798_), .A3(new_n833_), .A4(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n427_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT118), .B(G141gat), .Z(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1344gat));
  INV_X1    g637(.A(new_n835_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n584_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT120), .B1(new_n835_), .B2(new_n583_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT119), .B(G148gat), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n843_), .B(new_n845_), .ZN(G1345gat));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n839_), .A2(new_n847_), .A3(new_n467_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT121), .B1(new_n835_), .B2(new_n626_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT61), .B(G155gat), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n850_), .B(new_n852_), .ZN(G1346gat));
  OAI21_X1  g652(.A(G162gat), .B1(new_n835_), .B2(new_n538_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n692_), .A2(G162gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n835_), .B2(new_n855_), .ZN(G1347gat));
  NAND2_X1  g655(.A1(new_n807_), .A2(new_n797_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n601_), .A2(new_n381_), .A3(new_n362_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n592_), .A3(new_n858_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n859_), .A2(KEYINPUT122), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n861_));
  INV_X1    g660(.A(G169gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n859_), .B2(KEYINPUT122), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n860_), .A2(new_n861_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT22), .B(G169gat), .Z(new_n866_));
  OAI22_X1  g665(.A1(new_n864_), .A2(new_n865_), .B1(new_n859_), .B2(new_n866_), .ZN(G1348gat));
  AND2_X1   g666(.A1(new_n781_), .A2(new_n798_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n620_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n601_), .A2(new_n362_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n870_), .A2(G176gat), .A3(new_n242_), .A4(new_n584_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n857_), .A2(new_n858_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n583_), .ZN(new_n873_));
  OAI22_X1  g672(.A1(new_n869_), .A2(new_n871_), .B1(G176gat), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1349gat));
  NOR3_X1   g675(.A1(new_n872_), .A2(new_n225_), .A3(new_n466_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n870_), .A2(new_n242_), .A3(new_n467_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n869_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(G183gat), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n877_), .B1(new_n879_), .B2(new_n880_), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n857_), .A2(new_n537_), .A3(new_n858_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n882_), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT124), .B1(new_n882_), .B2(G190gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n590_), .A2(new_n223_), .ZN(new_n885_));
  OAI22_X1  g684(.A1(new_n883_), .A2(new_n884_), .B1(new_n872_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1351gat));
  NAND3_X1  g687(.A1(new_n868_), .A2(new_n833_), .A3(new_n870_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n427_), .ZN(new_n890_));
  INV_X1    g689(.A(G197gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1352gat));
  NOR2_X1   g691(.A1(new_n889_), .A2(new_n583_), .ZN(new_n893_));
  INV_X1    g692(.A(G204gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1353gat));
  AOI21_X1  g694(.A(new_n466_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT126), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n889_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1354gat));
  OAI21_X1  g699(.A(G218gat), .B1(new_n889_), .B2(new_n538_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n692_), .A2(G218gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n889_), .B2(new_n902_), .ZN(G1355gat));
endmodule


