//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT97), .ZN(new_n206_));
  XOR2_X1   g005(.A(G64gat), .B(G92gat), .Z(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT96), .ZN(new_n210_));
  INV_X1    g009(.A(G204gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT87), .B1(new_n211_), .B2(G197gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT87), .ZN(new_n213_));
  INV_X1    g012(.A(G197gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(G204gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(G197gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n212_), .A2(new_n215_), .A3(KEYINPUT88), .A4(new_n216_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT21), .ZN(new_n222_));
  INV_X1    g021(.A(G218gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G211gat), .ZN(new_n224_));
  INV_X1    g023(.A(G211gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G218gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n222_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n212_), .A2(new_n215_), .A3(new_n222_), .A4(new_n216_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n226_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n214_), .A2(G204gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n216_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(KEYINPUT21), .B2(new_n231_), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n221_), .A2(new_n227_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT79), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(G183gat), .B2(G190gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n236_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n234_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n235_), .A2(KEYINPUT77), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT23), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n239_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n238_), .A2(KEYINPUT23), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n241_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(KEYINPUT79), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT78), .ZN(new_n251_));
  INV_X1    g050(.A(G169gat), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n252_), .A2(KEYINPUT22), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(KEYINPUT22), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n251_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(KEYINPUT22), .ZN(new_n256_));
  AOI21_X1  g055(.A(G176gat), .B1(new_n256_), .B2(KEYINPUT78), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n255_), .A2(new_n257_), .B1(G169gat), .B2(G176gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n242_), .A2(new_n250_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G176gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(KEYINPUT24), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT25), .B(G183gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G190gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n237_), .A2(new_n238_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n239_), .A2(KEYINPUT23), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n261_), .A2(KEYINPUT24), .A3(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .A4(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n233_), .A2(new_n259_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT92), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT20), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n271_), .B2(KEYINPUT20), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n248_), .B(KEYINPUT95), .C1(new_n261_), .C2(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n264_), .A2(KEYINPUT93), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n264_), .A2(KEYINPUT93), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n263_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT95), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n275_), .A2(new_n261_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n280_), .B1(new_n240_), .B2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n275_), .A2(new_n261_), .A3(new_n268_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n276_), .A2(new_n279_), .A3(new_n282_), .A4(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n266_), .A2(new_n267_), .A3(new_n249_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n253_), .A2(new_n254_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n260_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n268_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n233_), .B1(new_n284_), .B2(new_n288_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n273_), .A2(new_n274_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT19), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n210_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n271_), .A2(KEYINPUT20), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT92), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT20), .ZN(new_n297_));
  INV_X1    g096(.A(new_n289_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(KEYINPUT96), .A3(new_n292_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n259_), .A2(new_n270_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n221_), .A2(new_n227_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n232_), .A2(new_n228_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n284_), .A2(new_n288_), .A3(new_n233_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT20), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(new_n292_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n209_), .B1(new_n301_), .B2(new_n310_), .ZN(new_n311_));
  AOI211_X1 g110(.A(new_n309_), .B(new_n208_), .C1(new_n294_), .C2(new_n300_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n203_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G127gat), .B(G134gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT31), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n302_), .B(KEYINPUT30), .ZN(new_n319_));
  XOR2_X1   g118(.A(G71gat), .B(G99gat), .Z(new_n320_));
  NAND2_X1  g119(.A1(G227gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G15gat), .B(G43gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT80), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n322_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n319_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n318_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OR3_X1    g127(.A1(new_n328_), .A2(new_n327_), .A3(new_n326_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT83), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT2), .ZN(new_n333_));
  INV_X1    g132(.A(G141gat), .ZN(new_n334_));
  INV_X1    g133(.A(G148gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT3), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT2), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n330_), .A2(new_n331_), .A3(new_n338_), .ZN(new_n339_));
  OR3_X1    g138(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n333_), .A2(new_n337_), .A3(new_n339_), .A4(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n342_), .A2(KEYINPUT1), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(G155gat), .B2(G162gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n342_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n336_), .A2(new_n330_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n350_), .A2(KEYINPUT82), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT82), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n348_), .A2(G155gat), .A3(G162gat), .ZN(new_n354_));
  INV_X1    g153(.A(G155gat), .ZN(new_n355_));
  INV_X1    g154(.A(G162gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT1), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n354_), .B1(new_n357_), .B2(new_n343_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n351_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n346_), .B1(new_n352_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n317_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT82), .B1(new_n350_), .B2(new_n351_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n358_), .A2(new_n353_), .A3(new_n359_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n317_), .A3(new_n346_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n363_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT98), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n317_), .B1(new_n366_), .B2(new_n346_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n364_), .A2(new_n365_), .B1(new_n341_), .B2(new_n345_), .ZN(new_n374_));
  NOR4_X1   g173(.A1(new_n374_), .A2(KEYINPUT98), .A3(KEYINPUT4), .A4(new_n317_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n363_), .A2(KEYINPUT4), .A3(new_n367_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n368_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n369_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT0), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G57gat), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n384_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n385_), .A2(new_n386_), .A3(G85gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(G85gat), .B1(new_n385_), .B2(new_n386_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n380_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n389_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n391_), .B(new_n369_), .C1(new_n376_), .C2(new_n379_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n328_), .B1(new_n327_), .B2(new_n326_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n329_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n301_), .A2(new_n310_), .A3(new_n209_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n308_), .A2(new_n293_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n299_), .B2(new_n293_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n400_), .B2(new_n208_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G78gat), .B(G106gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n404_), .B(KEYINPUT90), .Z(new_n405_));
  INV_X1    g204(.A(KEYINPUT89), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n233_), .B1(KEYINPUT29), .B2(new_n361_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(KEYINPUT86), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT29), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n305_), .B(new_n406_), .C1(new_n374_), .C2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  AOI211_X1 g212(.A(new_n406_), .B(new_n411_), .C1(new_n407_), .C2(KEYINPUT86), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n405_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT84), .B1(new_n361_), .B2(KEYINPUT29), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n374_), .A2(new_n418_), .A3(new_n409_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G22gat), .B(G50gat), .Z(new_n420_));
  AND3_X1   g219(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n416_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n417_), .A2(new_n419_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n420_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n416_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n423_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n305_), .B1(new_n374_), .B2(new_n409_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT89), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n408_), .A2(new_n412_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n404_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n415_), .A2(new_n430_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT91), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT91), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n415_), .A2(new_n430_), .A3(new_n439_), .A4(new_n436_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n413_), .A2(new_n414_), .A3(new_n405_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n405_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n429_), .B(new_n423_), .C1(new_n441_), .C2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n438_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n445_));
  NOR4_X1   g244(.A1(new_n314_), .A2(new_n396_), .A3(new_n403_), .A4(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n209_), .A2(KEYINPUT32), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n390_), .A2(new_n392_), .B1(new_n400_), .B2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n299_), .A2(KEYINPUT96), .A3(new_n292_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT96), .B1(new_n299_), .B2(new_n292_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n310_), .B(new_n447_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n311_), .A2(new_n312_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n392_), .A2(KEYINPUT99), .A3(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n363_), .A2(new_n367_), .A3(new_n378_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n389_), .A2(new_n457_), .A3(KEYINPUT100), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT100), .B1(new_n389_), .B2(new_n457_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n377_), .A2(new_n368_), .ZN(new_n460_));
  OAI22_X1  g259(.A1(new_n458_), .A2(new_n459_), .B1(new_n376_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n455_), .B1(new_n392_), .B2(KEYINPUT99), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n453_), .B1(new_n454_), .B2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT101), .B1(new_n465_), .B2(new_n445_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n313_), .A2(new_n394_), .A3(new_n445_), .A4(new_n402_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n310_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n208_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n464_), .A2(new_n469_), .A3(new_n397_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n449_), .A2(new_n452_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT101), .ZN(new_n473_));
  INV_X1    g272(.A(new_n445_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n466_), .A2(new_n467_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n329_), .A2(new_n395_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n446_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G190gat), .B(G218gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(G134gat), .B(G162gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(KEYINPUT36), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  AND2_X1   g283(.A1(G85gat), .A2(G92gat), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(KEYINPUT9), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT65), .B(G85gat), .Z(new_n487_));
  INV_X1    g286(.A(G92gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n486_), .B1(new_n489_), .B2(KEYINPUT9), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT6), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT10), .B(G99gat), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT64), .B(G106gat), .Z(new_n495_));
  OAI211_X1 g294(.A(new_n490_), .B(new_n492_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G85gat), .B(G92gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT66), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT7), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n492_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT68), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n492_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n492_), .A2(new_n506_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n501_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n499_), .B1(new_n509_), .B2(new_n498_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n496_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT70), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT70), .B(new_n496_), .C1(new_n505_), .C2(new_n510_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G29gat), .B(G36gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G43gat), .B(G50gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT15), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT72), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n496_), .B(new_n517_), .C1(new_n505_), .C2(new_n510_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .A4(new_n523_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n519_), .A2(new_n521_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT34), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n530_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n483_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n525_), .B(new_n526_), .C1(new_n528_), .C2(new_n530_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n481_), .B(KEYINPUT36), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n478_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G120gat), .B(G148gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT5), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G176gat), .B(G204gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G230gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G57gat), .B(G64gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n549_));
  XOR2_X1   g348(.A(G71gat), .B(G78gat), .Z(new_n550_));
  OR2_X1    g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n550_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n548_), .A2(KEYINPUT11), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n511_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n511_), .A2(new_n555_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n547_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT69), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(KEYINPUT69), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(KEYINPUT12), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n557_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n513_), .A2(KEYINPUT12), .A3(new_n514_), .A4(new_n555_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n564_), .A3(new_n547_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n546_), .B1(new_n561_), .B2(new_n565_), .ZN(new_n566_));
  AND4_X1   g365(.A1(new_n565_), .A2(new_n559_), .A3(new_n560_), .A4(new_n546_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT13), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n566_), .A2(KEYINPUT13), .A3(new_n567_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(G8gat), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(G22gat), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(G15gat), .ZN(new_n576_));
  INV_X1    g375(.A(G15gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(G22gat), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT73), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT73), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G1gat), .B(G8gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n582_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n518_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n517_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT74), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n585_), .B(new_n517_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(G229gat), .A3(G233gat), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n587_), .A2(KEYINPUT74), .A3(new_n588_), .A4(new_n589_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n592_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(G113gat), .B(G141gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT75), .ZN(new_n598_));
  XOR2_X1   g397(.A(G169gat), .B(G197gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT76), .ZN(new_n602_));
  INV_X1    g401(.A(new_n600_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n592_), .A2(new_n594_), .A3(new_n595_), .A4(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n596_), .A2(KEYINPUT76), .A3(new_n600_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n572_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n585_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(new_n554_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT17), .ZN(new_n613_));
  XOR2_X1   g412(.A(G127gat), .B(G155gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n612_), .A2(new_n613_), .A3(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(KEYINPUT17), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n612_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n541_), .A2(new_n608_), .A3(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT103), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n202_), .B1(new_n624_), .B2(new_n393_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT104), .ZN(new_n626_));
  INV_X1    g425(.A(new_n608_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n478_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n534_), .A2(KEYINPUT37), .A3(new_n538_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT37), .B1(new_n534_), .B2(new_n538_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(new_n621_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n628_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n202_), .A3(new_n393_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT38), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n626_), .A2(new_n637_), .ZN(G1324gat));
  NOR2_X1   g437(.A1(new_n314_), .A2(new_n403_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G8gat), .B1(new_n623_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT39), .ZN(new_n641_));
  INV_X1    g440(.A(new_n639_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n573_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g444(.A(new_n477_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n577_), .B1(new_n624_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n635_), .A2(new_n577_), .A3(new_n646_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(G1326gat));
  NAND2_X1  g451(.A1(new_n624_), .A2(new_n445_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G22gat), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n655_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n635_), .A2(new_n575_), .A3(new_n445_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(G1327gat));
  NOR2_X1   g458(.A1(new_n539_), .A2(new_n622_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n628_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G29gat), .B1(new_n661_), .B2(new_n393_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT106), .B(KEYINPUT43), .C1(new_n478_), .C2(new_n631_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n476_), .A2(new_n477_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n446_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n631_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n671_));
  NOR4_X1   g470(.A1(new_n478_), .A2(KEYINPUT107), .A3(KEYINPUT43), .A4(new_n631_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n663_), .B(new_n669_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n627_), .A2(new_n622_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(KEYINPUT44), .A3(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n675_), .A2(G29gat), .A3(new_n393_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n674_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n662_), .B1(new_n676_), .B2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n661_), .A2(new_n681_), .A3(new_n642_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n674_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n473_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n686_));
  AOI211_X1 g485(.A(KEYINPUT101), .B(new_n445_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n646_), .B1(new_n688_), .B2(new_n467_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n632_), .B1(new_n689_), .B2(new_n446_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT106), .B1(new_n690_), .B2(KEYINPUT43), .ZN(new_n691_));
  INV_X1    g490(.A(new_n663_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT107), .B1(new_n690_), .B2(KEYINPUT43), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n667_), .A2(new_n670_), .A3(new_n668_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n685_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n678_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n675_), .B(new_n642_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(G36gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(G36gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n684_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(KEYINPUT46), .B(new_n684_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  AND2_X1   g506(.A1(new_n646_), .A2(G43gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n679_), .A2(new_n675_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT111), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT111), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n679_), .A2(new_n711_), .A3(new_n675_), .A4(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G43gat), .B1(new_n661_), .B2(new_n646_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT112), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT47), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n713_), .A2(new_n715_), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1330gat));
  NAND3_X1  g519(.A1(new_n679_), .A2(new_n445_), .A3(new_n675_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G50gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n474_), .A2(G50gat), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT113), .Z(new_n724_));
  NAND2_X1  g523(.A1(new_n661_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1331gat));
  NAND4_X1  g525(.A1(new_n541_), .A2(new_n622_), .A3(new_n607_), .A4(new_n572_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n394_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n607_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n478_), .A2(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(KEYINPUT114), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(KEYINPUT114), .ZN(new_n732_));
  INV_X1    g531(.A(new_n572_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n633_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n393_), .A2(new_n384_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n728_), .B1(new_n735_), .B2(new_n736_), .ZN(G1332gat));
  OAI21_X1  g536(.A(G64gat), .B1(new_n727_), .B2(new_n639_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT48), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n639_), .A2(G64gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n735_), .B2(new_n740_), .ZN(G1333gat));
  OAI21_X1  g540(.A(G71gat), .B1(new_n727_), .B2(new_n477_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT49), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n477_), .A2(G71gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n735_), .B2(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n727_), .B2(new_n474_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT50), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n474_), .A2(G78gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n735_), .B2(new_n748_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT115), .Z(G1335gat));
  AND2_X1   g549(.A1(new_n734_), .A2(new_n660_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n393_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n733_), .A2(new_n622_), .A3(new_n729_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n673_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n394_), .A2(new_n487_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n752_), .B1(new_n754_), .B2(new_n755_), .ZN(G1336gat));
  AOI21_X1  g555(.A(G92gat), .B1(new_n751_), .B2(new_n642_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n642_), .A2(G92gat), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT116), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n757_), .B1(new_n754_), .B2(new_n759_), .ZN(G1337gat));
  NAND2_X1  g559(.A1(new_n754_), .A2(new_n646_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G99gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n751_), .A2(new_n493_), .A3(new_n646_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g564(.A1(new_n673_), .A2(new_n445_), .A3(new_n753_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G106gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT117), .B1(new_n767_), .B2(KEYINPUT52), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n766_), .A2(new_n769_), .A3(new_n770_), .A4(G106gat), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n767_), .A2(KEYINPUT52), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n768_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n474_), .A2(new_n495_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n751_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n773_), .A2(new_n778_), .A3(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n565_), .A2(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n563_), .A2(new_n564_), .A3(KEYINPUT55), .A4(new_n547_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n563_), .A2(new_n564_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n547_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n782_), .A2(new_n783_), .A3(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n545_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT119), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n787_), .A2(new_n790_), .A3(KEYINPUT56), .A4(new_n545_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n545_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n789_), .A2(new_n791_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n567_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n593_), .A2(new_n588_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n589_), .A2(new_n587_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n797_), .B(new_n600_), .C1(new_n588_), .C2(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n604_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n796_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT58), .B1(new_n795_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT120), .B1(new_n803_), .B2(new_n631_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n545_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(KEYINPUT119), .B2(new_n788_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n801_), .B1(new_n807_), .B2(new_n791_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n805_), .B(new_n632_), .C1(new_n808_), .C2(KEYINPUT58), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(KEYINPUT58), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n804_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n800_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n567_), .A2(new_n607_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n793_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n792_), .B2(new_n815_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n787_), .A2(new_n545_), .B1(new_n814_), .B2(new_n793_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n812_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT57), .B1(new_n818_), .B2(new_n539_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(KEYINPUT57), .A3(new_n539_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n818_), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n539_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n819_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n811_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n811_), .B2(new_n824_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n621_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n733_), .A2(new_n622_), .A3(new_n607_), .A4(new_n631_), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT54), .Z(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n642_), .A2(new_n445_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n393_), .A3(new_n646_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT59), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n811_), .A2(new_n824_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n621_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n831_), .A2(new_n839_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n835_), .A3(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n837_), .A2(new_n729_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G113gat), .ZN(new_n844_));
  OR3_X1    g643(.A1(new_n836_), .A2(G113gat), .A3(new_n607_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1340gat));
  NAND3_X1  g645(.A1(new_n837_), .A2(new_n572_), .A3(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G120gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n836_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n733_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n850_));
  AND2_X1   g649(.A1(KEYINPUT60), .A2(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n852_), .ZN(G1341gat));
  NAND3_X1  g652(.A1(new_n837_), .A2(new_n622_), .A3(new_n842_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G127gat), .ZN(new_n855_));
  OR3_X1    g654(.A1(new_n836_), .A2(G127gat), .A3(new_n621_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1342gat));
  AOI21_X1  g656(.A(G134gat), .B1(new_n849_), .B2(new_n540_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n837_), .A2(new_n842_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT124), .B(G134gat), .Z(new_n860_));
  NOR2_X1   g659(.A1(new_n631_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n858_), .B1(new_n859_), .B2(new_n861_), .ZN(G1343gat));
  NAND2_X1  g661(.A1(new_n838_), .A2(KEYINPUT122), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n811_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n830_), .B1(new_n865_), .B2(new_n621_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n642_), .A2(new_n474_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n868_), .A2(new_n394_), .A3(new_n646_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n866_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n729_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n572_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g674(.A1(new_n832_), .A2(new_n622_), .A3(new_n869_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT125), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n832_), .A2(new_n878_), .A3(new_n622_), .A4(new_n869_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT61), .B(G155gat), .Z(new_n880_));
  AND3_X1   g679(.A1(new_n877_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n877_), .B2(new_n879_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1346gat));
  NAND3_X1  g682(.A1(new_n871_), .A2(new_n356_), .A3(new_n540_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n866_), .A2(new_n631_), .A3(new_n870_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n356_), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n639_), .A2(new_n396_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n474_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n840_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G169gat), .B1(new_n890_), .B2(new_n607_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n892_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n890_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n286_), .A3(new_n729_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n894_), .A3(new_n896_), .ZN(G1348gat));
  NAND3_X1  g696(.A1(new_n840_), .A2(new_n572_), .A3(new_n889_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n572_), .A2(G176gat), .A3(new_n474_), .A4(new_n887_), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n899_), .A2(G176gat), .B1(new_n866_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  OAI221_X1 g702(.A(KEYINPUT126), .B1(new_n866_), .B2(new_n900_), .C1(new_n899_), .C2(G176gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1349gat));
  NAND2_X1  g704(.A1(new_n895_), .A2(new_n622_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n263_), .ZN(new_n907_));
  INV_X1    g706(.A(G183gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n906_), .ZN(G1350gat));
  NAND2_X1  g708(.A1(new_n895_), .A2(new_n632_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G190gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n540_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n890_), .B2(new_n912_), .ZN(G1351gat));
  NAND3_X1  g712(.A1(new_n477_), .A2(new_n445_), .A3(new_n394_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n866_), .A2(new_n639_), .A3(new_n914_), .ZN(new_n915_));
  AND3_X1   g714(.A1(new_n915_), .A2(G197gat), .A3(new_n729_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G197gat), .B1(new_n915_), .B2(new_n729_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1352gat));
  NAND2_X1  g717(.A1(new_n915_), .A2(new_n572_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G204gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n915_), .A2(new_n211_), .A3(new_n572_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1353gat));
  AOI21_X1  g721(.A(new_n621_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n915_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT127), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n924_), .A2(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n915_), .A2(new_n926_), .A3(new_n923_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1354gat));
  NAND3_X1  g729(.A1(new_n915_), .A2(new_n223_), .A3(new_n540_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n915_), .A2(new_n632_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n223_), .ZN(G1355gat));
endmodule


