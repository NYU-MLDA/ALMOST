//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_;
  INV_X1    g000(.A(G85gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  AND3_X1   g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n207_), .B1(new_n212_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT8), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n207_), .B(new_n221_), .C1(new_n212_), .C2(new_n218_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT64), .B1(new_n227_), .B2(new_n215_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229_));
  NOR4_X1   g028(.A1(new_n225_), .A2(new_n226_), .A3(new_n229_), .A4(G106gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n232_), .A2(new_n204_), .A3(new_n206_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n209_), .A2(new_n211_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n224_), .B1(new_n231_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n237_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT10), .B(G99gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n229_), .B1(new_n240_), .B2(G106gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n227_), .A2(KEYINPUT64), .A3(new_n215_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n243_), .A3(KEYINPUT66), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n223_), .A2(new_n238_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT68), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n223_), .A2(new_n238_), .A3(new_n247_), .A4(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G29gat), .B(G36gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G43gat), .B(G50gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n238_), .A2(KEYINPUT70), .A3(new_n244_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT70), .B1(new_n238_), .B2(new_n244_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n223_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n252_), .B(KEYINPUT15), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT73), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G232gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n260_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT35), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G190gat), .B(G218gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G134gat), .B(G162gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n259_), .A2(new_n266_), .B1(KEYINPUT36), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n269_), .A2(KEYINPUT36), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n264_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n273_));
  OR3_X1    g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT74), .B(KEYINPUT37), .Z(new_n280_));
  NOR2_X1   g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G15gat), .B(G22gat), .ZN(new_n284_));
  INV_X1    g083(.A(G1gat), .ZN(new_n285_));
  INV_X1    g084(.A(G8gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT14), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n284_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n287_), .A2(new_n288_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G1gat), .B(G8gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n291_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G231gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT69), .B(G71gat), .ZN(new_n297_));
  INV_X1    g096(.A(G78gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G57gat), .B(G64gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n300_), .A2(KEYINPUT11), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n300_), .A2(KEYINPUT11), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n299_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n296_), .B(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G127gat), .B(G155gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT77), .ZN(new_n309_));
  XOR2_X1   g108(.A(G183gat), .B(G211gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  AND2_X1   g112(.A1(new_n313_), .A2(KEYINPUT17), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n307_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n313_), .A2(KEYINPUT17), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n307_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n283_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT12), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n306_), .A2(new_n320_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n306_), .A2(new_n249_), .B1(new_n256_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n246_), .A2(new_n305_), .A3(new_n248_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n320_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n249_), .A2(new_n306_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n324_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n323_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G120gat), .B(G148gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT5), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G176gat), .B(G204gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT71), .ZN(new_n337_));
  INV_X1    g136(.A(new_n335_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n326_), .A2(new_n330_), .A3(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n331_), .A2(KEYINPUT71), .A3(new_n335_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT13), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT72), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT20), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n351_), .A2(KEYINPUT83), .B1(KEYINPUT23), .B2(new_n347_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(KEYINPUT83), .B2(new_n351_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT24), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G169gat), .ZN(new_n357_));
  INV_X1    g156(.A(G176gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT24), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n356_), .B1(new_n359_), .B2(new_n354_), .ZN(new_n360_));
  INV_X1    g159(.A(G190gat), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n361_), .A2(KEYINPUT81), .A3(KEYINPUT26), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n361_), .A2(KEYINPUT81), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(KEYINPUT26), .B2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT25), .B(G183gat), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n360_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT84), .B(G176gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G169gat), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n367_), .A2(new_n368_), .B1(G169gat), .B2(G176gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n349_), .B2(KEYINPUT23), .ZN(new_n371_));
  INV_X1    g170(.A(G183gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n361_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n353_), .A2(new_n366_), .B1(new_n369_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G197gat), .B(G204gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT21), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT90), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT89), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT89), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n381_), .A3(KEYINPUT90), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G211gat), .B(G218gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n376_), .A2(new_n377_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n386_), .B1(new_n378_), .B2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n376_), .A2(KEYINPUT88), .A3(new_n377_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n384_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n380_), .A2(new_n382_), .A3(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n385_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n346_), .B1(new_n375_), .B2(new_n393_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n383_), .A2(new_n384_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n369_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n353_), .B2(new_n373_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n354_), .B1(new_n359_), .B2(KEYINPUT94), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(KEYINPUT94), .B2(new_n359_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G190gat), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n365_), .A2(new_n400_), .B1(new_n355_), .B2(new_n354_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n371_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n395_), .B(new_n392_), .C1(new_n397_), .C2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n394_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G226gat), .A2(G233gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT19), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n397_), .A2(new_n403_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n409_), .B2(new_n393_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n393_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n353_), .A2(new_n366_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n374_), .A2(new_n369_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n346_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n410_), .A2(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G8gat), .B(G36gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n408_), .A2(new_n416_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT96), .ZN(new_n424_));
  INV_X1    g223(.A(new_n416_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n407_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n394_), .B2(new_n404_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n421_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT96), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n408_), .A2(new_n416_), .A3(new_n429_), .A4(new_n422_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n424_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT27), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n427_), .B1(new_n415_), .B2(new_n410_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n432_), .B1(new_n434_), .B2(new_n422_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT101), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT99), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n353_), .A2(new_n373_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n437_), .B(new_n402_), .C1(new_n438_), .C2(new_n396_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT99), .B1(new_n397_), .B2(new_n403_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n393_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n426_), .B1(new_n441_), .B2(new_n415_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n405_), .A2(new_n407_), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n436_), .B1(new_n444_), .B2(new_n421_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n436_), .B(new_n421_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n435_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G155gat), .A2(G162gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(G155gat), .B2(G162gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n451_), .B(KEYINPUT87), .C1(G155gat), .C2(G162gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(G141gat), .A2(G148gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT3), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G141gat), .A2(G148gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT2), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n451_), .A2(KEYINPUT1), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n451_), .B2(KEYINPUT1), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n457_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n459_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n462_), .A2(new_n463_), .A3(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G22gat), .B(G50gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT28), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n470_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G78gat), .B(G106gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n474_), .B(KEYINPUT91), .Z(new_n475_));
  NAND2_X1  g274(.A1(G228gat), .A2(G233gat), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n467_), .A2(new_n459_), .A3(new_n468_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n454_), .A2(new_n455_), .B1(new_n460_), .B2(new_n458_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT29), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n411_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n463_), .B1(new_n462_), .B2(new_n469_), .ZN(new_n481_));
  OAI211_X1 g280(.A(G228gat), .B(G233gat), .C1(new_n481_), .C2(new_n393_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n475_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n473_), .B1(new_n483_), .B2(KEYINPUT92), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT93), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n482_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n475_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n488_), .A2(new_n483_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n473_), .B(new_n490_), .C1(new_n483_), .C2(KEYINPUT92), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n485_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n489_), .B1(new_n485_), .B2(new_n491_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G227gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G15gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT30), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n375_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G127gat), .B(G134gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G120gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT85), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n498_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G71gat), .B(G99gat), .ZN(new_n504_));
  INV_X1    g303(.A(G43gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT31), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n507_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G1gat), .B(G29gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(G85gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT0), .B(G57gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G225gat), .A2(G233gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT97), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n462_), .A2(new_n469_), .A3(new_n501_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n502_), .B1(new_n462_), .B2(new_n469_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT4), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n462_), .A2(new_n469_), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n501_), .B(KEYINPUT85), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n517_), .B1(new_n521_), .B2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n524_), .A2(new_n518_), .A3(new_n515_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n514_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n525_), .B1(new_n524_), .B2(new_n518_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n520_), .A2(KEYINPUT4), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n516_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n514_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n528_), .A3(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n510_), .A2(new_n537_), .ZN(new_n538_));
  AND4_X1   g337(.A1(new_n433_), .A2(new_n448_), .A3(new_n494_), .A4(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n424_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n524_), .A2(new_n518_), .A3(new_n516_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n514_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT98), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n515_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT98), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n545_), .A3(new_n514_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n543_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n535_), .A2(KEYINPUT33), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT33), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n533_), .A2(new_n549_), .A3(new_n528_), .A4(new_n534_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(KEYINPUT32), .B(new_n422_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n422_), .A2(KEYINPUT32), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n530_), .A2(new_n535_), .B1(new_n434_), .B2(new_n553_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n540_), .A2(new_n551_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n485_), .A2(new_n491_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n489_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n485_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT100), .B1(new_n555_), .B2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n448_), .A2(new_n560_), .A3(new_n433_), .A4(new_n536_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n554_), .A2(new_n552_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n548_), .A2(new_n550_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n547_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n563_), .B1(new_n566_), .B2(new_n431_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT100), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n494_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n561_), .A2(new_n562_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n539_), .B1(new_n570_), .B2(new_n510_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT78), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n252_), .B(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(new_n294_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n257_), .A2(new_n294_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n573_), .B(new_n294_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n575_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n576_), .A2(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G113gat), .B(G141gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT79), .ZN(new_n582_));
  XOR2_X1   g381(.A(G169gat), .B(G197gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT80), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT80), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n580_), .A2(new_n584_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR4_X1   g390(.A1(new_n319_), .A2(new_n345_), .A3(new_n571_), .A4(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n285_), .A3(new_n537_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT38), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n318_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n344_), .A2(new_n590_), .ZN(new_n597_));
  NOR4_X1   g396(.A1(new_n571_), .A2(new_n596_), .A3(new_n277_), .A4(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n285_), .B1(new_n598_), .B2(new_n537_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n594_), .B2(new_n593_), .ZN(G1324gat));
  NAND2_X1  g400(.A1(new_n448_), .A2(new_n433_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n286_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT102), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n603_), .A2(new_n604_), .A3(KEYINPUT39), .ZN(new_n605_));
  INV_X1    g404(.A(new_n602_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(G8gat), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n605_), .B1(new_n592_), .B2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n603_), .A2(new_n604_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT39), .B1(new_n603_), .B2(new_n604_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n608_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g411(.A(G15gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n510_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n598_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n592_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n598_), .B2(new_n560_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT42), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n592_), .A2(new_n619_), .A3(new_n560_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1327gat));
  NOR2_X1   g422(.A1(new_n571_), .A2(new_n591_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n276_), .A2(new_n318_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n344_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G29gat), .B1(new_n628_), .B2(new_n537_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n571_), .A2(new_n283_), .A3(KEYINPUT43), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n570_), .A2(new_n510_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n539_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT103), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n571_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n282_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT104), .B1(new_n638_), .B2(KEYINPUT43), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n282_), .B1(new_n571_), .B2(new_n636_), .ZN(new_n640_));
  AOI211_X1 g439(.A(KEYINPUT103), .B(new_n539_), .C1(new_n570_), .C2(new_n510_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT104), .B(KEYINPUT43), .C1(new_n640_), .C2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n631_), .B1(new_n639_), .B2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n597_), .A2(new_n318_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n647_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(new_n645_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n537_), .A2(G29gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n629_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  NOR3_X1   g455(.A1(new_n627_), .A2(G36gat), .A3(new_n606_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT45), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n653_), .A2(new_n602_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n661_));
  INV_X1    g460(.A(G36gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT107), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n665_), .B(new_n659_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  NOR2_X1   g468(.A1(new_n510_), .A2(new_n505_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n650_), .A2(new_n653_), .A3(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n505_), .B1(new_n627_), .B2(new_n510_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT47), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT47), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n675_), .A3(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1330gat));
  AOI21_X1  g476(.A(G50gat), .B1(new_n628_), .B2(new_n560_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n560_), .A2(G50gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n654_), .B2(new_n679_), .ZN(G1331gat));
  NOR2_X1   g479(.A1(new_n590_), .A2(new_n596_), .ZN(new_n681_));
  AND4_X1   g480(.A1(new_n634_), .A2(new_n345_), .A3(new_n276_), .A4(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(G57gat), .A3(new_n537_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT108), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n319_), .A2(new_n344_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n571_), .A2(new_n590_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G57gat), .B1(new_n688_), .B2(new_n537_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n683_), .A2(KEYINPUT108), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n684_), .A2(new_n689_), .A3(new_n690_), .ZN(G1332gat));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n682_), .B2(new_n602_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT48), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n688_), .A2(new_n692_), .A3(new_n602_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1333gat));
  INV_X1    g495(.A(G71gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n682_), .B2(new_n614_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT49), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n688_), .A2(new_n697_), .A3(new_n614_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1334gat));
  AOI21_X1  g500(.A(new_n298_), .B1(new_n682_), .B2(new_n560_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT50), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n688_), .A2(new_n298_), .A3(new_n560_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1335gat));
  NOR3_X1   g504(.A1(new_n344_), .A2(new_n590_), .A3(new_n318_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n644_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G85gat), .B1(new_n707_), .B2(new_n536_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n345_), .A2(new_n625_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n686_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n202_), .A3(new_n537_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n712_), .ZN(G1336gat));
  OAI21_X1  g512(.A(G92gat), .B1(new_n707_), .B2(new_n606_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n203_), .A3(new_n602_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1337gat));
  NOR3_X1   g515(.A1(new_n710_), .A2(new_n510_), .A3(new_n240_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n644_), .A2(new_n614_), .A3(new_n706_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G99gat), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(G1338gat));
  NAND3_X1  g520(.A1(new_n711_), .A2(new_n215_), .A3(new_n560_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n640_), .B2(new_n641_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n630_), .B1(new_n725_), .B2(new_n642_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n706_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n726_), .A2(new_n494_), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT110), .B1(new_n728_), .B2(new_n215_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n730_), .B(G106gat), .C1(new_n707_), .C2(new_n494_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n729_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n722_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT53), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n722_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1339gat));
  INV_X1    g538(.A(KEYINPUT119), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n283_), .A2(new_n344_), .A3(new_n681_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT54), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n574_), .A2(new_n579_), .A3(new_n577_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n584_), .B1(new_n578_), .B2(new_n575_), .ZN(new_n744_));
  AOI22_X1  g543(.A1(new_n586_), .A2(new_n587_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(new_n339_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n256_), .A2(new_n321_), .ZN(new_n747_));
  AND4_X1   g546(.A1(new_n323_), .A2(new_n325_), .A3(new_n327_), .A4(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n325_), .A2(new_n327_), .A3(new_n747_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n329_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(KEYINPUT55), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n749_), .A2(new_n752_), .A3(new_n329_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n335_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n753_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n323_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n326_), .B1(new_n758_), .B2(new_n752_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(KEYINPUT56), .A4(new_n335_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n756_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n338_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n764_), .B2(KEYINPUT56), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n746_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT116), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT58), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n769_), .B(new_n746_), .C1(new_n763_), .C2(new_n765_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n768_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n282_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n766_), .A2(new_n768_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n771_), .A2(KEYINPUT117), .A3(new_n282_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT111), .B(KEYINPUT56), .Z(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT112), .B1(new_n764_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783_));
  INV_X1    g582(.A(new_n781_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n754_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n764_), .A2(KEYINPUT113), .A3(KEYINPUT56), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n780_), .A2(new_n782_), .A3(new_n785_), .A4(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n590_), .A2(new_n339_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n342_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n787_), .A2(new_n788_), .B1(new_n789_), .B2(new_n745_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n778_), .B1(new_n790_), .B2(new_n277_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n790_), .A2(new_n277_), .A3(new_n778_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(KEYINPUT114), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n790_), .A2(new_n277_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n778_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n777_), .A2(new_n793_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n318_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n777_), .A2(KEYINPUT118), .A3(new_n793_), .A4(new_n796_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n742_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n602_), .A2(new_n560_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(new_n537_), .A3(new_n614_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n740_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n776_), .A2(new_n775_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT117), .B1(new_n771_), .B2(new_n282_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n793_), .A2(new_n796_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n798_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(new_n596_), .A3(new_n800_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n742_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n803_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(KEYINPUT119), .A3(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n804_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(G113gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n590_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n794_), .A2(new_n778_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n807_), .A2(new_n818_), .A3(new_n792_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n811_), .B1(new_n819_), .B2(new_n318_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n813_), .A3(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n801_), .A2(new_n803_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(G113gat), .B1(new_n825_), .B2(new_n591_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n817_), .A2(new_n826_), .ZN(G1340gat));
  INV_X1    g626(.A(new_n345_), .ZN(new_n828_));
  OAI21_X1  g627(.A(G120gat), .B1(new_n825_), .B2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n344_), .A2(KEYINPUT60), .ZN(new_n830_));
  MUX2_X1   g629(.A(new_n830_), .B(KEYINPUT60), .S(G120gat), .Z(new_n831_));
  NAND2_X1  g630(.A1(new_n815_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n829_), .A2(new_n832_), .ZN(G1341gat));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n596_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n822_), .B(new_n835_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n804_), .A2(new_n318_), .A3(new_n814_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n834_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT121), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(new_n841_), .A3(new_n834_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n837_), .B1(new_n840_), .B2(new_n842_), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n815_), .A2(new_n844_), .A3(new_n277_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G134gat), .B1(new_n825_), .B2(new_n283_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1343gat));
  NOR4_X1   g646(.A1(new_n602_), .A2(new_n494_), .A3(new_n536_), .A4(new_n614_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n812_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n591_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT122), .B(G141gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1344gat));
  INV_X1    g651(.A(new_n849_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n345_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g654(.A1(new_n849_), .A2(new_n596_), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT61), .B(G155gat), .Z(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1346gat));
  OR3_X1    g657(.A1(new_n849_), .A2(G162gat), .A3(new_n276_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G162gat), .B1(new_n849_), .B2(new_n283_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1347gat));
  NAND2_X1  g660(.A1(new_n602_), .A2(new_n538_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n560_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n820_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n590_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n867_));
  INV_X1    g666(.A(new_n368_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n866_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT62), .B1(new_n866_), .B2(G169gat), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1348gat));
  OR2_X1    g670(.A1(new_n864_), .A2(new_n344_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n801_), .A2(new_n560_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n828_), .A2(new_n358_), .A3(new_n862_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n872_), .A2(new_n367_), .B1(new_n873_), .B2(new_n874_), .ZN(G1349gat));
  NOR3_X1   g674(.A1(new_n864_), .A2(new_n365_), .A3(new_n596_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT123), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n873_), .A2(new_n602_), .A3(new_n538_), .A4(new_n318_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n372_), .B2(new_n878_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n864_), .B2(new_n283_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n277_), .A2(new_n400_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n864_), .B2(new_n881_), .ZN(G1351gat));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n494_), .A2(new_n537_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(new_n602_), .A3(new_n510_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n886_));
  AOI211_X1 g685(.A(KEYINPUT125), .B(G197gat), .C1(new_n886_), .C2(new_n590_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888_));
  INV_X1    g687(.A(new_n885_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n812_), .A2(new_n590_), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(G197gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n888_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n887_), .A2(new_n892_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n812_), .A2(G197gat), .A3(new_n590_), .A4(new_n889_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT124), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n886_), .A2(new_n896_), .A3(G197gat), .A4(new_n590_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n883_), .B1(new_n893_), .B2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n897_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n900_), .B(KEYINPUT126), .C1(new_n892_), .C2(new_n887_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n886_), .A2(new_n345_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g703(.A(new_n886_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n596_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT63), .B(G211gat), .Z(new_n908_));
  AND3_X1   g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n906_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n907_), .B1(new_n906_), .B2(new_n908_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(G1354gat));
  OR3_X1    g711(.A1(new_n905_), .A2(G218gat), .A3(new_n276_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G218gat), .B1(new_n905_), .B2(new_n283_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1355gat));
endmodule


