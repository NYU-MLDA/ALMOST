//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT80), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G71gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G99gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT75), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT77), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT23), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n220_), .B(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n210_), .A2(KEYINPUT76), .A3(new_n213_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n216_), .A2(new_n224_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT22), .B(G169gat), .Z(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(G176gat), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n230_), .A2(KEYINPUT78), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT79), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n223_), .A2(new_n218_), .A3(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n217_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n233_), .B(new_n234_), .C1(G183gat), .C2(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(KEYINPUT78), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n231_), .A2(new_n207_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n205_), .A2(new_n228_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n205_), .B1(new_n228_), .B2(new_n237_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT82), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n240_), .B(new_n242_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n244_), .B1(new_n245_), .B2(KEYINPUT82), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  OR3_X1    g048(.A1(new_n238_), .A2(new_n239_), .A3(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G15gat), .B(G43gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT81), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT30), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT31), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n249_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n250_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G1gat), .B(G29gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(G85gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G57gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n271_));
  OAI22_X1  g070(.A1(new_n265_), .A2(new_n266_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n271_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT86), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n267_), .A2(new_n268_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n273_), .B(new_n276_), .C1(new_n275_), .C2(new_n274_), .ZN(new_n277_));
  AND2_X1   g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n265_), .B(KEYINPUT84), .Z(new_n282_));
  AOI22_X1  g081(.A1(new_n278_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n280_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n282_), .B(new_n283_), .C1(KEYINPUT1), .C2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n248_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n245_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(KEYINPUT4), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n248_), .A2(new_n291_), .A3(new_n286_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT96), .Z(new_n294_));
  NAND3_X1  g093(.A1(new_n290_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT97), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n290_), .A2(KEYINPUT97), .A3(new_n292_), .A4(new_n294_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n287_), .A2(new_n289_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n293_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n264_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n296_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n303_), .A2(new_n263_), .A3(new_n300_), .A4(new_n298_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n259_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT21), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G197gat), .B(G204gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT89), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310_));
  AOI211_X1 g109(.A(new_n307_), .B(new_n308_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n307_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n308_), .A2(KEYINPUT88), .ZN(new_n314_));
  INV_X1    g113(.A(G197gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G204gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT21), .B1(new_n316_), .B2(KEYINPUT88), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n313_), .B(new_n310_), .C1(new_n314_), .C2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G228gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT87), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n319_), .B(new_n321_), .C1(new_n288_), .C2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT90), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT90), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(new_n326_), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n325_), .A2(new_n327_), .B1(KEYINPUT29), .B2(new_n286_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n323_), .B1(new_n328_), .B2(new_n320_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n332_), .B(new_n323_), .C1(new_n328_), .C2(new_n320_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT91), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n286_), .A2(KEYINPUT29), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G22gat), .B(G50gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT28), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n338_), .B(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n335_), .A2(new_n342_), .ZN(new_n343_));
  OAI22_X1  g142(.A1(new_n331_), .A2(new_n334_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT27), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G226gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT19), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n224_), .B1(G183gat), .B2(G190gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n230_), .A3(new_n207_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n233_), .A2(new_n226_), .A3(new_n234_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT93), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n355_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n211_), .A2(new_n212_), .B1(new_n209_), .B2(new_n206_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT94), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT94), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n356_), .A2(new_n361_), .A3(new_n357_), .A4(new_n358_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n353_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT95), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(new_n324_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT20), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n237_), .A2(new_n228_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(new_n319_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n364_), .B1(new_n363_), .B2(new_n324_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n350_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n363_), .A2(new_n324_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT20), .B1(new_n367_), .B2(new_n319_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT92), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n374_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n372_), .A2(new_n375_), .A3(new_n349_), .A4(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n371_), .A2(new_n377_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n371_), .B2(new_n377_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n347_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n384_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n325_), .A2(new_n352_), .A3(new_n359_), .A4(new_n327_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n368_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n349_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n372_), .A2(new_n376_), .A3(new_n375_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n389_), .B1(new_n390_), .B2(new_n349_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n381_), .B(KEYINPUT98), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n347_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n386_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n306_), .A2(new_n346_), .A3(new_n385_), .A4(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT100), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n304_), .A2(KEYINPUT33), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n298_), .A2(new_n300_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n263_), .A4(new_n303_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n290_), .A2(new_n293_), .A3(new_n292_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n263_), .B1(new_n299_), .B2(new_n294_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n398_), .A2(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n383_), .A2(new_n384_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n302_), .A2(new_n304_), .B1(new_n408_), .B2(new_n391_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n371_), .A2(new_n377_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n345_), .B1(new_n406_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n394_), .A2(new_n385_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n305_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n345_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n259_), .B1(new_n413_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT99), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(KEYINPUT99), .B(new_n259_), .C1(new_n413_), .C2(new_n417_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n397_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G1gat), .B(G8gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT73), .ZN(new_n424_));
  OR2_X1    g223(.A1(G15gat), .A2(G22gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G15gat), .A2(G22gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G1gat), .A2(G8gat), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n425_), .A2(new_n426_), .B1(KEYINPUT14), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n424_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G43gat), .B(G50gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G29gat), .B(G36gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(KEYINPUT68), .ZN(new_n433_));
  INV_X1    g232(.A(G36gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(G29gat), .ZN(new_n435_));
  INV_X1    g234(.A(G29gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G36gat), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n435_), .A2(new_n437_), .A3(KEYINPUT68), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n431_), .B1(new_n433_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n437_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT68), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n432_), .A2(KEYINPUT68), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n430_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n429_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G229gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n429_), .A2(new_n445_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(new_n448_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n439_), .A2(KEYINPUT15), .A3(new_n444_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT15), .B1(new_n439_), .B2(new_n444_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n429_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n446_), .A2(new_n448_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G113gat), .B(G141gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(G169gat), .B(G197gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n454_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n422_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G99gat), .A2(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT6), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(G99gat), .A3(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n467_));
  INV_X1    g266(.A(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(G85gat), .ZN(new_n471_));
  INV_X1    g270(.A(G92gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G85gat), .A2(G92gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(KEYINPUT9), .A3(new_n474_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n474_), .A2(KEYINPUT9), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n466_), .A2(new_n470_), .A3(new_n475_), .A4(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n474_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI211_X1 g281(.A(KEYINPUT8), .B(new_n478_), .C1(new_n482_), .C2(new_n466_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT8), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  INV_X1    g284(.A(G99gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n468_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n464_), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n462_), .A2(KEYINPUT6), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n479_), .B(new_n487_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n478_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n484_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n477_), .B1(new_n483_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n477_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT8), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n490_), .A2(new_n484_), .A3(new_n491_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n445_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT70), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G232gat), .A2(G233gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n503_), .B(KEYINPUT34), .Z(new_n504_));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n494_), .A2(new_n501_), .A3(new_n502_), .A4(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n504_), .A2(new_n505_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n494_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n509_), .B(new_n510_), .C1(new_n508_), .C2(new_n511_), .ZN(new_n512_));
  OAI221_X1 g311(.A(new_n508_), .B1(new_n505_), .B2(new_n504_), .C1(new_n511_), .C2(KEYINPUT70), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G190gat), .B(G218gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G134gat), .B(G162gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT36), .Z(new_n517_));
  NAND3_X1  g316(.A1(new_n512_), .A2(new_n513_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT72), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n512_), .A2(new_n513_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n516_), .A2(KEYINPUT36), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT72), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n512_), .A2(new_n523_), .A3(new_n513_), .A4(new_n517_), .ZN(new_n524_));
  AND4_X1   g323(.A1(new_n461_), .A2(new_n519_), .A3(new_n522_), .A4(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT71), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n520_), .A2(KEYINPUT71), .A3(new_n521_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n518_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n525_), .B1(KEYINPUT37), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n429_), .B(new_n531_), .Z(new_n532_));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G71gat), .B(G78gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(KEYINPUT11), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n536_));
  INV_X1    g335(.A(new_n534_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n535_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(KEYINPUT74), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n532_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT17), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G127gat), .B(G155gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT16), .ZN(new_n546_));
  XOR2_X1   g345(.A(G183gat), .B(G211gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n543_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n544_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n542_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n530_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n540_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT64), .B1(new_n493_), .B2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n540_), .B(new_n477_), .C1(new_n483_), .C2(new_n492_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n493_), .A2(new_n557_), .A3(KEYINPUT64), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n556_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT65), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n493_), .A2(KEYINPUT12), .A3(new_n557_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n565_), .A2(new_n559_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT12), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n567_), .B1(new_n499_), .B2(new_n540_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT66), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT12), .B1(new_n493_), .B2(new_n557_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT66), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n566_), .A2(new_n569_), .A3(new_n572_), .A4(new_n555_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n563_), .A3(KEYINPUT65), .ZN(new_n574_));
  XOR2_X1   g373(.A(G120gat), .B(G148gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G176gat), .B(G204gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n564_), .A2(new_n574_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n564_), .B2(new_n574_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n582_), .A2(KEYINPUT13), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(KEYINPUT13), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n554_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n460_), .A2(new_n586_), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n587_), .A2(G1gat), .A3(new_n415_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n519_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT102), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n422_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n585_), .A2(new_n458_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n595_), .A2(new_n553_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G1gat), .B1(new_n597_), .B2(new_n415_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n590_), .A2(new_n591_), .A3(new_n598_), .ZN(G1324gat));
  INV_X1    g398(.A(KEYINPUT103), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n594_), .A2(new_n414_), .A3(new_n596_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n601_), .B2(G8gat), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n600_), .A3(G8gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n394_), .A2(new_n385_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n587_), .A2(G8gat), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n606_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n606_), .B2(new_n609_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1325gat));
  OAI21_X1  g412(.A(G15gat), .B1(new_n597_), .B2(new_n259_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT41), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n587_), .A2(G15gat), .A3(new_n259_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1326gat));
  OAI21_X1  g416(.A(G22gat), .B1(new_n597_), .B2(new_n346_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT42), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n346_), .A2(G22gat), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n619_), .B1(new_n587_), .B2(new_n620_), .ZN(G1327gat));
  NOR2_X1   g420(.A1(new_n552_), .A2(new_n592_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n585_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n460_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(G29gat), .B1(new_n625_), .B2(new_n305_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n595_), .A2(new_n552_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n530_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT43), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n422_), .A2(new_n628_), .A3(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n395_), .B(KEYINPUT100), .ZN(new_n635_));
  INV_X1    g434(.A(new_n421_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n404_), .A2(new_n405_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n637_));
  OAI22_X1  g436(.A1(new_n637_), .A2(new_n345_), .B1(new_n416_), .B2(new_n414_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT99), .B1(new_n638_), .B2(new_n259_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n636_), .B2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n634_), .B1(new_n640_), .B2(new_n530_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n627_), .B1(new_n632_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n640_), .B(new_n530_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n645_));
  OAI22_X1  g444(.A1(new_n422_), .A2(new_n628_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(KEYINPUT44), .A3(new_n627_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n415_), .A2(new_n436_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n626_), .B1(new_n649_), .B2(new_n650_), .ZN(G1328gat));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT46), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n644_), .A2(new_n414_), .A3(new_n648_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G36gat), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT45), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n414_), .B(KEYINPUT106), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(G36gat), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n460_), .A2(new_n658_), .A3(new_n623_), .A4(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n640_), .A2(new_n458_), .A3(new_n623_), .A4(new_n660_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT45), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n652_), .A2(new_n653_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n655_), .B1(new_n657_), .B2(new_n667_), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n654_), .B(new_n666_), .C1(new_n656_), .C2(G36gat), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1329gat));
  AND2_X1   g469(.A1(new_n258_), .A2(G43gat), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n644_), .A2(new_n648_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G43gat), .B1(new_n625_), .B2(new_n258_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n672_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n625_), .B2(new_n345_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n345_), .A2(G50gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n649_), .B2(new_n680_), .ZN(G1331gat));
  NOR3_X1   g480(.A1(new_n585_), .A2(new_n458_), .A3(new_n553_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n594_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G57gat), .B1(new_n683_), .B2(new_n415_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n585_), .A2(new_n458_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n640_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n554_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n415_), .A2(G57gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1332gat));
  OAI21_X1  g488(.A(G64gat), .B1(new_n683_), .B2(new_n659_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT48), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n659_), .A2(G64gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n687_), .B2(new_n692_), .ZN(G1333gat));
  OR3_X1    g492(.A1(new_n687_), .A2(G71gat), .A3(new_n259_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G71gat), .B1(new_n683_), .B2(new_n259_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n696_), .A2(new_n697_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n698_), .B2(new_n699_), .ZN(G1334gat));
  OAI21_X1  g499(.A(G78gat), .B1(new_n683_), .B2(new_n346_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT50), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n346_), .A2(G78gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n687_), .B2(new_n703_), .ZN(G1335gat));
  NAND2_X1  g503(.A1(new_n685_), .A2(new_n553_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G85gat), .B1(new_n707_), .B2(new_n415_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n686_), .A2(new_n622_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n471_), .A3(new_n305_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n708_), .A2(new_n711_), .ZN(G1336gat));
  OAI21_X1  g511(.A(G92gat), .B1(new_n707_), .B2(new_n659_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(new_n472_), .A3(new_n414_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1337gat));
  AOI21_X1  g514(.A(new_n486_), .B1(new_n706_), .B2(new_n258_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n258_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n709_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n716_), .A2(new_n718_), .B1(new_n719_), .B2(KEYINPUT51), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(KEYINPUT51), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1338gat));
  NAND3_X1  g521(.A1(new_n710_), .A2(new_n468_), .A3(new_n345_), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT52), .B(new_n468_), .C1(new_n706_), .C2(new_n345_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725_));
  INV_X1    g524(.A(new_n705_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n647_), .A2(new_n345_), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n727_), .B2(G106gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n723_), .B1(new_n724_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n723_), .B(new_n730_), .C1(new_n724_), .C2(new_n728_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1339gat));
  NAND2_X1  g533(.A1(new_n586_), .A2(new_n459_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n735_), .B(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n581_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n458_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n559_), .B(new_n565_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n568_), .A2(KEYINPUT66), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n556_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(KEYINPUT55), .A3(new_n573_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n741_), .A2(new_n742_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n555_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n744_), .A2(new_n745_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n745_), .B1(new_n744_), .B2(new_n748_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n579_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT56), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OAI211_X1 g552(.A(KEYINPUT56), .B(new_n579_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n740_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n457_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n453_), .B(new_n448_), .C1(new_n429_), .C2(new_n445_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n454_), .A2(new_n457_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT114), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n758_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n592_), .B1(new_n755_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(KEYINPUT57), .B(new_n592_), .C1(new_n755_), .C2(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n739_), .A2(new_n758_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n530_), .B1(new_n770_), .B2(KEYINPUT58), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(KEYINPUT115), .B(new_n530_), .C1(new_n770_), .C2(KEYINPUT58), .ZN(new_n774_));
  INV_X1    g573(.A(new_n769_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n744_), .A2(new_n748_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT113), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n744_), .A2(new_n745_), .A3(new_n748_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n579_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n754_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT58), .B(new_n775_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n770_), .A2(KEYINPUT116), .A3(KEYINPUT58), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n774_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n768_), .B1(new_n773_), .B2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n552_), .B1(new_n787_), .B2(KEYINPUT117), .ZN(new_n788_));
  INV_X1    g587(.A(new_n773_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n774_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n766_), .B(new_n767_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n738_), .B1(new_n788_), .B2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n607_), .A2(new_n305_), .A3(new_n346_), .A4(new_n258_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n787_), .A2(new_n552_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(new_n738_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n795_), .A2(new_n800_), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n796_), .A2(new_n797_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G113gat), .B1(new_n802_), .B2(new_n459_), .ZN(new_n803_));
  INV_X1    g602(.A(G113gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n796_), .A2(new_n804_), .A3(new_n458_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1340gat));
  OAI21_X1  g605(.A(G120gat), .B1(new_n802_), .B2(new_n585_), .ZN(new_n807_));
  INV_X1    g606(.A(G120gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n585_), .B2(KEYINPUT60), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n796_), .B(new_n809_), .C1(KEYINPUT60), .C2(new_n808_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(G1341gat));
  OAI21_X1  g610(.A(G127gat), .B1(new_n802_), .B2(new_n553_), .ZN(new_n812_));
  INV_X1    g611(.A(G127gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n796_), .A2(new_n813_), .A3(new_n552_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1342gat));
  OAI21_X1  g614(.A(G134gat), .B1(new_n802_), .B2(new_n628_), .ZN(new_n816_));
  INV_X1    g615(.A(G134gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n796_), .A2(new_n817_), .A3(new_n593_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1343gat));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n659_), .A2(new_n305_), .A3(new_n345_), .A4(new_n259_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT119), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n820_), .B1(new_n794_), .B2(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n735_), .B(new_n736_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n553_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n787_), .A2(KEYINPUT117), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(KEYINPUT120), .A3(new_n822_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n824_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n458_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g631(.A(new_n585_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g634(.A1(new_n830_), .A2(new_n552_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT61), .B(G155gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1346gat));
  AOI21_X1  g637(.A(G162gat), .B1(new_n830_), .B2(new_n593_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n530_), .A2(G162gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT121), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT122), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n830_), .A2(new_n841_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  INV_X1    g645(.A(new_n593_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n845_), .B(new_n846_), .C1(G162gat), .C2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n844_), .A2(new_n849_), .ZN(G1347gat));
  NOR3_X1   g649(.A1(new_n659_), .A2(new_n305_), .A3(new_n259_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n346_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n799_), .A2(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT124), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n459_), .A2(new_n229_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n458_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT123), .B1(new_n856_), .B2(G169gat), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n854_), .A2(new_n855_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n857_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n856_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(KEYINPUT62), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(G1348gat));
  NAND2_X1  g662(.A1(new_n828_), .A2(new_n346_), .ZN(new_n864_));
  INV_X1    g663(.A(G176gat), .ZN(new_n865_));
  INV_X1    g664(.A(new_n851_), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n585_), .A4(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n854_), .A2(new_n833_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n865_), .ZN(G1349gat));
  NOR3_X1   g668(.A1(new_n864_), .A2(new_n553_), .A3(new_n866_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(G183gat), .B1(new_n870_), .B2(new_n871_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n553_), .A2(new_n211_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n872_), .A2(new_n873_), .B1(new_n854_), .B2(new_n874_), .ZN(G1350gat));
  NAND3_X1  g674(.A1(new_n854_), .A2(new_n212_), .A3(new_n593_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n854_), .A2(new_n530_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n222_), .ZN(G1351gat));
  NOR3_X1   g677(.A1(new_n659_), .A2(new_n416_), .A3(new_n258_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n828_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n459_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n315_), .ZN(G1352gat));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n585_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1353gat));
  INV_X1    g684(.A(new_n880_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n553_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT127), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n888_), .B(new_n890_), .ZN(G1354gat));
  OR3_X1    g690(.A1(new_n880_), .A2(G218gat), .A3(new_n847_), .ZN(new_n892_));
  OAI21_X1  g691(.A(G218gat), .B1(new_n880_), .B2(new_n628_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1355gat));
endmodule


