//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OR3_X1    g003(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT23), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n204_), .A2(new_n205_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT82), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT22), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT83), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT84), .B(G176gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n215_), .B1(KEYINPUT83), .B2(KEYINPUT22), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n207_), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n210_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n214_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT21), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n226_), .A2(new_n227_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT20), .B1(new_n225_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G226gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT19), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n209_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n208_), .B1(new_n240_), .B2(new_n211_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT22), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G169gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n216_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT92), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(new_n219_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n222_), .A2(new_n210_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n241_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n239_), .B1(new_n234_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n225_), .A2(new_n235_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT93), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n248_), .A2(new_n251_), .A3(new_n234_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n251_), .B1(new_n248_), .B2(new_n234_), .ZN(new_n253_));
  OAI211_X1 g052(.A(KEYINPUT20), .B(new_n250_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n254_), .A2(KEYINPUT94), .A3(new_n238_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT94), .B1(new_n254_), .B2(new_n238_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n249_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G64gat), .B(G92gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n264_), .B(new_n249_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT27), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT89), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n234_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n232_), .A2(KEYINPUT89), .A3(new_n233_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n248_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n238_), .B1(new_n270_), .B2(new_n236_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT98), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI211_X1 g072(.A(KEYINPUT98), .B(new_n238_), .C1(new_n270_), .C2(new_n236_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n273_), .B(new_n274_), .C1(new_n238_), .C2(new_n254_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n262_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n265_), .A2(new_n276_), .A3(KEYINPUT27), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n266_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT85), .B(KEYINPUT86), .Z(new_n280_));
  NAND2_X1  g079(.A1(G227gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G71gat), .B(G99gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G15gat), .B(G43gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n224_), .B(KEYINPUT30), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT87), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n286_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT31), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n288_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G127gat), .B(G134gat), .ZN(new_n292_));
  INV_X1    g091(.A(G113gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(G120gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n291_), .B(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n290_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n290_), .A2(new_n296_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n301_), .B(new_n302_), .C1(new_n305_), .C2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n303_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n302_), .B(KEYINPUT1), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n310_), .B(new_n306_), .C1(new_n311_), .C2(new_n300_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n295_), .A2(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n294_), .A2(G120gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n294_), .A2(G120gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n315_), .A2(new_n312_), .A3(new_n309_), .A4(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n317_), .A3(KEYINPUT4), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G225gat), .A2(G233gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n318_), .B(new_n320_), .C1(KEYINPUT4), .C2(new_n314_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n314_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(KEYINPUT96), .B(KEYINPUT0), .Z(new_n324_));
  XNOR2_X1  g123(.A(G1gat), .B(G29gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G57gat), .B(G85gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n321_), .A2(new_n330_), .A3(new_n322_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n299_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n313_), .A2(KEYINPUT29), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G228gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT88), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n234_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n268_), .A2(new_n335_), .A3(new_n269_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n337_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n339_), .A2(KEYINPUT90), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT90), .B1(new_n339_), .B2(new_n340_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n338_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G78gat), .B(G106gat), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n343_), .A2(new_n345_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT91), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n313_), .A2(KEYINPUT29), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n351_), .B(KEYINPUT28), .Z(new_n352_));
  XOR2_X1   g151(.A(G22gat), .B(G50gat), .Z(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  OAI22_X1  g153(.A1(new_n347_), .A2(new_n348_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n343_), .A2(new_n345_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n352_), .B(new_n353_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n356_), .A2(new_n349_), .A3(new_n346_), .A4(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n279_), .A2(new_n334_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT99), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n358_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n266_), .A2(new_n362_), .A3(new_n277_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n332_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n275_), .A2(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n366_), .B(new_n332_), .C1(new_n257_), .C2(new_n365_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT33), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n331_), .A2(new_n368_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n318_), .B(new_n319_), .C1(KEYINPUT4), .C2(new_n314_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n314_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n328_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT97), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n321_), .A2(KEYINPUT33), .A3(new_n330_), .A4(new_n322_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n369_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n263_), .A2(new_n265_), .A3(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n372_), .A2(KEYINPUT97), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n367_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n363_), .A2(new_n364_), .B1(new_n378_), .B2(new_n362_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n299_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n361_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n362_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n263_), .A2(new_n265_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n265_), .A2(new_n276_), .A3(KEYINPUT27), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n385_), .A2(new_n359_), .A3(new_n364_), .A4(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(KEYINPUT99), .A3(new_n299_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n360_), .B1(new_n381_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G232gat), .A2(G233gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n391_), .B(KEYINPUT69), .Z(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT34), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT35), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT66), .ZN(new_n400_));
  AND3_X1   g199(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n400_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G99gat), .A2(G106gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(KEYINPUT66), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n399_), .A2(new_n403_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G85gat), .A2(G92gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(G85gat), .A2(G92gat), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n411_), .A2(new_n412_), .A3(KEYINPUT8), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT7), .ZN(new_n415_));
  INV_X1    g214(.A(G99gat), .ZN(new_n416_));
  INV_X1    g215(.A(G106gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n418_), .A2(new_n406_), .A3(new_n407_), .A4(new_n396_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n411_), .A2(new_n412_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT8), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n414_), .A2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(G29gat), .A2(G36gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G29gat), .A2(G36gat), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n424_), .A2(new_n425_), .A3(KEYINPUT70), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT70), .ZN(new_n427_));
  INV_X1    g226(.A(G29gat), .ZN(new_n428_));
  INV_X1    g227(.A(G36gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G29gat), .A2(G36gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(G43gat), .B1(new_n426_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT70), .B1(new_n424_), .B2(new_n425_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n435_));
  INV_X1    g234(.A(G43gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n433_), .A2(G50gat), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G50gat), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n436_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT10), .B(G99gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT64), .B1(new_n443_), .B2(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT64), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n416_), .A2(KEYINPUT10), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n416_), .A2(KEYINPUT10), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n445_), .B(new_n417_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n403_), .A2(new_n408_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT9), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n410_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n412_), .B1(new_n452_), .B2(KEYINPUT65), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n411_), .A2(KEYINPUT9), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT65), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n410_), .A2(new_n455_), .A3(new_n451_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n449_), .A2(new_n450_), .A3(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n423_), .A2(new_n438_), .A3(new_n442_), .A4(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n393_), .A2(new_n394_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT71), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n442_), .A2(new_n438_), .A3(KEYINPUT15), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT15), .B1(new_n442_), .B2(new_n438_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n458_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT68), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n423_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n414_), .A2(new_n422_), .A3(KEYINPUT68), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n467_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n462_), .B1(new_n466_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT15), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n440_), .A2(new_n441_), .A3(new_n439_), .ZN(new_n474_));
  AOI21_X1  g273(.A(G50gat), .B1(new_n433_), .B2(new_n437_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n463_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n414_), .A2(KEYINPUT68), .A3(new_n422_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT68), .B1(new_n414_), .B2(new_n422_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n458_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(new_n480_), .A3(KEYINPUT71), .ZN(new_n481_));
  AOI211_X1 g280(.A(new_n395_), .B(new_n461_), .C1(new_n472_), .C2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n395_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n472_), .A2(new_n481_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT72), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n461_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n459_), .A2(KEYINPUT72), .A3(new_n460_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI211_X1 g288(.A(KEYINPUT73), .B(new_n484_), .C1(new_n485_), .C2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT73), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n477_), .A2(new_n480_), .A3(KEYINPUT71), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT71), .B1(new_n477_), .B2(new_n480_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n487_), .B(new_n488_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n491_), .B1(new_n494_), .B2(new_n395_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n483_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G190gat), .B(G218gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT74), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(G134gat), .ZN(new_n499_));
  INV_X1    g298(.A(G162gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT75), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n496_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n496_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n501_), .B(KEYINPUT36), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n506_), .B(KEYINPUT37), .C1(new_n507_), .C2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n496_), .A2(KEYINPUT76), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n487_), .A2(new_n488_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n472_), .B2(new_n481_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT73), .B1(new_n514_), .B2(new_n484_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n494_), .A2(new_n491_), .A3(new_n395_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT76), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n483_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n512_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT77), .B1(new_n520_), .B2(new_n508_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT77), .ZN(new_n522_));
  AOI211_X1 g321(.A(new_n522_), .B(new_n509_), .C1(new_n512_), .C2(new_n519_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n506_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT37), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n511_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT78), .B(G15gat), .ZN(new_n527_));
  INV_X1    g326(.A(G22gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(G1gat), .ZN(new_n530_));
  INV_X1    g329(.A(G8gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT14), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G1gat), .B(G8gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT79), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n533_), .B(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G57gat), .B(G64gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT11), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT67), .ZN(new_n541_));
  INV_X1    g340(.A(G71gat), .ZN(new_n542_));
  INV_X1    g341(.A(G78gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n544_), .B(new_n545_), .C1(new_n539_), .C2(KEYINPUT11), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n541_), .A2(new_n546_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n538_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G127gat), .B(G155gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT16), .ZN(new_n554_));
  XOR2_X1   g353(.A(G183gat), .B(G211gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n552_), .B(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n550_), .A2(KEYINPUT17), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n526_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n423_), .A2(new_n458_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n549_), .B2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n541_), .B(new_n546_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n480_), .A2(KEYINPUT12), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n549_), .A2(new_n563_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n564_), .A2(new_n566_), .A3(new_n567_), .A4(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n565_), .B(new_n563_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n570_), .B2(new_n567_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G176gat), .ZN(new_n574_));
  INV_X1    g373(.A(G204gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n576_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT13), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(KEYINPUT13), .A3(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n442_), .A2(new_n438_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n536_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n536_), .B2(new_n477_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT81), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n536_), .B(new_n584_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(G229gat), .A3(G233gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(new_n215_), .ZN(new_n595_));
  INV_X1    g394(.A(G197gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n597_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n583_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n390_), .A2(new_n561_), .A3(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n530_), .A3(new_n332_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT38), .ZN(new_n606_));
  INV_X1    g405(.A(new_n360_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT99), .B1(new_n388_), .B2(new_n299_), .ZN(new_n608_));
  AOI211_X1 g407(.A(new_n361_), .B(new_n380_), .C1(new_n382_), .C2(new_n387_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n607_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n560_), .A2(new_n602_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT100), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n524_), .A2(KEYINPUT101), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n518_), .B1(new_n517_), .B2(new_n483_), .ZN(new_n614_));
  AOI211_X1 g413(.A(KEYINPUT76), .B(new_n482_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n508_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n522_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n520_), .A2(KEYINPUT77), .A3(new_n508_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(new_n506_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n613_), .A2(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n611_), .A2(KEYINPUT100), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n610_), .A2(new_n612_), .A3(new_n622_), .A4(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G1gat), .B1(new_n624_), .B2(new_n364_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n606_), .A2(new_n625_), .ZN(G1324gat));
  OAI21_X1  g425(.A(G8gat), .B1(new_n624_), .B2(new_n278_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT39), .B1(new_n627_), .B2(KEYINPUT102), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(KEYINPUT102), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n604_), .A2(new_n531_), .A3(new_n279_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n630_), .A2(KEYINPUT40), .A3(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n624_), .B2(new_n299_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT41), .Z(new_n638_));
  INV_X1    g437(.A(G15gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n604_), .A2(new_n639_), .A3(new_n380_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(G1326gat));
  NAND3_X1  g440(.A1(new_n604_), .A2(new_n528_), .A3(new_n359_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G22gat), .B1(new_n624_), .B2(new_n362_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT103), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n643_), .A2(KEYINPUT103), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n643_), .A2(KEYINPUT103), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT42), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n642_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT104), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n652_), .B(new_n642_), .C1(new_n646_), .C2(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1327gat));
  OAI21_X1  g453(.A(KEYINPUT43), .B1(new_n390_), .B2(new_n526_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  INV_X1    g455(.A(new_n526_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n610_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n603_), .A2(new_n560_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(KEYINPUT44), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  INV_X1    g463(.A(new_n660_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n666_), .B2(KEYINPUT105), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n428_), .B1(new_n668_), .B2(new_n332_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n390_), .A2(new_n622_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n660_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n671_), .A2(G29gat), .A3(new_n364_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n669_), .A2(KEYINPUT106), .A3(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT106), .B1(new_n669_), .B2(new_n672_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1328gat));
  AOI21_X1  g474(.A(new_n429_), .B1(new_n668_), .B2(new_n279_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n671_), .A2(G36gat), .A3(new_n278_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n677_), .B(new_n678_), .Z(new_n679_));
  NOR2_X1   g478(.A1(new_n676_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT46), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n676_), .B2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1329gat));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n663_), .A2(new_n667_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G43gat), .B1(new_n686_), .B2(new_n299_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n670_), .A2(new_n436_), .A3(new_n380_), .A4(new_n660_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n685_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n299_), .B1(new_n663_), .B2(new_n667_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n685_), .B(new_n688_), .C1(new_n690_), .C2(new_n436_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n689_), .A2(new_n692_), .ZN(G1330gat));
  OAI21_X1  g492(.A(G50gat), .B1(new_n686_), .B2(new_n362_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n359_), .A2(new_n439_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n671_), .B2(new_n695_), .ZN(G1331gat));
  NAND2_X1  g495(.A1(new_n560_), .A2(new_n601_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n610_), .A2(new_n583_), .A3(new_n622_), .A4(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(G57gat), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n364_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n583_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n561_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(KEYINPUT108), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(KEYINPUT108), .ZN(new_n705_));
  NOR4_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n600_), .A4(new_n390_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n332_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n701_), .B1(new_n707_), .B2(new_n700_), .ZN(G1332gat));
  INV_X1    g507(.A(G64gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n706_), .A2(new_n709_), .A3(new_n279_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G64gat), .B1(new_n699_), .B2(new_n278_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT48), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1333gat));
  NAND3_X1  g512(.A1(new_n706_), .A2(new_n542_), .A3(new_n380_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G71gat), .B1(new_n699_), .B2(new_n299_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1334gat));
  OAI21_X1  g516(.A(G78gat), .B1(new_n699_), .B2(new_n362_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT109), .Z(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n706_), .A2(new_n543_), .A3(new_n359_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1335gat));
  NOR3_X1   g521(.A1(new_n560_), .A2(new_n600_), .A3(new_n702_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n670_), .A2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT110), .ZN(new_n725_));
  AOI21_X1  g524(.A(G85gat), .B1(new_n725_), .B2(new_n332_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n659_), .A2(new_n723_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT111), .Z(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(new_n364_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n729_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g529(.A(G92gat), .B1(new_n725_), .B2(new_n279_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n728_), .A2(new_n278_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(G92gat), .ZN(G1337gat));
  OAI211_X1 g532(.A(new_n725_), .B(new_n380_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G99gat), .B1(new_n727_), .B2(new_n299_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738_));
  INV_X1    g537(.A(new_n723_), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n362_), .B(new_n739_), .C1(new_n655_), .C2(new_n658_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n740_), .B2(new_n417_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT112), .B(G106gat), .C1(new_n727_), .C2(new_n362_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(KEYINPUT52), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n725_), .A2(new_n417_), .A3(new_n359_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n738_), .B(new_n745_), .C1(new_n740_), .C2(new_n417_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n743_), .A2(new_n744_), .A3(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g547(.A(new_n505_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n702_), .B(new_n510_), .C1(new_n749_), .C2(KEYINPUT37), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n751_), .A2(new_n698_), .A3(new_n752_), .A4(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n753_), .B(new_n754_), .C1(new_n750_), .C2(new_n697_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n569_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT55), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n564_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(G230gat), .A3(G233gat), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n569_), .A2(new_n759_), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n763_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n576_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(KEYINPUT56), .A3(new_n576_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(KEYINPUT115), .A3(new_n770_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n770_), .A2(KEYINPUT115), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n600_), .A4(new_n577_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n586_), .A2(KEYINPUT116), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n586_), .A2(KEYINPUT116), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n588_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n591_), .A2(new_n589_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n597_), .A3(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n778_), .A2(KEYINPUT117), .A3(new_n598_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT117), .B1(new_n778_), .B2(new_n598_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n579_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n773_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n613_), .B2(new_n621_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT57), .B1(new_n784_), .B2(KEYINPUT118), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n620_), .B1(new_n619_), .B2(new_n506_), .ZN(new_n786_));
  AOI211_X1 g585(.A(KEYINPUT101), .B(new_n505_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n782_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n769_), .A2(new_n770_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n577_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n793_), .B(new_n794_), .Z(new_n795_));
  NAND2_X1  g594(.A1(new_n657_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n785_), .A2(new_n791_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n758_), .B1(new_n797_), .B2(new_n559_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n279_), .A2(new_n364_), .A3(new_n299_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n798_), .A2(new_n359_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(G113gat), .B1(new_n801_), .B2(new_n600_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n797_), .A2(new_n559_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n758_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n362_), .A3(new_n799_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n359_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n799_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n601_), .A2(new_n293_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n802_), .B1(new_n812_), .B2(new_n813_), .ZN(G1340gat));
  INV_X1    g613(.A(KEYINPUT60), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n702_), .B2(G120gat), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n801_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n807_), .A2(new_n817_), .A3(new_n583_), .A4(new_n810_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G120gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n801_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1341gat));
  AOI21_X1  g620(.A(G127gat), .B1(new_n801_), .B2(new_n560_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n560_), .A2(G127gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n812_), .B2(new_n823_), .ZN(G1342gat));
  AOI21_X1  g623(.A(new_n809_), .B1(new_n808_), .B2(new_n799_), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n798_), .A2(KEYINPUT59), .A3(new_n359_), .A4(new_n800_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n657_), .A2(G134gat), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n622_), .ZN(new_n829_));
  AOI21_X1  g628(.A(G134gat), .B1(new_n801_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT120), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832_));
  INV_X1    g631(.A(G134gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n806_), .B2(new_n622_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n832_), .B(new_n834_), .C1(new_n811_), .C2(new_n827_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n835_), .ZN(G1343gat));
  NOR2_X1   g635(.A1(new_n380_), .A2(new_n364_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n805_), .A2(new_n363_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n600_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n583_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g641(.A(KEYINPUT61), .B(G155gat), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n838_), .A2(new_n560_), .A3(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n805_), .A2(new_n363_), .A3(new_n837_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n843_), .B1(new_n846_), .B2(new_n559_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT121), .B(KEYINPUT122), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n845_), .A2(new_n847_), .A3(new_n849_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1346gat));
  AOI21_X1  g652(.A(G162gat), .B1(new_n838_), .B2(new_n829_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n846_), .A2(new_n500_), .A3(new_n526_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1347gat));
  NAND3_X1  g655(.A1(new_n808_), .A2(new_n333_), .A3(new_n279_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n857_), .A2(new_n601_), .A3(new_n245_), .ZN(new_n858_));
  NOR4_X1   g657(.A1(new_n798_), .A2(new_n334_), .A3(new_n359_), .A4(new_n278_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n215_), .B1(new_n859_), .B2(new_n600_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT62), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n860_), .A2(KEYINPUT62), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1348gat));
  NOR2_X1   g662(.A1(new_n857_), .A2(new_n702_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n219_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(G176gat), .B2(new_n864_), .ZN(G1349gat));
  NAND2_X1  g665(.A1(new_n859_), .A2(new_n560_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(KEYINPUT123), .B2(G183gat), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n202_), .B1(new_n869_), .B2(G183gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n867_), .B2(new_n870_), .ZN(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n857_), .B2(new_n526_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n859_), .A2(new_n829_), .A3(new_n203_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1351gat));
  NOR2_X1   g673(.A1(new_n798_), .A2(new_n278_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n359_), .A2(new_n364_), .A3(new_n299_), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(KEYINPUT124), .Z(new_n877_));
  AND3_X1   g676(.A1(new_n875_), .A2(new_n600_), .A3(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT125), .B1(new_n878_), .B2(G197gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(G197gat), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n875_), .A2(new_n877_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n881_), .B(new_n596_), .C1(new_n882_), .C2(new_n601_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n879_), .A2(new_n880_), .A3(new_n883_), .ZN(G1352gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n702_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n575_), .ZN(G1353gat));
  NAND3_X1  g685(.A1(new_n875_), .A2(new_n560_), .A3(new_n877_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  AND2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n887_), .B2(new_n888_), .ZN(G1354gat));
  OAI21_X1  g690(.A(KEYINPUT126), .B1(new_n882_), .B2(new_n622_), .ZN(new_n892_));
  INV_X1    g691(.A(G218gat), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n875_), .A2(new_n894_), .A3(new_n829_), .A4(new_n877_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(new_n893_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n657_), .A2(G218gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT127), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n875_), .A2(new_n877_), .A3(new_n898_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n896_), .A2(new_n899_), .ZN(G1355gat));
endmodule


