//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT71), .ZN(new_n205_));
  INV_X1    g004(.A(G36gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G29gat), .ZN(new_n207_));
  INV_X1    g006(.A(G29gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G36gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n207_), .A2(new_n209_), .A3(KEYINPUT71), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n205_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(new_n209_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n204_), .A2(KEYINPUT71), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(new_n202_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(KEYINPUT6), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT6), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(KEYINPUT65), .ZN(new_n230_));
  OAI22_X1  g029(.A1(new_n228_), .A2(new_n230_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(KEYINPUT65), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(KEYINPUT6), .ZN(new_n233_));
  AND2_X1   g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n226_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G85gat), .ZN(new_n237_));
  INV_X1    g036(.A(G92gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G85gat), .A2(G92gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n220_), .B1(new_n236_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n225_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT66), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n224_), .A2(new_n246_), .A3(new_n225_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n234_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n245_), .B(new_n247_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n241_), .A2(new_n220_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n223_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n239_), .A2(KEYINPUT9), .A3(new_n240_), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n240_), .A2(KEYINPUT9), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n231_), .A2(new_n235_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n242_), .A2(new_n252_), .A3(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G232gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT69), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n219_), .A2(new_n261_), .B1(new_n262_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n261_), .A2(KEYINPUT67), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n242_), .A2(new_n252_), .A3(new_n260_), .A4(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n217_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n266_), .A2(new_n262_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G190gat), .B(G218gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G134gat), .B(G162gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(KEYINPUT36), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n267_), .B(new_n272_), .C1(new_n262_), .C2(new_n266_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n275_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n278_), .B(KEYINPUT36), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n275_), .A2(new_n280_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n284_), .B1(new_n285_), .B2(KEYINPUT72), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n275_), .A2(new_n287_), .A3(new_n280_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n282_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G225gat), .A2(G233gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT3), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT2), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT86), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(KEYINPUT1), .B2(new_n297_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(KEYINPUT1), .B2(new_n297_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n291_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(new_n293_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G113gat), .B(G120gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n300_), .A2(new_n310_), .A3(new_n304_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(KEYINPUT4), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT4), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n305_), .A2(new_n313_), .A3(new_n308_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n290_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G1gat), .B(G29gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G57gat), .B(G85gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  INV_X1    g119(.A(new_n290_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n322_));
  OR3_X1    g121(.A1(new_n315_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n320_), .B1(new_n315_), .B2(new_n322_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G197gat), .A2(G204gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT87), .B(G204gat), .Z(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n330_), .B2(G197gat), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n331_), .A2(KEYINPUT21), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G211gat), .B(G218gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n330_), .A2(G197gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT21), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(G197gat), .B2(G204gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n333_), .A2(new_n336_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n332_), .A2(new_n338_), .B1(new_n331_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT25), .B(G183gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G190gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT23), .ZN(new_n348_));
  OR3_X1    g147(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n348_), .A2(KEYINPUT92), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(KEYINPUT92), .B1(new_n348_), .B2(new_n349_), .ZN(new_n351_));
  OAI221_X1 g150(.A(new_n344_), .B1(new_n345_), .B2(new_n346_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(new_n347_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(new_n354_), .B2(new_n347_), .ZN(new_n356_));
  OAI21_X1  g155(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n357_));
  OR3_X1    g156(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n328_), .B1(new_n341_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n348_), .A2(new_n349_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT79), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n342_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n367_), .B2(G183gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n343_), .A2(new_n368_), .ZN(new_n369_));
  OAI22_X1  g168(.A1(new_n366_), .A2(new_n369_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n363_), .B1(new_n364_), .B2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n370_), .A2(new_n364_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n340_), .B(new_n359_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n361_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n359_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n341_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n360_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n328_), .B1(new_n382_), .B2(new_n340_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n383_), .A3(new_n377_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n384_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n390_), .B1(new_n379_), .B2(new_n384_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n327_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OR3_X1    g193(.A1(new_n374_), .A2(KEYINPUT98), .A3(new_n378_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n381_), .A2(new_n383_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT98), .B1(new_n396_), .B2(new_n378_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n374_), .A2(new_n378_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n395_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT99), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n391_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n379_), .A2(new_n384_), .A3(new_n390_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(KEYINPUT27), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n400_), .B1(new_n399_), .B2(new_n391_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n326_), .B(new_n394_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n380_), .A2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G71gat), .B(G99gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT81), .ZN(new_n410_));
  INV_X1    g209(.A(G15gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT80), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT82), .ZN(new_n414_));
  AND2_X1   g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n412_), .B(new_n416_), .ZN(new_n417_));
  OAI211_X1 g216(.A(KEYINPUT30), .B(new_n359_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n408_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n419_), .A2(KEYINPUT84), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(KEYINPUT84), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n408_), .A2(new_n418_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n417_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n422_), .A2(KEYINPUT83), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT83), .B1(new_n422_), .B2(new_n423_), .ZN(new_n425_));
  OAI22_X1  g224(.A1(new_n420_), .A2(new_n421_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT85), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n419_), .B(KEYINPUT84), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n428_), .B(new_n429_), .C1(new_n425_), .C2(new_n424_), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n308_), .B(KEYINPUT31), .Z(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n340_), .B1(new_n305_), .B2(KEYINPUT29), .ZN(new_n435_));
  INV_X1    g234(.A(G228gat), .ZN(new_n436_));
  INV_X1    g235(.A(G233gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n438_), .B1(new_n442_), .B2(new_n340_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT90), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n434_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT28), .B1(new_n305_), .B2(KEYINPUT29), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT28), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n300_), .A2(new_n448_), .A3(new_n441_), .A4(new_n304_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G22gat), .B(G50gat), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n447_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n440_), .A2(KEYINPUT90), .A3(new_n443_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n446_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n433_), .B(KEYINPUT88), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR4_X1   g257(.A1(new_n453_), .A2(new_n456_), .A3(new_n444_), .A4(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n444_), .A2(new_n458_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n447_), .A2(new_n449_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n450_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n447_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n456_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n444_), .A2(new_n458_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n460_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n455_), .B1(new_n459_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n431_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n426_), .A2(KEYINPUT85), .A3(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n432_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n468_), .B1(new_n470_), .B2(new_n432_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n406_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n385_), .B2(KEYINPUT97), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT97), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT32), .B(new_n390_), .C1(new_n385_), .C2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n477_), .B2(new_n399_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n325_), .ZN(new_n479_));
  OAI211_X1 g278(.A(KEYINPUT33), .B(new_n320_), .C1(new_n315_), .C2(new_n322_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT95), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT33), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n324_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n392_), .A2(new_n393_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n309_), .A2(new_n321_), .A3(new_n311_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n320_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT96), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n312_), .A2(new_n290_), .A3(new_n314_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(KEYINPUT96), .A3(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n484_), .B(new_n485_), .C1(new_n488_), .C2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n479_), .B1(new_n482_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n432_), .A2(new_n470_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n468_), .A3(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n289_), .B1(new_n473_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G127gat), .B(G155gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT16), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G183gat), .B(G211gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT75), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G231gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n507_));
  XOR2_X1   g306(.A(G71gat), .B(G78gat), .Z(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n507_), .A2(new_n508_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n505_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n504_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n503_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n513_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G1gat), .B(G8gat), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT74), .ZN(new_n522_));
  NOR2_X1   g321(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(KEYINPUT73), .A2(G15gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(G22gat), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(G22gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n525_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(new_n528_), .B2(new_n523_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT14), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(G1gat), .B2(G8gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n522_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  AOI211_X1 g333(.A(KEYINPUT74), .B(new_n532_), .C1(new_n526_), .C2(new_n529_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n521_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(G22gat), .B1(new_n524_), .B2(new_n525_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n528_), .A2(new_n523_), .A3(new_n527_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n533_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT74), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n530_), .A2(new_n522_), .A3(new_n533_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(new_n520_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n519_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n515_), .A2(new_n518_), .A3(new_n542_), .A4(new_n536_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n501_), .A2(new_n502_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n536_), .A2(new_n542_), .A3(new_n217_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n217_), .B1(new_n536_), .B2(new_n542_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n543_), .A2(new_n271_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n217_), .A2(new_n218_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT15), .B1(new_n211_), .B2(new_n216_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n536_), .B(new_n542_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n548_), .B(KEYINPUT76), .Z(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n551_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G113gat), .B(G141gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G169gat), .B(G197gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n551_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT64), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n268_), .A2(new_n270_), .A3(new_n513_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n513_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n568_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n514_), .A2(new_n261_), .A3(KEYINPUT12), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(new_n570_), .B2(KEYINPUT12), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n268_), .A2(new_n270_), .A3(new_n513_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n567_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n571_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT5), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n580_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n571_), .B(new_n582_), .C1(new_n573_), .C2(new_n575_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n581_), .A2(KEYINPUT13), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT13), .B1(new_n581_), .B2(new_n583_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n496_), .A2(new_n547_), .A3(new_n565_), .A4(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(G1gat), .B1(new_n587_), .B2(new_n326_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT101), .Z(new_n589_));
  INV_X1    g388(.A(new_n565_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n473_), .B2(new_n495_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n285_), .A2(new_n283_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(KEYINPUT37), .A3(new_n281_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n289_), .B2(KEYINPUT37), .ZN(new_n594_));
  INV_X1    g393(.A(new_n547_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n591_), .A2(new_n586_), .A3(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n597_), .A2(G1gat), .A3(new_n326_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT38), .Z(new_n599_));
  NAND2_X1  g398(.A1(new_n589_), .A2(new_n599_), .ZN(G1324gat));
  OR2_X1    g399(.A1(new_n403_), .A2(new_n404_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n601_), .A2(new_n394_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G8gat), .B1(new_n587_), .B2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT39), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n597_), .A2(G8gat), .A3(new_n602_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT40), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(G1325gat));
  OAI21_X1  g407(.A(G15gat), .B1(new_n587_), .B2(new_n494_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT41), .Z(new_n610_));
  INV_X1    g409(.A(new_n494_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n411_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n597_), .B2(new_n612_), .ZN(G1326gat));
  OAI21_X1  g412(.A(G22gat), .B1(new_n587_), .B2(new_n468_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT42), .ZN(new_n615_));
  INV_X1    g414(.A(new_n468_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n527_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT102), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n615_), .B1(new_n597_), .B2(new_n618_), .ZN(G1327gat));
  NAND2_X1  g418(.A1(new_n595_), .A2(new_n289_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n586_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n494_), .A2(new_n616_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n432_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n405_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n493_), .A2(new_n468_), .A3(new_n494_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n565_), .B(new_n622_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT104), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n591_), .A2(new_n629_), .A3(new_n622_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(G29gat), .B1(new_n631_), .B2(new_n325_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n595_), .A2(new_n586_), .A3(new_n565_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT103), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n473_), .A2(new_n495_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n637_), .B2(new_n594_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n593_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n285_), .A2(KEYINPUT72), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n288_), .A3(new_n283_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n281_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT37), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  AOI211_X1 g443(.A(KEYINPUT43), .B(new_n644_), .C1(new_n473_), .C2(new_n495_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n635_), .B1(new_n638_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n594_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT43), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n637_), .A2(new_n636_), .A3(new_n594_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(KEYINPUT44), .A3(new_n635_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n648_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n326_), .A2(new_n208_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n632_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  INV_X1    g455(.A(new_n602_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n648_), .A2(new_n657_), .A3(new_n653_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(G36gat), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n602_), .A2(G36gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n628_), .A2(new_n630_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT105), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n628_), .A2(new_n630_), .A3(new_n664_), .A4(new_n660_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n662_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n663_), .B1(new_n662_), .B2(new_n665_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n659_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(KEYINPUT46), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  OAI221_X1 g470(.A(new_n659_), .B1(new_n669_), .B2(KEYINPUT46), .C1(new_n667_), .C2(new_n666_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1329gat));
  INV_X1    g472(.A(G43gat), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n494_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n648_), .A2(new_n653_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n648_), .A2(new_n653_), .A3(KEYINPUT107), .A4(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n631_), .A2(new_n611_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n674_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT47), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n678_), .A2(new_n684_), .A3(new_n679_), .A4(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1330gat));
  INV_X1    g485(.A(G50gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n631_), .A2(new_n687_), .A3(new_n616_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n654_), .A2(KEYINPUT108), .A3(new_n616_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT108), .B1(new_n654_), .B2(new_n616_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(G1331gat));
  NOR3_X1   g491(.A1(new_n595_), .A2(new_n586_), .A3(new_n565_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n496_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n326_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n565_), .B1(new_n473_), .B2(new_n495_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n621_), .A3(new_n596_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n326_), .A2(G57gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n695_), .B1(new_n697_), .B2(new_n698_), .ZN(G1332gat));
  NAND3_X1  g498(.A1(new_n496_), .A2(new_n657_), .A3(new_n693_), .ZN(new_n700_));
  XOR2_X1   g499(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(G64gat), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n700_), .B2(G64gat), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n602_), .A2(G64gat), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT110), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n703_), .A2(new_n704_), .B1(new_n697_), .B2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT111), .Z(G1333gat));
  OAI21_X1  g507(.A(G71gat), .B1(new_n694_), .B2(new_n494_), .ZN(new_n709_));
  XOR2_X1   g508(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n494_), .A2(G71gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n697_), .B2(new_n712_), .ZN(G1334gat));
  OAI21_X1  g512(.A(G78gat), .B1(new_n694_), .B2(new_n468_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT50), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n468_), .A2(G78gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n697_), .B2(new_n716_), .ZN(G1335gat));
  NAND3_X1  g516(.A1(new_n621_), .A2(new_n595_), .A3(new_n590_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n652_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n326_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n620_), .A2(new_n586_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n696_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n237_), .A3(new_n325_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n721_), .A2(new_n725_), .ZN(G1336gat));
  OAI21_X1  g525(.A(G92gat), .B1(new_n720_), .B2(new_n602_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n724_), .A2(new_n238_), .A3(new_n657_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1337gat));
  NAND3_X1  g528(.A1(new_n611_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n723_), .A2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT113), .Z(new_n732_));
  OAI21_X1  g531(.A(G99gat), .B1(new_n720_), .B2(new_n494_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(G1338gat));
  INV_X1    g535(.A(KEYINPUT115), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n468_), .B(new_n718_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(new_n223_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n652_), .A2(new_n616_), .A3(new_n719_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n739_), .A2(KEYINPUT52), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n737_), .B(new_n743_), .C1(new_n738_), .C2(new_n223_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n724_), .A2(new_n223_), .A3(new_n616_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT53), .B1(new_n742_), .B2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n739_), .A2(KEYINPUT52), .A3(new_n741_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n744_), .A4(new_n745_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(G1339gat));
  NAND4_X1  g550(.A1(new_n644_), .A2(new_n586_), .A3(new_n547_), .A4(new_n590_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n596_), .A2(new_n590_), .A3(new_n586_), .A4(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT119), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n574_), .A2(new_n567_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n243_), .A2(new_n244_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n241_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n765_), .A2(new_n220_), .B1(new_n259_), .B2(new_n258_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n269_), .B1(new_n766_), .B2(new_n252_), .ZN(new_n767_));
  AND4_X1   g566(.A1(new_n269_), .A2(new_n242_), .A3(new_n252_), .A4(new_n260_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n514_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT12), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n761_), .A2(new_n771_), .A3(KEYINPUT55), .A4(new_n572_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n574_), .B(new_n572_), .C1(new_n570_), .C2(KEYINPUT12), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n568_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n760_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n580_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n580_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  INV_X1    g579(.A(new_n583_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n556_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n556_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n552_), .A2(new_n555_), .A3(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n784_), .A3(new_n562_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT117), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n782_), .A2(new_n784_), .A3(new_n787_), .A4(new_n562_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n564_), .A3(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n780_), .B1(new_n781_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n564_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n550_), .A2(new_n556_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n561_), .B1(new_n792_), .B2(new_n555_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n787_), .B1(new_n793_), .B2(new_n782_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n791_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(KEYINPUT118), .A3(new_n583_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n778_), .A2(new_n779_), .B1(new_n790_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n594_), .B1(new_n797_), .B2(KEYINPUT58), .ZN(new_n798_));
  INV_X1    g597(.A(new_n779_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n580_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n791_), .ZN(new_n801_));
  AND4_X1   g600(.A1(KEYINPUT118), .A2(new_n801_), .A3(new_n583_), .A4(new_n786_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT118), .B1(new_n795_), .B2(new_n583_), .ZN(new_n803_));
  OAI22_X1  g602(.A1(new_n799_), .A2(new_n800_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n758_), .B1(new_n798_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n805_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n797_), .A2(KEYINPUT58), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(KEYINPUT119), .A4(new_n594_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n565_), .A2(new_n583_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n789_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n642_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT57), .B(new_n642_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n807_), .A2(new_n810_), .A3(new_n816_), .A4(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n757_), .B1(new_n818_), .B2(new_n595_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n602_), .A2(new_n325_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n471_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n819_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G113gat), .B1(new_n823_), .B2(new_n565_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT59), .B1(new_n819_), .B2(new_n822_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n819_), .C2(new_n822_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n816_), .B(new_n817_), .C1(new_n806_), .C2(new_n798_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n757_), .B1(new_n595_), .B2(new_n830_), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n820_), .A2(KEYINPUT59), .A3(new_n624_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT121), .B1(new_n829_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n836_), .B(new_n833_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n565_), .A2(G113gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n824_), .B1(new_n838_), .B2(new_n839_), .ZN(G1340gat));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n586_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n823_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n586_), .B(new_n833_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n841_), .ZN(G1341gat));
  AOI21_X1  g644(.A(G127gat), .B1(new_n823_), .B2(new_n547_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n547_), .A2(G127gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n838_), .B2(new_n847_), .ZN(G1342gat));
  AOI21_X1  g647(.A(G134gat), .B1(new_n823_), .B2(new_n289_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n594_), .A2(G134gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n838_), .B2(new_n850_), .ZN(G1343gat));
  NOR2_X1   g650(.A1(new_n819_), .A2(new_n623_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n821_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n565_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n621_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g657(.A1(new_n853_), .A2(new_n595_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT61), .B(G155gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1346gat));
  OR3_X1    g660(.A1(new_n853_), .A2(G162gat), .A3(new_n642_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G162gat), .B1(new_n853_), .B2(new_n644_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n602_), .A2(new_n325_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n611_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n590_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT122), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n468_), .ZN(new_n869_));
  OAI21_X1  g668(.A(G169gat), .B1(new_n869_), .B2(new_n831_), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n865_), .A2(new_n471_), .ZN(new_n873_));
  OR3_X1    g672(.A1(new_n831_), .A2(KEYINPUT124), .A3(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT124), .B1(new_n831_), .B2(new_n873_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT22), .B(G169gat), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n874_), .A2(new_n565_), .A3(new_n875_), .A4(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n872_), .B(new_n877_), .C1(new_n870_), .C2(new_n878_), .ZN(G1348gat));
  NAND3_X1  g678(.A1(new_n874_), .A2(new_n621_), .A3(new_n875_), .ZN(new_n880_));
  INV_X1    g679(.A(G176gat), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n819_), .A2(new_n616_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n866_), .A2(new_n881_), .A3(new_n586_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n880_), .A2(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(G1349gat));
  NAND2_X1  g683(.A1(new_n874_), .A2(new_n875_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n885_), .A2(new_n342_), .A3(new_n595_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n866_), .A2(new_n595_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G183gat), .B1(new_n882_), .B2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1350gat));
  OAI21_X1  g688(.A(G190gat), .B1(new_n885_), .B2(new_n644_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n289_), .A2(new_n343_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT125), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n885_), .B2(new_n892_), .ZN(G1351gat));
  AND2_X1   g692(.A1(new_n852_), .A2(new_n865_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n565_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g695(.A1(new_n852_), .A2(new_n865_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n586_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(G204gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n330_), .B2(new_n898_), .ZN(G1353gat));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n595_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n894_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n903_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n901_), .B1(new_n897_), .B2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n907_), .B(new_n909_), .ZN(G1354gat));
  OR3_X1    g709(.A1(new_n897_), .A2(G218gat), .A3(new_n642_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G218gat), .B1(new_n897_), .B2(new_n644_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1355gat));
endmodule


