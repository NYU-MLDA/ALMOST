//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT80), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G127gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G134gat), .ZN(new_n207_));
  INV_X1    g006(.A(G134gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(G127gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT80), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G113gat), .B(G120gat), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n205_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n205_), .B2(new_n210_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT83), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n220_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT2), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n226_), .B1(G141gat), .B2(G148gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(KEYINPUT2), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n225_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT84), .B1(new_n222_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(KEYINPUT2), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n226_), .A2(G141gat), .A3(G148gat), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n232_), .A2(new_n233_), .B1(new_n224_), .B2(new_n223_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n219_), .A2(new_n221_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT84), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n217_), .B1(new_n231_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT82), .ZN(new_n239_));
  OR3_X1    g038(.A1(new_n216_), .A2(new_n239_), .A3(KEYINPUT1), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n239_), .B1(new_n216_), .B2(KEYINPUT1), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n216_), .A2(KEYINPUT1), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n240_), .A2(new_n215_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n223_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n228_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n214_), .B1(new_n238_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n217_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n236_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n212_), .A2(new_n213_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(new_n245_), .A3(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n247_), .A2(KEYINPUT4), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n245_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n214_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n202_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G1gat), .B(G29gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(G85gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G57gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n202_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n265_));
  OR3_X1    g064(.A1(new_n258_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n263_), .B1(new_n258_), .B2(new_n265_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n252_), .B(KEYINPUT31), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT79), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(G43gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(KEYINPUT79), .A3(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(G15gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT30), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n281_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n275_), .A2(new_n276_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT78), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT23), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(G176gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n285_), .B(new_n287_), .C1(new_n294_), .C2(KEYINPUT24), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT24), .B1(new_n291_), .B2(new_n292_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n286_), .B(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT78), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G183gat), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT26), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n301_), .A2(KEYINPUT25), .B1(new_n303_), .B2(G190gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(KEYINPUT76), .B(G190gat), .Z(new_n305_));
  OAI211_X1 g104(.A(new_n302_), .B(new_n304_), .C1(new_n305_), .C2(new_n303_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n294_), .A2(KEYINPUT24), .A3(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n295_), .A2(new_n299_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(G169gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n305_), .A2(G183gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n298_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT81), .Z(new_n315_));
  AND3_X1   g114(.A1(new_n282_), .A2(new_n284_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n315_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n269_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n255_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G22gat), .B(G50gat), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n321_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G78gat), .ZN(new_n325_));
  INV_X1    g124(.A(G204gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n326_), .A2(G197gat), .ZN(new_n327_));
  INV_X1    g126(.A(G197gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n328_), .A2(G204gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT21), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G211gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(G218gat), .ZN(new_n332_));
  INV_X1    g131(.A(G218gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(G211gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n326_), .B2(G197gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n326_), .A2(G197gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n328_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n330_), .B(new_n335_), .C1(new_n340_), .C2(KEYINPUT21), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT88), .B1(new_n332_), .B2(new_n334_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n333_), .A2(G211gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n331_), .A2(G218gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT88), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n342_), .A2(new_n340_), .A3(KEYINPUT21), .A4(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n325_), .B(new_n349_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n320_), .B1(new_n251_), .B2(new_n245_), .ZN(new_n351_));
  OAI21_X1  g150(.A(G78gat), .B1(new_n351_), .B2(new_n348_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(G106gat), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(G106gat), .B1(new_n350_), .B2(new_n352_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n324_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n352_), .ZN(new_n357_));
  INV_X1    g156(.A(G106gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n321_), .B(new_n322_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n353_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n349_), .A2(new_n363_), .B1(G228gat), .B2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n356_), .A2(new_n366_), .A3(new_n361_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT20), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n287_), .B1(G183gat), .B2(G190gat), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n372_), .A2(new_n311_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT89), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(KEYINPUT24), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT24), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(KEYINPUT89), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n293_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n286_), .A2(KEYINPUT23), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n297_), .A2(G183gat), .A3(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT90), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n307_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n388_), .A2(new_n293_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n303_), .A2(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT26), .ZN(new_n392_));
  AND2_X1   g191(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n390_), .B(new_n392_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n389_), .B(new_n395_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n374_), .B1(new_n387_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n371_), .B1(new_n397_), .B2(new_n349_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT97), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT19), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n309_), .A2(new_n348_), .A3(new_n313_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n398_), .A2(new_n399_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n395_), .B1(new_n388_), .B2(new_n293_), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n379_), .A2(new_n293_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(KEYINPUT90), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n373_), .B1(new_n407_), .B2(new_n386_), .ZN(new_n408_));
  OAI211_X1 g207(.A(KEYINPUT20), .B(new_n403_), .C1(new_n408_), .C2(new_n348_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT97), .B1(new_n409_), .B2(new_n401_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n314_), .A2(new_n349_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n348_), .B(new_n374_), .C1(new_n387_), .C2(new_n396_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n411_), .A2(new_n412_), .A3(KEYINPUT20), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n404_), .B(new_n410_), .C1(new_n402_), .C2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT18), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n416_), .B(new_n417_), .Z(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n409_), .A2(new_n401_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n411_), .A2(new_n412_), .A3(KEYINPUT20), .A4(new_n402_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(KEYINPUT91), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT91), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n409_), .A2(new_n424_), .A3(new_n401_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n419_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n420_), .B1(KEYINPUT98), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(KEYINPUT98), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT27), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n423_), .A2(new_n419_), .A3(new_n425_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n431_), .A2(new_n426_), .A3(KEYINPUT27), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AOI211_X1 g232(.A(new_n318_), .B(new_n370_), .C1(new_n430_), .C2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n414_), .A2(KEYINPUT32), .A3(new_n418_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n423_), .A2(new_n425_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT32), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n436_), .B1(new_n437_), .B2(new_n419_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n438_), .A3(new_n268_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT92), .B1(new_n431_), .B2(new_n426_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n418_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT92), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n423_), .A2(new_n419_), .A3(new_n425_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT96), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n254_), .A2(new_n202_), .A3(new_n257_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n247_), .A2(new_n264_), .A3(new_n253_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(KEYINPUT95), .A3(new_n262_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT95), .B1(new_n448_), .B2(new_n262_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n446_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n451_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n453_), .A2(KEYINPUT96), .A3(new_n447_), .A4(new_n449_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(KEYINPUT33), .B(new_n263_), .C1(new_n258_), .C2(new_n265_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT94), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n267_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n457_), .B1(new_n267_), .B2(new_n458_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n455_), .B(new_n456_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n439_), .B1(new_n445_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n370_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n268_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT27), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT98), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n441_), .A2(new_n467_), .B1(new_n419_), .B2(new_n414_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n468_), .B2(new_n428_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n465_), .B1(new_n469_), .B2(new_n432_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n464_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n316_), .A2(new_n317_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n434_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT73), .B(G8gat), .Z(new_n474_));
  INV_X1    g273(.A(G1gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G8gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n476_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G29gat), .B(G36gat), .Z(new_n484_));
  XOR2_X1   g283(.A(G43gat), .B(G50gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n483_), .B(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G229gat), .A2(G233gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n486_), .B(KEYINPUT15), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(new_n482_), .A3(new_n481_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n487_), .A2(new_n489_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G113gat), .B(G141gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT74), .ZN(new_n495_));
  XOR2_X1   g294(.A(G169gat), .B(G197gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n493_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n483_), .B(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G78gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n325_), .A3(new_n503_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n505_), .A2(new_n506_), .B1(KEYINPUT11), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(KEYINPUT11), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n505_), .A2(new_n506_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n501_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n514_));
  XOR2_X1   g313(.A(G127gat), .B(G155gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT16), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G183gat), .B(G211gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n513_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(KEYINPUT17), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n513_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT10), .B(G99gat), .Z(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n358_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(KEYINPUT9), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT6), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n528_), .A2(KEYINPUT9), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n525_), .A2(new_n529_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT65), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n527_), .A2(new_n535_), .A3(new_n528_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n528_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT65), .B1(new_n537_), .B2(new_n526_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT7), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n530_), .A2(KEYINPUT6), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n530_), .A2(KEYINPUT6), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n542_), .B(new_n543_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT64), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n539_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(KEYINPUT8), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT8), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n542_), .A2(new_n543_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT64), .B1(new_n551_), .B2(new_n531_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n552_), .B2(new_n539_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT67), .B1(new_n549_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n548_), .A2(KEYINPUT8), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n550_), .A3(new_n539_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n534_), .B1(new_n554_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n511_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n534_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n560_), .B1(new_n563_), .B2(new_n511_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n511_), .ZN(new_n565_));
  OAI22_X1  g364(.A1(new_n559_), .A2(new_n562_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT68), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n511_), .B(new_n533_), .C1(new_n549_), .C2(new_n553_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n568_), .B1(new_n571_), .B2(new_n565_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n558_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n557_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n533_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n561_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n533_), .B1(new_n549_), .B2(new_n553_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n511_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n571_), .B2(new_n560_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT68), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n576_), .A2(new_n580_), .A3(new_n581_), .A4(new_n567_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n569_), .A2(new_n572_), .A3(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G120gat), .B(G148gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n569_), .A2(new_n572_), .A3(new_n582_), .A4(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT13), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT72), .ZN(new_n594_));
  INV_X1    g393(.A(new_n491_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT70), .B1(new_n559_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT70), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n575_), .A2(new_n597_), .A3(new_n491_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT34), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(KEYINPUT35), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n563_), .B2(new_n486_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(KEYINPUT35), .B(new_n601_), .C1(new_n604_), .C2(KEYINPUT71), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n599_), .A2(new_n605_), .A3(new_n603_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n599_), .B2(new_n603_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n594_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(G190gat), .B(G218gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n612_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  OAI221_X1 g416(.A(new_n594_), .B1(new_n617_), .B2(new_n613_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n616_), .A2(KEYINPUT37), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT37), .B1(new_n616_), .B2(new_n618_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n523_), .B(new_n593_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n473_), .A2(new_n499_), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n475_), .A3(new_n268_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n624_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(KEYINPUT38), .A3(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT100), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT38), .B1(new_n625_), .B2(new_n626_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n616_), .A2(new_n618_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n593_), .A2(new_n498_), .A3(new_n523_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n473_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n475_), .B1(new_n632_), .B2(new_n268_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n628_), .A2(new_n634_), .ZN(G1324gat));
  NAND2_X1  g434(.A1(new_n430_), .A2(new_n433_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n622_), .A2(new_n474_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n637_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G8gat), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(KEYINPUT39), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(KEYINPUT39), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n638_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g443(.A(new_n472_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n279_), .B1(new_n632_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT41), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n622_), .A2(new_n279_), .A3(new_n645_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1326gat));
  INV_X1    g448(.A(G22gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n632_), .B2(new_n370_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT42), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n622_), .A2(new_n650_), .A3(new_n370_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1327gat));
  INV_X1    g453(.A(new_n318_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n636_), .A2(new_n463_), .A3(new_n655_), .ZN(new_n656_));
  AOI22_X1  g455(.A1(new_n465_), .A2(new_n636_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(new_n645_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n593_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n630_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n659_), .A2(new_n660_), .A3(new_n523_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n658_), .A2(new_n498_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G29gat), .B1(new_n662_), .B2(new_n268_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n619_), .A2(new_n620_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n645_), .B1(new_n464_), .B2(new_n470_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n664_), .B(new_n665_), .C1(new_n666_), .C2(new_n434_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n658_), .A2(KEYINPUT101), .A3(new_n664_), .A4(new_n665_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n665_), .ZN(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT43), .B1(new_n473_), .B2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n670_), .A3(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n593_), .A2(new_n498_), .A3(new_n522_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n673_), .A2(KEYINPUT44), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT44), .B1(new_n673_), .B2(new_n675_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n268_), .A2(G29gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n663_), .B1(new_n678_), .B2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n662_), .A2(new_n681_), .A3(new_n637_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT45), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n676_), .A2(new_n677_), .A3(new_n636_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(new_n681_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n683_), .B(KEYINPUT46), .C1(new_n684_), .C2(new_n681_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1329gat));
  NAND2_X1  g488(.A1(new_n662_), .A2(new_n645_), .ZN(new_n690_));
  INV_X1    g489(.A(G43gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT102), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR4_X1   g493(.A1(new_n676_), .A2(new_n677_), .A3(new_n691_), .A4(new_n472_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT47), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n678_), .A2(G43gat), .A3(new_n645_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n693_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1330gat));
  INV_X1    g499(.A(G50gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n662_), .A2(new_n701_), .A3(new_n370_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n677_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n673_), .A2(KEYINPUT44), .A3(new_n675_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n370_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(new_n706_), .A3(G50gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(G50gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n702_), .B1(new_n707_), .B2(new_n708_), .ZN(G1331gat));
  NOR2_X1   g508(.A1(new_n473_), .A2(new_n498_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT37), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n630_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n616_), .A2(KEYINPUT37), .A3(new_n618_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n522_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n710_), .A2(new_n714_), .A3(new_n659_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n268_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n659_), .A2(new_n499_), .A3(new_n523_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n473_), .A2(new_n630_), .A3(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(G57gat), .A3(new_n268_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT104), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(KEYINPUT104), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n717_), .A2(new_n721_), .A3(new_n722_), .ZN(G1332gat));
  OR3_X1    g522(.A1(new_n715_), .A2(G64gat), .A3(new_n636_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n719_), .A2(new_n637_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G64gat), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT105), .B(KEYINPUT48), .Z(new_n729_));
  AND2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n729_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n724_), .B1(new_n730_), .B2(new_n731_), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n719_), .B2(new_n645_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT49), .Z(new_n735_));
  NAND2_X1  g534(.A1(new_n645_), .A2(new_n733_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT107), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n715_), .B2(new_n737_), .ZN(G1334gat));
  AOI21_X1  g537(.A(new_n325_), .B1(new_n719_), .B2(new_n370_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT50), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n716_), .A2(new_n325_), .A3(new_n370_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1335gat));
  NOR3_X1   g541(.A1(new_n660_), .A2(new_n593_), .A3(new_n523_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n710_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(G85gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n268_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n593_), .A2(new_n498_), .A3(new_n523_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n673_), .A2(new_n268_), .A3(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n749_), .B2(new_n746_), .ZN(G1336gat));
  AOI21_X1  g549(.A(G92gat), .B1(new_n745_), .B2(new_n637_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT108), .Z(new_n752_));
  NAND4_X1  g551(.A1(new_n673_), .A2(G92gat), .A3(new_n637_), .A4(new_n748_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1337gat));
  NAND3_X1  g553(.A1(new_n745_), .A2(new_n645_), .A3(new_n524_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n673_), .A2(new_n645_), .A3(new_n748_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n756_), .A2(KEYINPUT109), .A3(G99gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT109), .B1(new_n756_), .B2(G99gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n755_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT51), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT111), .Z(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n759_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n762_), .B(new_n755_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n745_), .A2(new_n358_), .A3(new_n370_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n673_), .A2(new_n370_), .A3(new_n748_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(G106gat), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n767_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n569_), .A2(new_n777_), .A3(new_n582_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n576_), .A2(new_n580_), .A3(KEYINPUT55), .A4(new_n567_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n566_), .A2(new_n568_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n782_), .B2(new_n589_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n784_), .B(new_n588_), .C1(new_n778_), .C2(new_n781_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n497_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n488_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n492_), .A2(new_n788_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n493_), .A2(new_n497_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n591_), .B2(new_n790_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n591_), .A2(new_n786_), .A3(new_n790_), .ZN(new_n792_));
  OAI22_X1  g591(.A1(new_n783_), .A2(new_n785_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT58), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  OAI221_X1 g594(.A(new_n795_), .B1(new_n792_), .B2(new_n791_), .C1(new_n783_), .C2(new_n785_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n665_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n591_), .A2(new_n498_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n782_), .A2(new_n589_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n784_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n782_), .A2(KEYINPUT56), .A3(new_n589_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n799_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n592_), .A2(new_n790_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n660_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(KEYINPUT114), .A3(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT57), .B(new_n660_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n798_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT114), .B1(new_n806_), .B2(new_n807_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n522_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n714_), .A2(new_n813_), .A3(new_n499_), .A4(new_n593_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT113), .ZN(new_n815_));
  INV_X1    g614(.A(new_n621_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n813_), .A4(new_n499_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n621_), .B2(new_n498_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n812_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n636_), .A2(new_n463_), .A3(new_n268_), .A4(new_n645_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT116), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT59), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n797_), .A2(new_n665_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n809_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n806_), .A2(new_n807_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n798_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n522_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n820_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n823_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n825_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837_), .B2(new_n499_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n823_), .ZN(new_n841_));
  AOI211_X1 g640(.A(KEYINPUT117), .B(new_n841_), .C1(new_n812_), .C2(new_n820_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n499_), .A2(G113gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n838_), .B1(new_n844_), .B2(new_n845_), .ZN(G1340gat));
  OAI21_X1  g645(.A(G120gat), .B1(new_n837_), .B2(new_n593_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n848_));
  AOI21_X1  g647(.A(G120gat), .B1(new_n659_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n848_), .B2(G120gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT120), .B1(new_n843_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852_));
  INV_X1    g651(.A(new_n850_), .ZN(new_n853_));
  NOR4_X1   g652(.A1(new_n840_), .A2(new_n842_), .A3(new_n852_), .A4(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n847_), .B1(new_n851_), .B2(new_n854_), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n837_), .B2(new_n522_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n843_), .A2(new_n206_), .A3(new_n523_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1342gat));
  XOR2_X1   g657(.A(KEYINPUT121), .B(G134gat), .Z(new_n859_));
  NOR3_X1   g658(.A1(new_n837_), .A2(new_n671_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G134gat), .B1(new_n843_), .B2(new_n630_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1343gat));
  AOI21_X1  g661(.A(new_n645_), .B1(new_n812_), .B2(new_n820_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n637_), .A2(new_n463_), .A3(new_n269_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n498_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g667(.A1(new_n865_), .A2(new_n593_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT122), .B(G148gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1345gat));
  NOR2_X1   g670(.A1(new_n865_), .A2(new_n522_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT61), .B(G155gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  OR3_X1    g673(.A1(new_n865_), .A2(G162gat), .A3(new_n660_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G162gat), .B1(new_n865_), .B2(new_n671_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1347gat));
  INV_X1    g676(.A(KEYINPUT22), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n637_), .A2(new_n655_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT123), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n370_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n832_), .A2(new_n878_), .A3(new_n498_), .A4(new_n881_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n882_), .A2(KEYINPUT62), .A3(new_n289_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(KEYINPUT62), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n832_), .A2(new_n498_), .A3(new_n881_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n289_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n883_), .B1(new_n884_), .B2(new_n887_), .ZN(G1348gat));
  NAND2_X1  g687(.A1(new_n832_), .A2(new_n881_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n290_), .B1(new_n889_), .B2(new_n593_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT124), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n892_), .B(new_n290_), .C1(new_n889_), .C2(new_n593_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n370_), .B1(new_n812_), .B2(new_n820_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n880_), .A2(new_n290_), .A3(new_n593_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n891_), .A2(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  OR2_X1    g695(.A1(new_n393_), .A2(new_n394_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n522_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n880_), .A2(new_n522_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n894_), .A2(new_n899_), .ZN(new_n900_));
  OAI221_X1 g699(.A(KEYINPUT125), .B1(new_n889_), .B2(new_n898_), .C1(new_n900_), .C2(G183gat), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n889_), .A2(new_n898_), .ZN(new_n903_));
  AOI21_X1  g702(.A(G183gat), .B1(new_n894_), .B2(new_n899_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n901_), .A2(new_n905_), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n889_), .B2(new_n671_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n630_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n889_), .B2(new_n908_), .ZN(G1351gat));
  NOR3_X1   g708(.A1(new_n636_), .A2(new_n463_), .A3(new_n268_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n863_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n912_), .B(new_n498_), .C1(KEYINPUT126), .C2(G197gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT126), .B(G197gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(new_n911_), .B2(new_n499_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1352gat));
  NOR2_X1   g715(.A1(new_n911_), .A2(new_n593_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(new_n326_), .ZN(G1353gat));
  AOI21_X1  g717(.A(new_n522_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n912_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT127), .Z(new_n922_));
  XNOR2_X1  g721(.A(new_n920_), .B(new_n922_), .ZN(G1354gat));
  OAI21_X1  g722(.A(G218gat), .B1(new_n911_), .B2(new_n671_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n630_), .A2(new_n333_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n911_), .B2(new_n925_), .ZN(G1355gat));
endmodule


