//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT21), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(KEYINPUT21), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  INV_X1    g007(.A(KEYINPUT85), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NOR3_X1   g011(.A1(KEYINPUT82), .A2(G169gat), .A3(G176gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n210_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n210_), .B1(G169gat), .B2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT82), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n211_), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n214_), .A2(new_n219_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT80), .B1(new_n229_), .B2(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G183gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT25), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(G183gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT80), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n227_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G190gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT26), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G190gat), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n230_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n229_), .A2(G183gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n232_), .A2(KEYINPUT25), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(KEYINPUT81), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n226_), .B1(new_n236_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT83), .B(G176gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT22), .B(G169gat), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n248_), .A2(new_n249_), .B1(G169gat), .B2(G176gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n232_), .A2(new_n237_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n217_), .A2(new_n218_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT84), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n217_), .A2(new_n251_), .A3(KEYINPUT84), .A4(new_n218_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n209_), .B1(new_n247_), .B2(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n214_), .A2(new_n219_), .A3(new_n225_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT81), .B1(new_n241_), .B2(new_n245_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n231_), .A2(new_n235_), .A3(new_n227_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(KEYINPUT85), .A3(new_n256_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n208_), .B1(new_n258_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT19), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT25), .B(G183gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n228_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT95), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n210_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n219_), .B2(new_n270_), .ZN(new_n271_));
  AND4_X1   g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n225_), .B(new_n268_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n250_), .A2(new_n252_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n206_), .B(new_n207_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT20), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n264_), .A2(new_n266_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n266_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n258_), .A2(new_n263_), .A3(new_n208_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT20), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(KEYINPUT96), .B(KEYINPUT18), .Z(new_n284_));
  XNOR2_X1  g083(.A(G8gat), .B(G36gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n278_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n280_), .A2(new_n282_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n266_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n258_), .A2(new_n263_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n276_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n277_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n279_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n290_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n202_), .B1(new_n289_), .B2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n291_), .A2(new_n266_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n279_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n288_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n292_), .A2(new_n296_), .A3(new_n290_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(KEYINPUT27), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT103), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G22gat), .B(G50gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n307_), .B(KEYINPUT28), .Z(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT2), .ZN(new_n313_));
  AND3_X1   g112(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT90), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(KEYINPUT90), .B(new_n313_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT91), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT91), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT89), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NOR4_X1   g129(.A1(KEYINPUT89), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n325_), .B(new_n326_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n312_), .B1(new_n320_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n311_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(new_n328_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n310_), .A2(new_n334_), .A3(new_n311_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT87), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n336_), .A2(new_n337_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT88), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n336_), .A2(KEYINPUT88), .A3(new_n342_), .A4(new_n337_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT92), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n333_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n333_), .B2(new_n347_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n309_), .B1(new_n351_), .B2(KEYINPUT29), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT29), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(new_n308_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G78gat), .B(G106gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G228gat), .A2(G233gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT93), .Z(new_n358_));
  NOR3_X1   g157(.A1(new_n349_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n208_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n333_), .A2(new_n347_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT29), .ZN(new_n362_));
  INV_X1    g161(.A(new_n358_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(new_n276_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n356_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(KEYINPUT92), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n333_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(KEYINPUT29), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n363_), .B1(new_n368_), .B2(new_n276_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n356_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n364_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(KEYINPUT94), .B(new_n355_), .C1(new_n365_), .C2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n355_), .A2(KEYINPUT94), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n360_), .A2(new_n356_), .A3(new_n364_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n370_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT94), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n352_), .A2(new_n354_), .A3(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .A4(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n298_), .A2(new_n303_), .A3(KEYINPUT103), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n306_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G15gat), .B(G43gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  AND3_X1   g186(.A1(new_n258_), .A2(new_n263_), .A3(KEYINPUT30), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT30), .B1(new_n258_), .B2(new_n263_), .ZN(new_n389_));
  OR3_X1    g188(.A1(new_n388_), .A2(new_n389_), .A3(KEYINPUT86), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT86), .B1(new_n388_), .B2(new_n389_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n387_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n387_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G134gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G127gat), .ZN(new_n396_));
  INV_X1    g195(.A(G127gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G134gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G120gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G113gat), .ZN(new_n401_));
  INV_X1    g200(.A(G113gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G120gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n399_), .A2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n396_), .A2(new_n398_), .A3(new_n401_), .A4(new_n403_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n407_), .B(KEYINPUT31), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  OR3_X1    g208(.A1(new_n392_), .A2(new_n394_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n409_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT101), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414_));
  INV_X1    g213(.A(new_n407_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n366_), .A2(new_n414_), .A3(new_n367_), .A4(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT97), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n405_), .A2(new_n406_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n333_), .A3(new_n347_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT98), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT98), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n423_), .A2(new_n333_), .A3(new_n347_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n366_), .A2(new_n367_), .A3(new_n415_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(KEYINPUT4), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n351_), .A2(new_n415_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n419_), .A2(new_n430_), .B1(new_n431_), .B2(new_n417_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G1gat), .B(G29gat), .Z(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT0), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G57gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G85gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n413_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n428_), .A2(new_n429_), .A3(new_n417_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n428_), .A2(new_n429_), .A3(KEYINPUT4), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n416_), .A2(new_n418_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G85gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n435_), .B(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(KEYINPUT101), .A3(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n438_), .B(new_n436_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n437_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n412_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n382_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT102), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n416_), .A2(new_n417_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n431_), .B2(KEYINPUT4), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n428_), .A2(new_n429_), .A3(new_n418_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n443_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT100), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n436_), .B1(new_n431_), .B2(new_n418_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT100), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n430_), .A2(new_n417_), .A3(new_n416_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n456_), .A2(new_n460_), .B1(new_n445_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n288_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n302_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n445_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n464_), .B1(new_n465_), .B2(KEYINPUT33), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n462_), .A2(new_n466_), .B1(new_n373_), .B2(new_n379_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n299_), .A2(new_n300_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n292_), .A2(new_n296_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n290_), .A2(KEYINPUT32), .ZN(new_n470_));
  MUX2_X1   g269(.A(new_n468_), .B(new_n469_), .S(new_n470_), .Z(new_n471_));
  NAND3_X1  g270(.A1(new_n430_), .A2(new_n418_), .A3(new_n416_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n436_), .B1(new_n472_), .B2(new_n438_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n445_), .B1(new_n473_), .B2(KEYINPUT101), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n432_), .A2(new_n413_), .A3(new_n436_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n471_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n412_), .B1(new_n467_), .B2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n373_), .B(new_n379_), .C1(new_n446_), .C2(new_n304_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n451_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n456_), .A2(new_n460_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n289_), .A2(new_n297_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n432_), .A2(KEYINPUT33), .A3(new_n436_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n445_), .A2(new_n461_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n476_), .A2(new_n484_), .A3(new_n380_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n412_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n451_), .A3(new_n478_), .A4(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n450_), .B1(new_n479_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT9), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(G85gat), .A3(G92gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G85gat), .B(G92gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT10), .B(G99gat), .ZN(new_n493_));
  OAI221_X1 g292(.A(new_n491_), .B1(new_n492_), .B2(new_n490_), .C1(G106gat), .C2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n499_), .A2(KEYINPUT8), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n494_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n497_), .A2(new_n498_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT65), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT65), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n499_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n505_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT64), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n492_), .B(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(KEYINPUT8), .A3(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(KEYINPUT8), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n506_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G29gat), .B(G36gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT15), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT35), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT34), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n517_), .A2(new_n521_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n492_), .A2(KEYINPUT64), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n492_), .A2(KEYINPUT64), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(KEYINPUT8), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n504_), .B1(new_n509_), .B2(new_n499_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n529_), .B1(new_n508_), .B2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n504_), .B1(new_n494_), .B2(new_n500_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n515_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n520_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n526_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n525_), .A2(new_n522_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT70), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(KEYINPUT70), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n526_), .A2(KEYINPUT70), .A3(new_n534_), .A4(new_n536_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G190gat), .B(G218gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n539_), .A2(KEYINPUT36), .A3(new_n540_), .A4(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(KEYINPUT36), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n540_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n545_), .ZN(new_n549_));
  AOI211_X1 g348(.A(KEYINPUT71), .B(new_n549_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n544_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n544_), .B(KEYINPUT37), .C1(new_n548_), .C2(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT76), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G127gat), .B(G155gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT17), .Z(new_n563_));
  XNOR2_X1  g362(.A(G71gat), .B(G78gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(G57gat), .B(G64gat), .Z(new_n565_));
  INV_X1    g364(.A(KEYINPUT11), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G57gat), .B(G64gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT11), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n564_), .A3(KEYINPUT11), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT72), .B(G15gat), .ZN(new_n573_));
  INV_X1    g372(.A(G22gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(G1gat), .ZN(new_n576_));
  INV_X1    g375(.A(G8gat), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT14), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G1gat), .B(G8gat), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT73), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n583_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n563_), .B1(new_n572_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n572_), .B2(new_n587_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT67), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n572_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT74), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n592_), .A2(new_n586_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n594_));
  NOR3_X1   g393(.A1(new_n593_), .A2(new_n562_), .A3(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n592_), .B2(new_n586_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n589_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n556_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n572_), .A2(new_n590_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT67), .B1(new_n570_), .B2(new_n571_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT12), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT68), .B1(new_n601_), .B2(new_n533_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT68), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n591_), .A2(new_n603_), .A3(KEYINPUT12), .A4(new_n517_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n570_), .A2(new_n571_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n517_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n517_), .A2(new_n606_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(G230gat), .ZN(new_n611_));
  INV_X1    g410(.A(G233gat), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n605_), .A2(new_n610_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n607_), .B2(KEYINPUT66), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT66), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n609_), .A2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n616_), .B1(new_n607_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621_));
  INV_X1    g420(.A(G204gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT5), .B(G176gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT69), .Z(new_n626_));
  AND2_X1   g425(.A1(new_n620_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n615_), .A2(new_n619_), .A3(new_n625_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OR3_X1    g428(.A1(new_n627_), .A2(KEYINPUT13), .A3(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT13), .B1(new_n627_), .B2(new_n629_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n581_), .A2(new_n582_), .A3(new_n520_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT78), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT78), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n581_), .A2(new_n635_), .A3(new_n582_), .A4(new_n520_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n520_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n634_), .A2(new_n636_), .B1(new_n583_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G229gat), .A2(G233gat), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT79), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n634_), .A2(new_n636_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n583_), .A2(new_n521_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n639_), .A3(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT79), .B1(new_n638_), .B2(new_n639_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G113gat), .B(G141gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(G169gat), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(G197gat), .Z(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n642_), .A2(new_n646_), .A3(new_n645_), .A4(new_n650_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n632_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n489_), .A2(new_n598_), .A3(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n576_), .A3(new_n446_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n446_), .A2(new_n471_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n453_), .A2(KEYINPUT100), .A3(new_n455_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n458_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n483_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n482_), .A2(new_n481_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n380_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n478_), .B(new_n486_), .C1(new_n661_), .C2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT102), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n449_), .B1(new_n668_), .B2(new_n487_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n551_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n655_), .A2(new_n597_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G1gat), .B1(new_n672_), .B2(new_n447_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n658_), .A2(new_n659_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n660_), .A2(new_n673_), .A3(new_n674_), .ZN(G1324gat));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  INV_X1    g475(.A(new_n551_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n306_), .A2(new_n381_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n489_), .A2(new_n677_), .A3(new_n679_), .A4(new_n671_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G8gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT39), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n678_), .A2(G8gat), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n489_), .A2(new_n598_), .A3(new_n656_), .A4(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT104), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n682_), .A2(new_n683_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n683_), .B1(new_n682_), .B2(new_n686_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n676_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n682_), .A2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT105), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n682_), .A2(new_n683_), .A3(new_n686_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(KEYINPUT40), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n689_), .A2(new_n693_), .ZN(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n672_), .B2(new_n486_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT41), .Z(new_n696_));
  INV_X1    g495(.A(G15gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n657_), .A2(new_n697_), .A3(new_n412_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1326gat));
  OAI21_X1  g498(.A(G22gat), .B1(new_n672_), .B2(new_n380_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT42), .ZN(new_n701_));
  INV_X1    g500(.A(new_n380_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n657_), .A2(new_n574_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1327gat));
  INV_X1    g503(.A(new_n597_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n677_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n489_), .A2(new_n656_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G29gat), .B1(new_n707_), .B2(new_n446_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n656_), .A2(new_n597_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT106), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n669_), .B2(new_n555_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n489_), .A2(new_n712_), .A3(new_n556_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n709_), .B(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n712_), .B1(new_n489_), .B2(new_n556_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n669_), .A2(KEYINPUT43), .A3(new_n555_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n719_), .B(KEYINPUT44), .C1(new_n720_), .C2(new_n721_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n722_), .A2(G29gat), .A3(new_n446_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n708_), .B1(new_n717_), .B2(new_n723_), .ZN(G1328gat));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n679_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G36gat), .B1(new_n716_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(G36gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n707_), .A2(new_n727_), .A3(new_n679_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT45), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n726_), .A2(KEYINPUT46), .A3(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1329gat));
  NAND3_X1  g533(.A1(new_n722_), .A2(G43gat), .A3(new_n412_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n707_), .A2(new_n412_), .ZN(new_n736_));
  OAI22_X1  g535(.A1(new_n716_), .A2(new_n735_), .B1(G43gat), .B2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g537(.A(G50gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n707_), .A2(new_n739_), .A3(new_n702_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n722_), .B(new_n702_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n741_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT108), .B1(new_n741_), .B2(G50gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(G1331gat));
  NOR3_X1   g543(.A1(new_n632_), .A2(new_n597_), .A3(new_n654_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n670_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G57gat), .B1(new_n746_), .B2(new_n447_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n654_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n489_), .A2(KEYINPUT109), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(new_n669_), .B2(new_n654_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n632_), .B1(new_n749_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n598_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n447_), .A2(G57gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n747_), .B1(new_n753_), .B2(new_n754_), .ZN(G1332gat));
  OAI21_X1  g554(.A(G64gat), .B1(new_n746_), .B2(new_n678_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT48), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n678_), .A2(G64gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n753_), .B2(new_n758_), .ZN(G1333gat));
  OR3_X1    g558(.A1(new_n753_), .A2(G71gat), .A3(new_n486_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n670_), .A2(new_n412_), .A3(new_n745_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G71gat), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT110), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT110), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(KEYINPUT49), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT49), .B1(new_n763_), .B2(new_n764_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n760_), .B1(new_n765_), .B2(new_n766_), .ZN(G1334gat));
  OAI21_X1  g566(.A(G78gat), .B1(new_n746_), .B2(new_n380_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT50), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT50), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n380_), .A2(G78gat), .ZN(new_n771_));
  OAI22_X1  g570(.A1(new_n769_), .A2(new_n770_), .B1(new_n753_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT111), .ZN(G1335gat));
  NOR2_X1   g572(.A1(new_n705_), .A2(new_n654_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n630_), .A2(new_n631_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n713_), .B2(new_n711_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778_), .B2(new_n447_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n752_), .A2(new_n706_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n446_), .A2(new_n442_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(G1336gat));
  OAI21_X1  g581(.A(G92gat), .B1(new_n778_), .B2(new_n678_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n678_), .A2(G92gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n780_), .B2(new_n784_), .ZN(G1337gat));
  NOR3_X1   g584(.A1(new_n780_), .A2(new_n493_), .A3(new_n486_), .ZN(new_n786_));
  INV_X1    g585(.A(G99gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n777_), .B2(new_n412_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1338gat));
  INV_X1    g590(.A(new_n776_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n702_), .B(new_n792_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n793_));
  XOR2_X1   g592(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n794_));
  AND3_X1   g593(.A1(new_n793_), .A2(G106gat), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n793_), .B2(G106gat), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n794_), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n380_), .B(new_n776_), .C1(new_n713_), .C2(new_n711_), .ZN(new_n800_));
  INV_X1    g599(.A(G106gat), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n797_), .B(new_n799_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n752_), .A2(new_n801_), .A3(new_n702_), .A4(new_n706_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT53), .B1(new_n798_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n793_), .A2(G106gat), .A3(new_n794_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(KEYINPUT113), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n803_), .A4(new_n802_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n805_), .A2(new_n810_), .ZN(G1339gat));
  NOR3_X1   g610(.A1(new_n382_), .A2(new_n486_), .A3(new_n447_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n615_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n605_), .A2(new_n610_), .A3(KEYINPUT55), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n613_), .A2(KEYINPUT114), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n605_), .A2(new_n610_), .A3(KEYINPUT55), .A4(new_n816_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n814_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n626_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT56), .ZN(new_n822_));
  INV_X1    g621(.A(new_n639_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n643_), .A2(new_n823_), .A3(new_n644_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n824_), .B(new_n651_), .C1(new_n823_), .C2(new_n638_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n653_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n820_), .A2(new_n827_), .A3(new_n626_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n822_), .A2(new_n628_), .A3(new_n826_), .A4(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n556_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n555_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT115), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n629_), .B1(new_n821_), .B2(KEYINPUT56), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n837_), .A2(KEYINPUT58), .A3(new_n826_), .A4(new_n828_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n834_), .A2(new_n836_), .A3(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n822_), .A2(new_n654_), .A3(new_n628_), .A4(new_n828_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n826_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n551_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n705_), .B1(new_n839_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n654_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n598_), .B2(new_n847_), .ZN(new_n848_));
  AND4_X1   g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n705_), .A4(new_n555_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n812_), .B1(new_n845_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n402_), .B1(new_n851_), .B2(new_n748_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT116), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n840_), .A2(new_n841_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n677_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n843_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n842_), .A2(KEYINPUT57), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n838_), .B1(new_n835_), .B2(KEYINPUT115), .ZN(new_n858_));
  AOI211_X1 g657(.A(new_n833_), .B(new_n555_), .C1(new_n830_), .C2(new_n829_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n856_), .B(new_n857_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n597_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n850_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n812_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n864_), .A2(KEYINPUT118), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(KEYINPUT118), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n867_));
  NOR3_X1   g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n851_), .A2(KEYINPUT59), .B1(new_n863_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n870_), .A2(new_n402_), .A3(new_n748_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n853_), .A2(new_n871_), .ZN(G1340gat));
  AOI21_X1  g671(.A(new_n400_), .B1(new_n869_), .B2(new_n775_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n850_), .B1(new_n860_), .B2(new_n597_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n864_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n400_), .A2(KEYINPUT60), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n400_), .B1(new_n632_), .B2(KEYINPUT60), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT119), .B1(new_n873_), .B2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n863_), .A2(new_n868_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n881_), .B(new_n775_), .C1(new_n875_), .C2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G120gat), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n878_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n880_), .A2(new_n886_), .ZN(G1341gat));
  OAI21_X1  g686(.A(G127gat), .B1(new_n870_), .B2(new_n597_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n875_), .A2(new_n397_), .A3(new_n705_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1342gat));
  OAI21_X1  g689(.A(G134gat), .B1(new_n870_), .B2(new_n555_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n875_), .A2(new_n395_), .A3(new_n551_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1343gat));
  NOR4_X1   g692(.A1(new_n679_), .A2(new_n380_), .A3(new_n447_), .A4(new_n412_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n863_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n654_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n775_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g699(.A1(new_n895_), .A2(new_n597_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT61), .B(G155gat), .Z(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  OR3_X1    g702(.A1(new_n895_), .A2(G162gat), .A3(new_n677_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G162gat), .B1(new_n895_), .B2(new_n555_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n678_), .A2(new_n448_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n863_), .A2(new_n380_), .A3(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n249_), .A3(new_n654_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n874_), .A2(new_n702_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n907_), .A2(new_n654_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT120), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n911_), .B1(new_n915_), .B2(G169gat), .ZN(new_n916_));
  AOI211_X1 g715(.A(KEYINPUT62), .B(new_n222_), .C1(new_n912_), .C2(new_n914_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n910_), .B1(new_n916_), .B2(new_n917_), .ZN(G1348gat));
  NOR2_X1   g717(.A1(new_n908_), .A2(new_n632_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n248_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT121), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n922_), .B(new_n248_), .C1(new_n908_), .C2(new_n632_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n919_), .A2(G176gat), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n921_), .A2(new_n923_), .A3(new_n924_), .ZN(G1349gat));
  NAND2_X1  g724(.A1(new_n909_), .A2(new_n705_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(G183gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n267_), .B1(KEYINPUT122), .B2(G183gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n926_), .B2(new_n929_), .ZN(G1350gat));
  NOR2_X1   g729(.A1(new_n908_), .A2(new_n555_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n551_), .A2(new_n228_), .ZN(new_n932_));
  OAI22_X1  g731(.A1(new_n931_), .A2(new_n237_), .B1(new_n908_), .B2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  OAI221_X1 g734(.A(KEYINPUT123), .B1(new_n908_), .B2(new_n932_), .C1(new_n931_), .C2(new_n237_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1351gat));
  NOR2_X1   g736(.A1(new_n412_), .A2(new_n446_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n679_), .A2(new_n702_), .A3(new_n938_), .ZN(new_n939_));
  OAI21_X1  g738(.A(KEYINPUT124), .B1(new_n874_), .B2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941_));
  INV_X1    g740(.A(new_n939_), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n941_), .B(new_n942_), .C1(new_n845_), .C2(new_n850_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n940_), .A2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n654_), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT125), .B(G197gat), .Z(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n944_), .A2(new_n775_), .ZN(new_n948_));
  AOI21_X1  g747(.A(KEYINPUT126), .B1(new_n948_), .B2(G204gat), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n632_), .B1(new_n940_), .B2(new_n943_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n950_), .A2(new_n951_), .A3(new_n622_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953_));
  AND4_X1   g752(.A1(new_n953_), .A2(new_n944_), .A3(new_n622_), .A4(new_n775_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n953_), .B1(new_n950_), .B2(new_n622_), .ZN(new_n955_));
  OAI22_X1  g754(.A1(new_n949_), .A2(new_n952_), .B1(new_n954_), .B2(new_n955_), .ZN(G1353gat));
  OR2_X1    g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  NAND2_X1  g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  AND4_X1   g757(.A1(new_n705_), .A2(new_n944_), .A3(new_n957_), .A4(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n957_), .B1(new_n944_), .B2(new_n705_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n959_), .A2(new_n960_), .ZN(G1354gat));
  INV_X1    g760(.A(new_n944_), .ZN(new_n962_));
  OR3_X1    g761(.A1(new_n962_), .A2(G218gat), .A3(new_n677_), .ZN(new_n963_));
  OAI21_X1  g762(.A(G218gat), .B1(new_n962_), .B2(new_n555_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1355gat));
endmodule


