//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT66), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT10), .B(G99gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n210_), .B1(G106gat), .B2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n213_), .B1(new_n215_), .B2(KEYINPUT9), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n214_), .A2(KEYINPUT64), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT64), .B1(new_n214_), .B2(new_n217_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n216_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT65), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n216_), .B(new_n222_), .C1(new_n219_), .C2(new_n218_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n212_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n215_), .A2(new_n213_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT7), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT68), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(KEYINPUT67), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(KEYINPUT68), .B2(new_n229_), .ZN(new_n234_));
  OAI22_X1  g033(.A1(KEYINPUT67), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n232_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n228_), .B1(new_n210_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n226_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(new_n236_), .B2(new_n206_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n227_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT67), .B1(new_n242_), .B2(KEYINPUT7), .ZN(new_n243_));
  INV_X1    g042(.A(G99gat), .ZN(new_n244_));
  INV_X1    g043(.A(G106gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n233_), .A2(new_n229_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n248_), .A2(new_n232_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT69), .B1(new_n249_), .B2(new_n238_), .ZN(new_n250_));
  AOI211_X1 g049(.A(KEYINPUT71), .B(new_n237_), .C1(new_n241_), .C2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n234_), .A2(new_n235_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n243_), .A2(new_n246_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n206_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(new_n240_), .A3(new_n226_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n250_), .A2(new_n256_), .A3(KEYINPUT8), .ZN(new_n257_));
  INV_X1    g056(.A(new_n237_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n252_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n225_), .B1(new_n251_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G29gat), .B(G36gat), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n261_), .A2(KEYINPUT73), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(KEYINPUT73), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G43gat), .B(G50gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n262_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(KEYINPUT15), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT15), .ZN(new_n270_));
  INV_X1    g069(.A(new_n268_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n265_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n260_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G232gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT34), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(KEYINPUT35), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n257_), .A2(new_n258_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n225_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n267_), .A2(new_n268_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n277_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n276_), .A2(KEYINPUT35), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT72), .Z(new_n284_));
  NAND3_X1  g083(.A1(new_n274_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n274_), .B2(new_n282_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G190gat), .B(G218gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT74), .ZN(new_n289_));
  XOR2_X1   g088(.A(G134gat), .B(G162gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  OAI22_X1  g091(.A1(new_n286_), .A2(new_n287_), .B1(KEYINPUT36), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n274_), .A2(new_n282_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n284_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n292_), .A2(KEYINPUT36), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n285_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n293_), .A2(new_n298_), .B1(KEYINPUT36), .B2(new_n292_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT37), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n299_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G127gat), .B(G155gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT16), .ZN(new_n305_));
  XOR2_X1   g104(.A(G183gat), .B(G211gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT17), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G57gat), .B(G64gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G71gat), .B(G78gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(KEYINPUT11), .ZN(new_n313_));
  XOR2_X1   g112(.A(G71gat), .B(G78gat), .Z(new_n314_));
  INV_X1    g113(.A(G64gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G57gat), .ZN(new_n316_));
  INV_X1    g115(.A(G57gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G64gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n318_), .A3(KEYINPUT11), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n311_), .A2(KEYINPUT11), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n313_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT77), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G15gat), .B(G22gat), .ZN(new_n326_));
  INV_X1    g125(.A(G1gat), .ZN(new_n327_));
  INV_X1    g126(.A(G8gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT14), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G1gat), .B(G8gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G231gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  AOI211_X1 g133(.A(new_n309_), .B(new_n310_), .C1(new_n325_), .C2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n334_), .B2(new_n325_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n334_), .A2(new_n322_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n322_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n310_), .A3(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n339_), .A2(KEYINPUT76), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(KEYINPUT76), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n336_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n303_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT78), .ZN(new_n344_));
  XOR2_X1   g143(.A(G8gat), .B(G36gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT102), .ZN(new_n350_));
  INV_X1    g149(.A(G183gat), .ZN(new_n351_));
  INV_X1    g150(.A(G190gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT23), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT84), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(G183gat), .A3(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT85), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n363_), .A3(new_n360_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT83), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT25), .B(G183gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT26), .B(G190gat), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n366_), .A2(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n364_), .A3(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G211gat), .B(G218gat), .Z(new_n373_));
  INV_X1    g172(.A(G197gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(KEYINPUT94), .A3(G204gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT94), .ZN(new_n376_));
  INV_X1    g175(.A(G204gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n376_), .B1(new_n377_), .B2(G197gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT93), .B(G197gat), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n375_), .B(new_n378_), .C1(new_n379_), .C2(G204gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n373_), .B1(new_n380_), .B2(KEYINPUT21), .ZN(new_n381_));
  MUX2_X1   g180(.A(G197gat), .B(new_n379_), .S(G204gat), .Z(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(KEYINPUT21), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(KEYINPUT21), .A3(new_n373_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(G176gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT22), .ZN(new_n387_));
  OAI21_X1  g186(.A(G169gat), .B1(new_n387_), .B2(KEYINPUT86), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n387_), .A2(G169gat), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n386_), .B(new_n388_), .C1(new_n389_), .C2(KEYINPUT86), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n353_), .A2(new_n357_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n390_), .B(new_n366_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n372_), .A2(new_n385_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n358_), .B1(G183gat), .B2(G190gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT22), .B(G169gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n386_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n366_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT96), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  AOI211_X1 g202(.A(new_n359_), .B(new_n391_), .C1(new_n365_), .C2(new_n368_), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n369_), .B(KEYINPUT95), .Z(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n370_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n398_), .A2(new_n403_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT20), .B1(new_n407_), .B2(new_n385_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n395_), .A2(new_n397_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n397_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n372_), .A2(new_n393_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n383_), .A2(new_n384_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT20), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n407_), .B2(new_n385_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n350_), .B1(new_n409_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n410_), .A3(new_n415_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n395_), .A2(new_n408_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n418_), .B(new_n349_), .C1(new_n419_), .C2(new_n410_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(KEYINPUT27), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT103), .ZN(new_n422_));
  XOR2_X1   g221(.A(G155gat), .B(G162gat), .Z(new_n423_));
  INV_X1    g222(.A(KEYINPUT1), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(G141gat), .A2(G148gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT90), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G141gat), .A2(G148gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .A4(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n426_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT2), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n433_), .A2(new_n435_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n423_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n431_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT92), .B1(new_n440_), .B2(KEYINPUT29), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n412_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G228gat), .A2(G233gat), .ZN(new_n443_));
  INV_X1    g242(.A(G78gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(G106gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n442_), .B(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT91), .ZN(new_n449_));
  OR3_X1    g248(.A1(new_n440_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT28), .B1(new_n440_), .B2(KEYINPUT29), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G22gat), .B(G50gat), .Z(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n455_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n448_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n457_), .A3(new_n447_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT27), .ZN(new_n465_));
  INV_X1    g264(.A(new_n420_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n398_), .A2(new_n403_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n404_), .A2(new_n406_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n414_), .B1(new_n469_), .B2(new_n412_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n410_), .B1(new_n470_), .B2(new_n394_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n349_), .B1(new_n472_), .B2(new_n418_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n465_), .B1(new_n466_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT103), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n417_), .A2(new_n420_), .A3(new_n475_), .A4(KEYINPUT27), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n422_), .A2(new_n464_), .A3(new_n474_), .A4(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G15gat), .B(G43gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT87), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT30), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G227gat), .A2(G233gat), .ZN(new_n481_));
  INV_X1    g280(.A(G71gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(new_n244_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n411_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n411_), .A2(new_n484_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n480_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n487_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n480_), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n489_), .A2(new_n485_), .A3(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT89), .B1(new_n488_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n490_), .B1(new_n489_), .B2(new_n485_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n486_), .A2(new_n480_), .A3(new_n487_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G127gat), .B(G134gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT88), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G113gat), .B(G120gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n497_), .A2(KEYINPUT88), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(KEYINPUT88), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n499_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT31), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n492_), .A2(new_n496_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n501_), .A2(new_n431_), .A3(new_n439_), .A4(new_n504_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n440_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT98), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n509_), .B(KEYINPUT4), .C1(new_n510_), .C2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n505_), .A2(KEYINPUT98), .A3(new_n513_), .A4(new_n440_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n508_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G1gat), .B(G29gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(G85gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT0), .B(G57gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n510_), .A2(new_n509_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n508_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OR4_X1    g322(.A1(KEYINPUT101), .A2(new_n515_), .A3(new_n520_), .A4(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n512_), .A2(new_n514_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n508_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(new_n519_), .A3(new_n522_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n520_), .B1(new_n515_), .B2(new_n523_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT101), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n524_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n506_), .ZN(new_n532_));
  OAI211_X1 g331(.A(KEYINPUT89), .B(new_n532_), .C1(new_n488_), .C2(new_n491_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n507_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n477_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(KEYINPUT32), .B(new_n349_), .C1(new_n409_), .C2(new_n416_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n472_), .A2(new_n537_), .A3(new_n418_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n536_), .A2(new_n524_), .A3(new_n530_), .A4(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n519_), .B1(new_n521_), .B2(new_n508_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT100), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n512_), .A2(new_n508_), .A3(new_n514_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT33), .ZN(new_n544_));
  AOI22_X1  g343(.A1(new_n542_), .A2(new_n543_), .B1(new_n529_), .B2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n519_), .B1(new_n527_), .B2(new_n522_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(KEYINPUT99), .A3(KEYINPUT33), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT99), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n529_), .B2(new_n544_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n349_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n418_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(new_n471_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n420_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n539_), .B1(new_n550_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n464_), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n462_), .A2(new_n460_), .B1(new_n524_), .B2(new_n530_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n557_), .A2(new_n422_), .A3(new_n476_), .A4(new_n474_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n507_), .A2(new_n533_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n535_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n237_), .B1(new_n241_), .B2(new_n250_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n562_), .A2(new_n324_), .A3(new_n224_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT12), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n324_), .B1(new_n562_), .B2(new_n224_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n322_), .A2(new_n564_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n260_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n279_), .A2(new_n324_), .ZN(new_n572_));
  OAI211_X1 g371(.A(G230gat), .B(G233gat), .C1(new_n572_), .C2(new_n563_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n578_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n571_), .A2(new_n573_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT13), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n579_), .A2(KEYINPUT13), .A3(new_n581_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n332_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n281_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n267_), .A2(new_n332_), .A3(new_n268_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(KEYINPUT79), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT79), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n267_), .A2(new_n332_), .A3(new_n593_), .A4(new_n268_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n273_), .A2(new_n269_), .A3(new_n332_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n591_), .A3(new_n588_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G113gat), .B(G141gat), .Z(new_n599_));
  XOR2_X1   g398(.A(G169gat), .B(G197gat), .Z(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT80), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n598_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n595_), .A2(new_n597_), .A3(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT81), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT81), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n595_), .A2(new_n597_), .A3(new_n606_), .A4(new_n601_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n603_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(KEYINPUT82), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n607_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n603_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n610_), .A2(KEYINPUT82), .A3(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n561_), .A2(new_n586_), .A3(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n344_), .A2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n531_), .B(KEYINPUT104), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n327_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n293_), .A2(new_n298_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n292_), .A2(KEYINPUT36), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n561_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n586_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n342_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n608_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n628_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n623_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n632_), .B2(new_n531_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n617_), .A2(new_n618_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n619_), .A2(new_n633_), .A3(new_n634_), .ZN(G1324gat));
  NAND3_X1  g434(.A1(new_n422_), .A2(new_n476_), .A3(new_n474_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n615_), .A2(new_n328_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n631_), .A2(new_n636_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(G8gat), .ZN(new_n640_));
  AOI211_X1 g439(.A(KEYINPUT39), .B(new_n328_), .C1(new_n631_), .C2(new_n636_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1325gat));
  OAI21_X1  g443(.A(G15gat), .B1(new_n632_), .B2(new_n560_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n645_), .A2(KEYINPUT41), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(KEYINPUT41), .ZN(new_n647_));
  INV_X1    g446(.A(G15gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n560_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n615_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n646_), .A2(new_n647_), .A3(new_n650_), .ZN(G1326gat));
  OAI21_X1  g450(.A(G22gat), .B1(new_n632_), .B2(new_n464_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT42), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n464_), .A2(G22gat), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT106), .Z(new_n655_));
  NAND2_X1  g454(.A1(new_n615_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(G1327gat));
  NOR2_X1   g456(.A1(new_n299_), .A2(new_n625_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n614_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n531_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G29gat), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n586_), .A2(new_n625_), .A3(new_n608_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n466_), .A2(new_n473_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n665_), .A2(new_n547_), .A3(new_n549_), .A4(new_n545_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n463_), .B1(new_n666_), .B2(new_n539_), .ZN(new_n667_));
  AND4_X1   g466(.A1(new_n557_), .A2(new_n422_), .A3(new_n476_), .A4(new_n474_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n560_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n535_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n664_), .B1(new_n671_), .B2(new_n303_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n622_), .B(new_n302_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n561_), .A2(new_n673_), .A3(KEYINPUT43), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n663_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n671_), .A2(new_n664_), .A3(new_n303_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n561_), .B2(new_n673_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n676_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(new_n663_), .A3(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n677_), .A2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n616_), .A2(G29gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n662_), .B1(new_n683_), .B2(new_n684_), .ZN(G1328gat));
  AND2_X1   g484(.A1(new_n636_), .A2(KEYINPUT108), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n636_), .A2(KEYINPUT108), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(G36gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n659_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n677_), .A2(new_n636_), .A3(new_n682_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n690_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  OAI221_X1 g498(.A(new_n694_), .B1(new_n697_), .B2(KEYINPUT46), .C1(new_n695_), .C2(new_n690_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1329gat));
  INV_X1    g500(.A(G43gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n560_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n677_), .A2(new_n682_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n677_), .A2(new_n682_), .A3(KEYINPUT111), .A4(new_n703_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n659_), .B2(new_n560_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT47), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n706_), .A2(new_n711_), .A3(new_n707_), .A4(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1330gat));
  OR3_X1    g512(.A1(new_n659_), .A2(G50gat), .A3(new_n464_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n683_), .A2(new_n715_), .A3(new_n463_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G50gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n683_), .B2(new_n463_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1331gat));
  NAND4_X1  g518(.A1(new_n623_), .A2(new_n625_), .A3(new_n586_), .A4(new_n613_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(new_n317_), .A3(new_n531_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n616_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n586_), .A2(new_n608_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n561_), .A2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n344_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n726_), .B2(new_n725_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n721_), .B1(new_n728_), .B2(new_n317_), .ZN(G1332gat));
  OAI21_X1  g528(.A(G64gat), .B1(new_n720_), .B2(new_n688_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT48), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n725_), .A2(new_n315_), .A3(new_n689_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1333gat));
  OAI21_X1  g532(.A(G71gat), .B1(new_n720_), .B2(new_n560_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT49), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n725_), .A2(new_n482_), .A3(new_n649_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1334gat));
  OAI21_X1  g536(.A(G78gat), .B1(new_n720_), .B2(new_n464_), .ZN(new_n738_));
  XOR2_X1   g537(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n725_), .A2(new_n444_), .A3(new_n463_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1335gat));
  NAND3_X1  g541(.A1(new_n586_), .A2(new_n342_), .A3(new_n608_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n680_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n531_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n724_), .A2(new_n658_), .ZN(new_n747_));
  OR3_X1    g546(.A1(new_n747_), .A2(G85gat), .A3(new_n722_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1336gat));
  OAI21_X1  g548(.A(G92gat), .B1(new_n745_), .B2(new_n688_), .ZN(new_n750_));
  INV_X1    g549(.A(G92gat), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n636_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n747_), .B2(new_n752_), .ZN(G1337gat));
  OAI21_X1  g552(.A(G99gat), .B1(new_n745_), .B2(new_n560_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n560_), .A2(new_n211_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n747_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g556(.A1(new_n680_), .A2(new_n463_), .A3(new_n744_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n680_), .A2(KEYINPUT116), .A3(new_n463_), .A4(new_n744_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n760_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n761_), .ZN(new_n762_));
  AND4_X1   g561(.A1(new_n245_), .A2(new_n724_), .A3(new_n463_), .A4(new_n658_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n761_), .A2(G106gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(new_n767_), .B2(new_n760_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT53), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n760_), .A2(G106gat), .A3(new_n761_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n762_), .A4(new_n765_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n769_), .A2(new_n774_), .ZN(G1339gat));
  AND2_X1   g574(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n776_));
  NOR4_X1   g575(.A1(new_n609_), .A2(new_n612_), .A3(new_n342_), .A4(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n673_), .A2(new_n624_), .A3(new_n777_), .A4(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n624_), .A2(new_n777_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n303_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n626_), .A2(new_n581_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n570_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n571_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n566_), .A2(new_n569_), .A3(KEYINPUT55), .A4(new_n570_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n578_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n578_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n784_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n590_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n601_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n596_), .A2(new_n592_), .A3(new_n588_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n610_), .A2(new_n795_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n795_), .B1(new_n610_), .B2(new_n799_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n582_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n299_), .B1(new_n794_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n578_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n791_), .B(new_n580_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n581_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n807_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n811_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(KEYINPUT58), .C1(new_n808_), .C2(new_n809_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(new_n303_), .A3(new_n814_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n626_), .A2(new_n581_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n802_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(KEYINPUT57), .A3(new_n299_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n806_), .A2(new_n815_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n783_), .B1(new_n820_), .B2(new_n342_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n722_), .A2(new_n560_), .A3(new_n477_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(KEYINPUT120), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n821_), .A2(new_n823_), .A3(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n824_), .A2(KEYINPUT120), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n821_), .A2(new_n823_), .B1(new_n827_), .B2(new_n825_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G113gat), .B1(new_n829_), .B2(new_n613_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT57), .B1(new_n818_), .B2(new_n299_), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n805_), .B(new_n622_), .C1(new_n817_), .C2(new_n802_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n625_), .B1(new_n835_), .B2(new_n815_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT119), .B(new_n822_), .C1(new_n836_), .C2(new_n783_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n608_), .A2(G113gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n832_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n830_), .A2(new_n839_), .ZN(G1340gat));
  OAI21_X1  g639(.A(G120gat), .B1(new_n829_), .B2(new_n624_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT60), .ZN(new_n842_));
  AOI21_X1  g641(.A(G120gat), .B1(new_n586_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(G120gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(KEYINPUT121), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(KEYINPUT121), .B2(new_n843_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n832_), .A2(new_n837_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n841_), .A2(new_n847_), .ZN(G1341gat));
  OAI21_X1  g647(.A(G127gat), .B1(new_n829_), .B2(new_n342_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n342_), .A2(G127gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n832_), .A2(new_n837_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1342gat));
  AND4_X1   g651(.A1(G134gat), .A2(new_n826_), .A3(new_n303_), .A4(new_n828_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n832_), .A2(new_n837_), .A3(new_n622_), .ZN(new_n854_));
  INV_X1    g653(.A(G134gat), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT122), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n854_), .A2(new_n858_), .A3(new_n855_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n853_), .B1(new_n857_), .B2(new_n859_), .ZN(G1343gat));
  INV_X1    g659(.A(new_n821_), .ZN(new_n861_));
  NOR4_X1   g660(.A1(new_n689_), .A2(new_n464_), .A3(new_n649_), .A4(new_n722_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n608_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT123), .B(G141gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n863_), .A2(new_n624_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g667(.A1(new_n863_), .A2(new_n342_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n869_), .B(new_n870_), .Z(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n863_), .B2(new_n673_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n299_), .A2(G162gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n863_), .B2(new_n873_), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n616_), .A2(new_n560_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n689_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT124), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n689_), .A2(new_n878_), .A3(new_n875_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n877_), .A2(new_n464_), .A3(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n821_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n626_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G169gat), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n882_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n886_));
  INV_X1    g685(.A(new_n399_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n885_), .B(new_n886_), .C1(new_n887_), .C2(new_n882_), .ZN(G1348gat));
  NAND2_X1  g687(.A1(new_n881_), .A2(new_n586_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g689(.A(G183gat), .B1(new_n881_), .B2(new_n625_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n881_), .A2(new_n625_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n892_), .B(new_n893_), .C1(new_n405_), .C2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n405_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT125), .B1(new_n896_), .B2(new_n891_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1350gat));
  AND3_X1   g697(.A1(new_n881_), .A2(new_n622_), .A3(new_n370_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n352_), .B1(new_n881_), .B2(new_n303_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1351gat));
  NAND2_X1  g700(.A1(new_n560_), .A2(new_n557_), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT126), .Z(new_n903_));
  NOR3_X1   g702(.A1(new_n821_), .A2(new_n688_), .A3(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n626_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n586_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g707(.A(KEYINPUT63), .B(G211gat), .C1(new_n904_), .C2(new_n625_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n904_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n342_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT63), .B(G211gat), .Z(new_n912_));
  AOI21_X1  g711(.A(new_n909_), .B1(new_n911_), .B2(new_n912_), .ZN(G1354gat));
  AND3_X1   g712(.A1(new_n904_), .A2(G218gat), .A3(new_n303_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n904_), .A2(new_n622_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916_));
  AOI21_X1  g715(.A(G218gat), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT127), .B1(new_n910_), .B2(new_n299_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n914_), .B1(new_n917_), .B2(new_n918_), .ZN(G1355gat));
endmodule


