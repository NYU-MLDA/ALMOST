//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT86), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT85), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n203_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT83), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n210_), .A2(KEYINPUT84), .A3(KEYINPUT25), .A4(G183gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(KEYINPUT84), .A2(G183gat), .ZN(new_n212_));
  OAI221_X1 g011(.A(new_n211_), .B1(new_n210_), .B2(G183gat), .C1(KEYINPUT25), .C2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT26), .B(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT23), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n206_), .A2(new_n207_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n209_), .A2(new_n215_), .A3(new_n217_), .A4(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT22), .B(G169gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n203_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT83), .B(G183gat), .Z(new_n225_));
  OAI21_X1  g024(.A(new_n217_), .B1(G190gat), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G71gat), .B(G99gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G43gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n228_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT88), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT88), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT87), .B1(new_n234_), .B2(new_n235_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT87), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n238_), .B(new_n240_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G15gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT30), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n243_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n233_), .B(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n248_), .A2(KEYINPUT90), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(KEYINPUT90), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT18), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G64gat), .B(G92gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n254_), .B(new_n255_), .Z(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G226gat), .A2(G233gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT21), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G211gat), .B(G218gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G197gat), .B(G204gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT92), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n262_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G211gat), .B(G218gat), .Z(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n263_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n261_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(KEYINPUT92), .B2(new_n263_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n270_), .A2(KEYINPUT21), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT93), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n264_), .A2(new_n262_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT21), .B1(new_n270_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT93), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n266_), .A2(new_n261_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n272_), .A2(new_n277_), .A3(new_n227_), .A4(new_n221_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n217_), .B1(G183gat), .B2(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n224_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n208_), .B1(G169gat), .B2(G176gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT25), .B(G183gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n214_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n204_), .A2(new_n219_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n217_), .A3(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n281_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n269_), .A2(new_n271_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n279_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT97), .B1(new_n278_), .B2(KEYINPUT20), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n260_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n259_), .A2(KEYINPUT20), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n287_), .A2(new_n288_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT98), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n272_), .A2(new_n277_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n228_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n297_), .B(new_n299_), .C1(new_n296_), .C2(new_n295_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n256_), .B1(new_n292_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G29gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G85gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT0), .B(G57gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT3), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT2), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(KEYINPUT91), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT91), .B1(new_n312_), .B2(new_n314_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n310_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n309_), .B1(KEYINPUT1), .B2(new_n307_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n319_), .B1(KEYINPUT1), .B2(new_n307_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n311_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n313_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n234_), .A2(new_n235_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n237_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n318_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n310_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n312_), .A2(new_n314_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT91), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n326_), .B1(new_n329_), .B2(new_n315_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n322_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n325_), .B1(new_n332_), .B2(new_n243_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n306_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n243_), .B1(new_n318_), .B2(new_n322_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n318_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT4), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n318_), .A2(new_n322_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n243_), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT4), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n335_), .B1(new_n343_), .B2(new_n334_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n334_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n333_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n306_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n341_), .B1(new_n333_), .B2(KEYINPUT4), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n347_), .B(new_n348_), .C1(new_n349_), .C2(new_n334_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT33), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n344_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n292_), .A2(new_n300_), .A3(new_n256_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n334_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(new_n346_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(KEYINPUT33), .A3(new_n348_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n302_), .A2(new_n352_), .A3(new_n353_), .A4(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n306_), .B1(new_n354_), .B2(new_n346_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n350_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n256_), .A2(KEYINPUT32), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n292_), .A2(new_n300_), .A3(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n290_), .A2(new_n260_), .A3(new_n291_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n295_), .A2(KEYINPUT20), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n259_), .B1(new_n363_), .B2(new_n299_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n359_), .B(new_n361_), .C1(new_n365_), .C2(new_n360_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n357_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT29), .B1(new_n330_), .B2(new_n331_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n288_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n298_), .A2(new_n369_), .A3(new_n368_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT94), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n298_), .A2(new_n369_), .A3(KEYINPUT94), .A4(new_n368_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n370_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT95), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n339_), .A2(KEYINPUT29), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G22gat), .B(G50gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT28), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n379_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n375_), .A2(new_n377_), .ZN(new_n384_));
  AOI211_X1 g183(.A(new_n376_), .B(new_n370_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n385_));
  OAI22_X1  g184(.A1(new_n378_), .A2(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n373_), .A2(new_n374_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n370_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n376_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n375_), .A2(new_n377_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(KEYINPUT95), .A3(new_n391_), .A4(new_n382_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n386_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n367_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT99), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n359_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n397_));
  XOR2_X1   g196(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n398_));
  INV_X1    g197(.A(new_n353_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(new_n301_), .ZN(new_n400_));
  OAI211_X1 g199(.A(KEYINPUT27), .B(new_n353_), .C1(new_n365_), .C2(new_n256_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n395_), .A2(new_n396_), .B1(new_n397_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n393_), .B1(new_n366_), .B2(new_n357_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT99), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n252_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT101), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n401_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(new_n393_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n394_), .A2(KEYINPUT101), .A3(new_n400_), .A4(new_n401_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n359_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .A4(new_n248_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n406_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G29gat), .B(G36gat), .Z(new_n415_));
  XOR2_X1   g214(.A(G43gat), .B(G50gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT15), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G15gat), .B(G22gat), .ZN(new_n419_));
  INV_X1    g218(.A(G1gat), .ZN(new_n420_));
  INV_X1    g219(.A(G8gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT14), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT77), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n419_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n423_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G1gat), .B(G8gat), .ZN(new_n426_));
  OR3_X1    g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n418_), .A2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n427_), .A2(new_n428_), .A3(new_n417_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G229gat), .A2(G233gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n417_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n435_), .B1(new_n431_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G113gat), .B(G141gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G169gat), .B(G197gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n434_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(KEYINPUT81), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT81), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n438_), .A2(new_n446_), .A3(new_n442_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n448_), .B(KEYINPUT82), .Z(new_n449_));
  NOR2_X1   g248(.A1(new_n414_), .A2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(KEYINPUT10), .B(G99gat), .Z(new_n451_));
  INV_X1    g250(.A(G106gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT66), .B(G92gat), .ZN(new_n453_));
  INV_X1    g252(.A(G85gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(KEYINPUT9), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n451_), .A2(new_n452_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G99gat), .A2(G106gat), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G85gat), .A2(G92gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT9), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n456_), .A2(new_n461_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT67), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT69), .B(KEYINPUT7), .ZN(new_n470_));
  INV_X1    g269(.A(G99gat), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT68), .B1(new_n471_), .B2(new_n452_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n452_), .A3(KEYINPUT68), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n470_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n457_), .ZN(new_n476_));
  AND2_X1   g275(.A1(KEYINPUT71), .A2(KEYINPUT6), .ZN(new_n477_));
  NOR2_X1   g276(.A1(KEYINPUT71), .A2(KEYINPUT6), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT71), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n458_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(KEYINPUT71), .A2(KEYINPUT6), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n457_), .A3(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n479_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n465_), .B1(new_n475_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT72), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(KEYINPUT8), .ZN(new_n488_));
  AND2_X1   g287(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n489_));
  NOR2_X1   g288(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT68), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n492_), .A2(G99gat), .A3(G106gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n472_), .B2(new_n493_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n459_), .A2(new_n484_), .A3(new_n460_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n462_), .A2(new_n497_), .A3(new_n463_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT70), .ZN(new_n501_));
  AOI211_X1 g300(.A(KEYINPUT70), .B(new_n498_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n488_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n487_), .B1(new_n486_), .B2(KEYINPUT8), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n469_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n418_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n417_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n507_), .B(KEYINPUT76), .C1(new_n508_), .C2(new_n506_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G232gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  OR3_X1    g312(.A1(new_n509_), .A2(KEYINPUT75), .A3(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n513_), .B1(new_n509_), .B2(KEYINPUT75), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT35), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G190gat), .B(G218gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G134gat), .B(G162gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n509_), .A2(new_n516_), .B1(KEYINPUT36), .B2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n514_), .A2(new_n515_), .A3(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n519_), .A2(KEYINPUT36), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n514_), .A2(new_n524_), .A3(new_n515_), .A4(new_n520_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT37), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n429_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G57gat), .B(G64gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT11), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT73), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G71gat), .B(G78gat), .Z(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(KEYINPUT11), .B2(new_n531_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n534_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n530_), .B(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(G127gat), .B(G155gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G183gat), .B(G211gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT17), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n538_), .A2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT80), .Z(new_n546_));
  INV_X1    g345(.A(new_n538_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT78), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(KEYINPUT78), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n548_), .A2(KEYINPUT17), .A3(new_n543_), .A4(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n546_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n528_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n537_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n506_), .A2(new_n558_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n479_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n464_), .B1(new_n560_), .B2(new_n494_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT72), .B1(new_n561_), .B2(new_n497_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(new_n502_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n565_), .A3(new_n488_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(new_n537_), .A3(new_n469_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n559_), .A2(KEYINPUT12), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n537_), .B1(new_n566_), .B2(new_n469_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n557_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n556_), .B1(new_n559_), .B2(new_n567_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n578_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n580_), .A2(KEYINPUT74), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT74), .B1(new_n580_), .B2(new_n581_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT13), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n553_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n450_), .A2(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n587_), .A2(G1gat), .A3(new_n411_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT38), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT102), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n523_), .A2(new_n525_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n414_), .A2(new_n591_), .ZN(new_n592_));
  AND4_X1   g391(.A1(new_n448_), .A2(new_n592_), .A3(new_n551_), .A4(new_n585_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(new_n359_), .ZN(new_n594_));
  OAI221_X1 g393(.A(new_n590_), .B1(KEYINPUT38), .B2(new_n588_), .C1(new_n420_), .C2(new_n594_), .ZN(G1324gat));
  INV_X1    g394(.A(new_n587_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n421_), .A3(new_n408_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT39), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n408_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(G8gat), .ZN(new_n600_));
  AOI211_X1 g399(.A(KEYINPUT39), .B(new_n421_), .C1(new_n593_), .C2(new_n408_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT40), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(G1325gat));
  NAND2_X1  g403(.A1(new_n593_), .A2(new_n252_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G15gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n607_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n587_), .A2(G15gat), .A3(new_n251_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(G1326gat));
  INV_X1    g410(.A(G22gat), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n593_), .B2(new_n393_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT42), .Z(new_n614_));
  NAND3_X1  g413(.A1(new_n596_), .A2(new_n612_), .A3(new_n393_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1327gat));
  NAND3_X1  g415(.A1(new_n585_), .A2(new_n448_), .A3(new_n552_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n397_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n404_), .B2(KEYINPUT99), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n367_), .A2(KEYINPUT99), .A3(new_n394_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n251_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n412_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n619_), .B1(new_n624_), .B2(new_n528_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n526_), .B(KEYINPUT37), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT43), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(KEYINPUT104), .ZN(new_n628_));
  AOI211_X1 g427(.A(new_n626_), .B(new_n628_), .C1(new_n623_), .C2(new_n412_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n618_), .B1(new_n625_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n624_), .A2(new_n528_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n619_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n628_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n528_), .B(new_n637_), .C1(new_n406_), .C2(new_n413_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n617_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n633_), .B1(new_n639_), .B2(KEYINPUT44), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n630_), .A2(KEYINPUT105), .A3(new_n631_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n632_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G29gat), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n411_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n551_), .A2(new_n526_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n450_), .A2(new_n585_), .A3(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(new_n411_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n642_), .A2(new_n644_), .B1(new_n643_), .B2(new_n647_), .ZN(G1328gat));
  NOR3_X1   g447(.A1(new_n646_), .A2(G36gat), .A3(new_n402_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT45), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n642_), .A2(new_n408_), .ZN(new_n653_));
  INV_X1    g452(.A(G36gat), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n651_), .B(new_n652_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n652_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n654_), .B1(new_n642_), .B2(new_n408_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(new_n650_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(G1329gat));
  NAND2_X1  g458(.A1(new_n639_), .A2(KEYINPUT44), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n248_), .A2(G43gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n626_), .B1(new_n623_), .B2(new_n412_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n638_), .B1(new_n662_), .B2(new_n619_), .ZN(new_n663_));
  AOI211_X1 g462(.A(new_n633_), .B(KEYINPUT44), .C1(new_n663_), .C2(new_n618_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT105), .B1(new_n630_), .B2(new_n631_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n660_), .B(new_n661_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT107), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n640_), .A2(new_n641_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n660_), .A4(new_n661_), .ZN(new_n670_));
  INV_X1    g469(.A(G43gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n671_), .B1(new_n646_), .B2(new_n251_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n667_), .A2(new_n670_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT47), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT47), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n667_), .A2(new_n670_), .A3(new_n675_), .A4(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1330gat));
  INV_X1    g476(.A(G50gat), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n394_), .A2(new_n678_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n646_), .A2(new_n394_), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n642_), .A2(new_n679_), .B1(new_n678_), .B2(new_n680_), .ZN(G1331gat));
  INV_X1    g480(.A(new_n585_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(new_n449_), .A3(new_n551_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n592_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n411_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n448_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n624_), .A2(new_n686_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT108), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n585_), .B1(new_n687_), .B2(KEYINPUT108), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n553_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n411_), .A2(G57gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n685_), .B1(new_n691_), .B2(new_n692_), .ZN(G1332gat));
  OAI21_X1  g492(.A(G64gat), .B1(new_n684_), .B2(new_n402_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT48), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n402_), .A2(G64gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n691_), .B2(new_n696_), .ZN(G1333gat));
  OR2_X1    g496(.A1(new_n251_), .A2(G71gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n592_), .A2(new_n683_), .A3(new_n252_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(G71gat), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(G71gat), .ZN(new_n702_));
  OAI22_X1  g501(.A1(new_n691_), .A2(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT110), .ZN(G1334gat));
  OAI21_X1  g503(.A(G78gat), .B1(new_n684_), .B2(new_n394_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT50), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n394_), .A2(G78gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n691_), .B2(new_n707_), .ZN(G1335gat));
  NAND3_X1  g507(.A1(new_n688_), .A2(new_n645_), .A3(new_n689_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n454_), .A3(new_n359_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n585_), .A2(new_n448_), .A3(new_n551_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n663_), .A2(new_n712_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n713_), .A2(KEYINPUT111), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(KEYINPUT111), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n714_), .A2(KEYINPUT112), .A3(new_n715_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n411_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n711_), .B1(new_n720_), .B2(new_n454_), .ZN(G1336gat));
  AOI21_X1  g520(.A(G92gat), .B1(new_n710_), .B2(new_n408_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(new_n719_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n408_), .A2(new_n453_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(G1337gat));
  NAND3_X1  g524(.A1(new_n710_), .A2(new_n248_), .A3(new_n451_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n251_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(new_n471_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g528(.A1(new_n663_), .A2(new_n393_), .A3(new_n712_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(G106gat), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT52), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n394_), .A2(G106gat), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n690_), .A2(KEYINPUT113), .A3(new_n645_), .A4(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  INV_X1    g534(.A(new_n733_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n709_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n731_), .A2(KEYINPUT52), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n732_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g540(.A1(new_n553_), .A2(new_n585_), .A3(new_n449_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n742_), .B(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT56), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n566_), .A2(new_n537_), .A3(new_n469_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n571_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n556_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT55), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n572_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n568_), .A2(new_n557_), .A3(new_n571_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n568_), .A2(KEYINPUT116), .A3(new_n557_), .A4(new_n571_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n751_), .A2(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n746_), .B1(new_n758_), .B2(new_n579_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n579_), .A2(new_n746_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT118), .B1(new_n758_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n756_), .A2(new_n757_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n572_), .A2(new_n752_), .ZN(new_n764_));
  AOI211_X1 g563(.A(KEYINPUT55), .B(new_n557_), .C1(new_n568_), .C2(new_n571_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n760_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n759_), .A2(new_n762_), .A3(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n430_), .A2(new_n432_), .A3(new_n435_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n433_), .B1(new_n431_), .B2(new_n436_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n442_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n444_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n574_), .B2(new_n579_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n769_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT58), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT119), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n528_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT58), .B1(new_n769_), .B2(new_n774_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT119), .B1(new_n780_), .B2(new_n626_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n769_), .A2(KEYINPUT58), .A3(new_n774_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT120), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n779_), .A2(new_n781_), .A3(KEYINPUT120), .A4(new_n782_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT117), .B1(new_n758_), .B2(new_n761_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n766_), .A2(new_n788_), .A3(new_n760_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n759_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n580_), .A2(new_n448_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT115), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n773_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n584_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(KEYINPUT57), .A3(new_n526_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n790_), .A2(new_n792_), .B1(new_n584_), .B2(new_n794_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n591_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n797_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n785_), .A2(new_n786_), .A3(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n745_), .B1(new_n802_), .B2(new_n552_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n409_), .A2(new_n410_), .A3(new_n248_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(new_n359_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT59), .B1(new_n803_), .B2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n551_), .B1(new_n801_), .B2(new_n783_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n745_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811_), .B2(new_n449_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n797_), .A2(new_n800_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n551_), .B1(new_n814_), .B2(new_n786_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n805_), .B1(new_n815_), .B2(new_n745_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(G113gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n448_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n812_), .A2(new_n819_), .ZN(G1340gat));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  INV_X1    g620(.A(G120gat), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n810_), .A2(new_n682_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n807_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n585_), .B2(KEYINPUT60), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(KEYINPUT60), .B2(new_n822_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n816_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n821_), .B1(new_n824_), .B2(new_n827_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n816_), .A2(new_n826_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n810_), .A2(new_n682_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n816_), .B2(KEYINPUT59), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n829_), .B(KEYINPUT121), .C1(new_n831_), .C2(new_n822_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n832_), .ZN(G1341gat));
  OAI21_X1  g632(.A(G127gat), .B1(new_n811_), .B2(new_n552_), .ZN(new_n834_));
  INV_X1    g633(.A(G127gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n817_), .A2(new_n835_), .A3(new_n551_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1342gat));
  OAI21_X1  g636(.A(G134gat), .B1(new_n811_), .B2(new_n626_), .ZN(new_n838_));
  INV_X1    g637(.A(G134gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n817_), .A2(new_n839_), .A3(new_n591_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1343gat));
  INV_X1    g640(.A(new_n803_), .ZN(new_n842_));
  NOR4_X1   g641(.A1(new_n252_), .A2(new_n394_), .A3(new_n411_), .A4(new_n408_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n448_), .A3(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g644(.A1(new_n842_), .A2(new_n682_), .A3(new_n843_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g646(.A1(new_n842_), .A2(new_n551_), .A3(new_n843_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  OAI211_X1 g649(.A(new_n528_), .B(new_n843_), .C1(new_n815_), .C2(new_n745_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(G162gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n526_), .A2(G162gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n842_), .A2(new_n843_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT122), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n852_), .A2(new_n854_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1347gat));
  NOR3_X1   g658(.A1(new_n251_), .A2(new_n402_), .A3(new_n359_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n860_), .A2(new_n394_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n809_), .B2(new_n745_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT123), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n864_), .B(new_n861_), .C1(new_n809_), .C2(new_n745_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n223_), .A3(new_n448_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n862_), .A2(new_n686_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n868_), .A2(new_n869_), .A3(G169gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n868_), .B2(G169gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n867_), .B1(new_n870_), .B2(new_n871_), .ZN(G1348gat));
  NAND2_X1  g671(.A1(new_n866_), .A2(new_n682_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n222_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n585_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT124), .B1(new_n876_), .B2(G176gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT125), .B1(new_n803_), .B2(new_n393_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n879_), .B(new_n394_), .C1(new_n815_), .C2(new_n745_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n878_), .A2(new_n860_), .A3(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n585_), .A2(new_n222_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n875_), .A2(new_n877_), .B1(new_n881_), .B2(new_n882_), .ZN(G1349gat));
  NAND4_X1  g682(.A1(new_n878_), .A2(new_n551_), .A3(new_n880_), .A4(new_n860_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n225_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n552_), .A2(new_n283_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n884_), .A2(new_n885_), .B1(new_n866_), .B2(new_n886_), .ZN(G1350gat));
  NAND3_X1  g686(.A1(new_n866_), .A2(new_n214_), .A3(new_n591_), .ZN(new_n888_));
  INV_X1    g687(.A(G190gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n626_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(G1351gat));
  NAND2_X1  g690(.A1(new_n251_), .A2(new_n397_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n408_), .B1(new_n892_), .B2(KEYINPUT126), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(KEYINPUT126), .B2(new_n892_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n842_), .A2(new_n448_), .A3(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g695(.A1(new_n842_), .A2(new_n682_), .A3(new_n894_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n899_), .A2(KEYINPUT127), .ZN(new_n900_));
  XOR2_X1   g699(.A(new_n899_), .B(KEYINPUT127), .Z(new_n901_));
  AOI21_X1  g700(.A(new_n552_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n842_), .A2(new_n894_), .A3(new_n902_), .ZN(new_n903_));
  MUX2_X1   g702(.A(new_n900_), .B(new_n901_), .S(new_n903_), .Z(G1354gat));
  NAND2_X1  g703(.A1(new_n842_), .A2(new_n894_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G218gat), .B1(new_n905_), .B2(new_n626_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n526_), .A2(G218gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n905_), .B2(new_n907_), .ZN(G1355gat));
endmodule


