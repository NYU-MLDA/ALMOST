//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT22), .ZN(new_n208_));
  OAI21_X1  g007(.A(G169gat), .B1(new_n208_), .B2(KEYINPUT82), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT22), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT83), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(KEYINPUT83), .A3(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT23), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n221_), .A2(new_n223_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT84), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n218_), .A2(new_n219_), .A3(new_n230_), .A4(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n215_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OR3_X1    g035(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT25), .B(G183gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT26), .B(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT81), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n239_), .A2(new_n244_), .A3(new_n224_), .A4(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT21), .ZN(new_n247_));
  AND2_X1   g046(.A1(G197gat), .A2(G204gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G197gat), .A2(G204gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT91), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT91), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n252_), .B(new_n247_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n248_), .A2(new_n249_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT21), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n251_), .A2(new_n253_), .A3(new_n255_), .A4(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n255_), .A2(new_n256_), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n233_), .A2(new_n246_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n258_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n242_), .A2(new_n224_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n211_), .A2(KEYINPUT22), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n208_), .A2(G169gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(new_n213_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n215_), .ZN(new_n265_));
  OAI22_X1  g064(.A1(new_n261_), .A2(new_n238_), .B1(new_n231_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT20), .B1(new_n260_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT19), .ZN(new_n269_));
  NOR3_X1   g068(.A1(new_n259_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n257_), .A2(new_n258_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(new_n233_), .A3(new_n246_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n260_), .B2(new_n266_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n271_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n207_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n275_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n269_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n233_), .A2(new_n246_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n260_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n266_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n274_), .B1(new_n282_), .B2(new_n272_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n283_), .A3(new_n271_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n207_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n279_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT94), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n277_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT27), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n279_), .A2(new_n284_), .A3(KEYINPUT94), .A4(new_n285_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n269_), .B1(new_n259_), .B2(new_n267_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n269_), .B2(new_n278_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n293_), .B2(new_n207_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n286_), .A2(KEYINPUT100), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT100), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n279_), .A2(new_n284_), .A3(new_n296_), .A4(new_n285_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n291_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G141gat), .ZN(new_n301_));
  INV_X1    g100(.A(G148gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(KEYINPUT1), .B2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(KEYINPUT1), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n305_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OR3_X1    g112(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(KEYINPUT89), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n304_), .A2(KEYINPUT89), .A3(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n313_), .B(new_n314_), .C1(new_n316_), .C2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n307_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n320_), .A2(new_n306_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n310_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G22gat), .B(G50gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT28), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n324_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT90), .B1(new_n322_), .B2(new_n323_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT90), .ZN(new_n331_));
  INV_X1    g130(.A(new_n321_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n314_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n315_), .B(KEYINPUT89), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n331_), .B(KEYINPUT29), .C1(new_n335_), .C2(new_n310_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n330_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n260_), .B1(new_n322_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n338_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n329_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT93), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n327_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n340_), .A2(new_n344_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n328_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n340_), .A2(new_n344_), .A3(new_n329_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n349_), .A2(new_n346_), .A3(new_n350_), .A4(new_n327_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n300_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n316_), .A2(new_n318_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n314_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n321_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n310_), .ZN(new_n361_));
  INV_X1    g160(.A(G127gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n362_), .A2(G134gat), .ZN(new_n363_));
  INV_X1    g162(.A(G134gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n364_), .A2(G127gat), .ZN(new_n365_));
  INV_X1    g164(.A(G113gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n366_), .A2(G120gat), .ZN(new_n367_));
  INV_X1    g166(.A(G120gat), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n368_), .A2(G113gat), .ZN(new_n369_));
  OAI22_X1  g168(.A1(new_n363_), .A2(new_n365_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G127gat), .B(G134gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G113gat), .B(G120gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n373_), .A3(KEYINPUT86), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n360_), .A2(new_n361_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n357_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n370_), .A2(new_n373_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n360_), .A2(new_n361_), .A3(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n374_), .A2(new_n376_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n381_), .B(KEYINPUT4), .C1(new_n382_), .C2(new_n322_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n360_), .A2(new_n361_), .A3(new_n380_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(new_n377_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n357_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G1gat), .B(G29gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G85gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT0), .B(G57gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n389_), .B(new_n390_), .Z(new_n391_));
  AND3_X1   g190(.A1(new_n384_), .A2(new_n387_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(G71gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(G99gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n280_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G15gat), .B(G43gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT85), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT30), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n400_), .B(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n382_), .B(KEYINPUT31), .Z(new_n405_));
  INV_X1    g204(.A(KEYINPUT87), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(KEYINPUT88), .A3(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n400_), .A2(new_n403_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n400_), .A2(new_n403_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n405_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT88), .B1(new_n404_), .B2(new_n407_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n395_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n356_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n205_), .A2(KEYINPUT32), .A3(new_n206_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n293_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT99), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT99), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n293_), .A2(new_n420_), .A3(new_n417_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n416_), .B(KEYINPUT98), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n279_), .A3(new_n284_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n394_), .A2(new_n419_), .A3(new_n421_), .A4(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n383_), .A2(new_n379_), .B1(new_n386_), .B2(new_n357_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n391_), .ZN(new_n428_));
  AND4_X1   g227(.A1(new_n391_), .A2(new_n384_), .A3(new_n387_), .A4(new_n426_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT97), .ZN(new_n431_));
  INV_X1    g230(.A(new_n357_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n383_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT96), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n383_), .A3(KEYINPUT96), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n391_), .B1(new_n386_), .B2(new_n432_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n431_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n433_), .A2(KEYINPUT96), .A3(new_n383_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT96), .B1(new_n433_), .B2(new_n383_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n431_), .B(new_n439_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n430_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n288_), .A2(new_n290_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n424_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n355_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n394_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n449_), .A2(KEYINPUT101), .A3(new_n291_), .A4(new_n298_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n395_), .A2(new_n291_), .A3(new_n354_), .A4(new_n298_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT101), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n448_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n412_), .A2(new_n413_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n415_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(G99gat), .B2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(G99gat), .ZN(new_n459_));
  INV_X1    g258(.A(G106gat), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n459_), .B(new_n460_), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n464_), .A2(new_n466_), .A3(KEYINPUT66), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT66), .B1(new_n464_), .B2(new_n466_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n462_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT68), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G85gat), .A2(G92gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(G85gat), .A2(G92gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT68), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT8), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n473_), .A2(new_n476_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n458_), .A2(new_n461_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT8), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n468_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n464_), .A2(new_n466_), .A3(KEYINPUT66), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT10), .B(G99gat), .Z(new_n485_));
  AOI22_X1  g284(.A1(new_n483_), .A2(new_n484_), .B1(new_n460_), .B2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n475_), .B1(new_n474_), .B2(KEYINPUT9), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT65), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n489_), .B2(new_n472_), .ZN(new_n490_));
  AND2_X1   g289(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n491_));
  NOR2_X1   g290(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n488_), .B(new_n472_), .C1(new_n491_), .C2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n487_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n486_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n482_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G36gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G29gat), .ZN(new_n499_));
  INV_X1    g298(.A(G29gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G36gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G50gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G43gat), .ZN(new_n504_));
  INV_X1    g303(.A(G43gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G50gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n499_), .A2(new_n501_), .A3(new_n504_), .A4(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT15), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n497_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT34), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n478_), .A2(new_n481_), .B1(new_n486_), .B2(new_n495_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n510_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n512_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(KEYINPUT35), .A3(new_n514_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n512_), .A2(new_n520_), .A3(new_n517_), .A4(new_n515_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n521_), .A3(KEYINPUT74), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G190gat), .B(G218gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(KEYINPUT36), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n522_), .A2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n519_), .A2(new_n521_), .A3(KEYINPUT74), .A4(new_n526_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n525_), .A2(KEYINPUT36), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n456_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT103), .ZN(new_n536_));
  AND2_X1   g335(.A1(G230gat), .A2(G233gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT70), .ZN(new_n538_));
  AND2_X1   g337(.A1(G71gat), .A2(G78gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G57gat), .B(G64gat), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(KEYINPUT11), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT69), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n542_), .B2(KEYINPUT11), .ZN(new_n545_));
  INV_X1    g344(.A(G64gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(G57gat), .ZN(new_n547_));
  INV_X1    g346(.A(G57gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(G64gat), .ZN(new_n549_));
  AND4_X1   g348(.A1(new_n544_), .A2(new_n547_), .A3(new_n549_), .A4(KEYINPUT11), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n543_), .B1(new_n545_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n549_), .A3(KEYINPUT11), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT69), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n549_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT11), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n547_), .A2(new_n549_), .A3(new_n544_), .A4(KEYINPUT11), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n553_), .A2(new_n556_), .A3(new_n541_), .A4(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n551_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n538_), .B1(new_n497_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n516_), .A2(KEYINPUT70), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n516_), .A2(new_n561_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n537_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n551_), .A2(new_n558_), .A3(KEYINPUT71), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT71), .B1(new_n551_), .B2(new_n558_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT12), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT72), .B1(new_n568_), .B2(new_n516_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n516_), .B2(new_n561_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT71), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n559_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n551_), .A2(new_n558_), .A3(KEYINPUT71), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT72), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n575_), .A2(new_n497_), .A3(new_n576_), .A4(KEYINPUT12), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n537_), .B1(new_n516_), .B2(new_n561_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n569_), .A2(new_n571_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n565_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G120gat), .B(G148gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n565_), .A2(new_n579_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT13), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G1gat), .A2(G8gat), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(KEYINPUT75), .A3(KEYINPUT14), .ZN(new_n592_));
  INV_X1    g391(.A(G15gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(G22gat), .ZN(new_n594_));
  INV_X1    g393(.A(G22gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(G15gat), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT75), .B1(new_n591_), .B2(KEYINPUT14), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT76), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n598_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT76), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G15gat), .B(G22gat), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .A4(new_n592_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G1gat), .B(G8gat), .Z(new_n604_));
  AND3_X1   g403(.A1(new_n599_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n599_), .B2(new_n603_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n575_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT17), .ZN(new_n612_));
  XOR2_X1   g411(.A(G127gat), .B(G155gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT16), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n611_), .A2(new_n612_), .A3(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n616_), .B(KEYINPUT17), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n609_), .A2(new_n561_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n609_), .A2(new_n561_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n618_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G229gat), .A2(G233gat), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n599_), .A2(new_n603_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n604_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n599_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT77), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT77), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n510_), .A2(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .A4(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n631_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n634_), .A2(new_n636_), .A3(KEYINPUT78), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT78), .B1(new_n634_), .B2(new_n636_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n626_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n607_), .A2(new_n511_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n636_), .A3(new_n625_), .ZN(new_n641_));
  XOR2_X1   g440(.A(G113gat), .B(G141gat), .Z(new_n642_));
  XNOR2_X1  g441(.A(G169gat), .B(G197gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n639_), .A2(new_n641_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n590_), .A2(new_n624_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n536_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT104), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(KEYINPUT104), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n395_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n456_), .A2(new_n650_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n534_), .A2(KEYINPUT37), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n532_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT37), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n660_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n624_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n590_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n659_), .A2(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n394_), .B(KEYINPUT102), .Z(new_n669_));
  NOR3_X1   g468(.A1(new_n668_), .A2(G1gat), .A3(new_n669_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n670_), .A2(KEYINPUT38), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(KEYINPUT38), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n658_), .A2(new_n671_), .A3(new_n672_), .ZN(G1324gat));
  OR3_X1    g472(.A1(new_n668_), .A2(G8gat), .A3(new_n300_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n536_), .A2(new_n299_), .A3(new_n653_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G8gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT105), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT39), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n679_), .A3(G8gat), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n677_), .A2(new_n678_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n677_), .B2(new_n680_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n674_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(KEYINPUT40), .B(new_n674_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  OAI21_X1  g486(.A(G15gat), .B1(new_n657_), .B2(new_n455_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n690_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n668_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n455_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n593_), .A3(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n691_), .A2(new_n692_), .A3(new_n695_), .ZN(G1326gat));
  NAND3_X1  g495(.A1(new_n693_), .A2(new_n595_), .A3(new_n354_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n354_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(G22gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G22gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1327gat));
  NAND2_X1  g501(.A1(new_n623_), .A2(new_n534_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT108), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n659_), .A2(new_n590_), .A3(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT109), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(KEYINPUT109), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(new_n500_), .A3(new_n394_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n711_));
  INV_X1    g510(.A(new_n664_), .ZN(new_n712_));
  AOI22_X1  g511(.A1(new_n447_), .A2(new_n355_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n694_), .B1(new_n713_), .B2(new_n450_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n711_), .B(new_n712_), .C1(new_n714_), .C2(new_n415_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT107), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n454_), .A2(new_n455_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n415_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n711_), .A4(new_n712_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT43), .B1(new_n456_), .B2(new_n664_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n716_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n666_), .A2(new_n624_), .A3(new_n650_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(KEYINPUT44), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT44), .B1(new_n723_), .B2(new_n724_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n669_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n710_), .B1(new_n728_), .B2(new_n500_), .ZN(G1328gat));
  NAND4_X1  g528(.A1(new_n706_), .A2(new_n498_), .A3(new_n299_), .A4(new_n707_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT45), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n726_), .A2(new_n727_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT110), .B1(new_n732_), .B2(new_n299_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n723_), .A2(new_n724_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n736_), .A2(KEYINPUT110), .A3(new_n299_), .A4(new_n725_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G36gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n731_), .B1(new_n733_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT111), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n740_), .A2(KEYINPUT111), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n736_), .A2(new_n299_), .A3(new_n725_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(G36gat), .A3(new_n737_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n747_), .A2(KEYINPUT111), .A3(new_n740_), .A4(new_n731_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n743_), .A2(new_n748_), .ZN(G1329gat));
  NAND3_X1  g548(.A1(new_n732_), .A2(G43gat), .A3(new_n694_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n505_), .B1(new_n708_), .B2(new_n455_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g552(.A1(new_n709_), .A2(new_n503_), .A3(new_n354_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n732_), .A2(KEYINPUT112), .A3(new_n354_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(G50gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT112), .B1(new_n732_), .B2(new_n354_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n756_), .B2(new_n757_), .ZN(G1331gat));
  NOR4_X1   g557(.A1(new_n456_), .A2(new_n665_), .A3(new_n651_), .A4(new_n590_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n669_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n548_), .A3(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n590_), .A2(new_n651_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n536_), .A2(new_n624_), .A3(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n763_), .A2(new_n394_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n764_), .B2(new_n548_), .ZN(G1332gat));
  AOI21_X1  g564(.A(new_n546_), .B1(new_n763_), .B2(new_n299_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT48), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n759_), .A2(new_n546_), .A3(new_n299_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1333gat));
  AOI21_X1  g568(.A(new_n397_), .B1(new_n763_), .B2(new_n694_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT49), .Z(new_n771_));
  NAND3_X1  g570(.A1(new_n759_), .A2(new_n397_), .A3(new_n694_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1334gat));
  INV_X1    g572(.A(G78gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n763_), .B2(new_n354_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT50), .Z(new_n776_));
  NAND3_X1  g575(.A1(new_n759_), .A2(new_n774_), .A3(new_n354_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1335gat));
  NAND2_X1  g577(.A1(new_n762_), .A2(new_n623_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT113), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n723_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n395_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n456_), .A2(new_n651_), .A3(new_n590_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n704_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n669_), .A2(G85gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n782_), .B1(new_n784_), .B2(new_n785_), .ZN(G1336gat));
  OAI21_X1  g585(.A(G92gat), .B1(new_n781_), .B2(new_n300_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n300_), .A2(G92gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n784_), .B2(new_n788_), .ZN(G1337gat));
  INV_X1    g588(.A(new_n784_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(new_n694_), .A3(new_n485_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT115), .Z(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n723_), .A2(new_n694_), .A3(new_n780_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(G99gat), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(new_n793_), .A3(G99gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g597(.A1(new_n790_), .A2(new_n460_), .A3(new_n354_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n723_), .A2(KEYINPUT116), .A3(new_n354_), .A4(new_n780_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(G106gat), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n781_), .B2(new_n355_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n801_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n802_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n799_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n625_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n636_), .A2(new_n626_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n646_), .B1(new_n811_), .B2(new_n640_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n647_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n647_), .A2(KEYINPUT118), .A3(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n589_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n588_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n569_), .A2(new_n571_), .A3(new_n577_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n537_), .B1(new_n821_), .B2(new_n563_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT12), .B1(new_n497_), .B2(new_n559_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n568_), .A2(new_n516_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n576_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n825_), .A2(KEYINPUT55), .A3(new_n569_), .A4(new_n578_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n579_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n822_), .A2(new_n826_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n585_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n820_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n819_), .B1(new_n834_), .B2(KEYINPUT117), .ZN(new_n835_));
  INV_X1    g634(.A(new_n820_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n833_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n829_), .B2(new_n585_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n836_), .B(KEYINPUT117), .C1(new_n837_), .C2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n661_), .B1(new_n835_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n838_), .B1(new_n842_), .B2(new_n833_), .ZN(new_n843_));
  AOI211_X1 g642(.A(KEYINPUT120), .B(KEYINPUT56), .C1(new_n829_), .C2(new_n585_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT119), .B1(new_n818_), .B2(new_n588_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n647_), .A2(KEYINPUT118), .A3(new_n813_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT118), .B1(new_n647_), .B2(new_n813_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT119), .B(new_n588_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  OAI22_X1  g648(.A1(new_n843_), .A2(new_n844_), .B1(new_n845_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n664_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n588_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n848_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n851_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n856_), .B(new_n857_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n809_), .A2(new_n841_), .B1(new_n852_), .B2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT57), .B(new_n661_), .C1(new_n835_), .C2(new_n840_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n624_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n664_), .A2(new_n590_), .A3(new_n624_), .A4(new_n650_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT122), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n841_), .A2(new_n809_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n850_), .A2(new_n851_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n712_), .A3(new_n858_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n860_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n623_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871_));
  INV_X1    g670(.A(new_n864_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n865_), .A2(new_n873_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n356_), .A2(new_n669_), .A3(new_n455_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G113gat), .B1(new_n877_), .B2(new_n651_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n861_), .A2(new_n864_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n875_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n879_), .A2(KEYINPUT59), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n876_), .B2(KEYINPUT59), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n650_), .A2(new_n366_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT123), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n878_), .B1(new_n882_), .B2(new_n884_), .ZN(G1340gat));
  OAI21_X1  g684(.A(new_n368_), .B1(new_n590_), .B2(KEYINPUT60), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n877_), .B(new_n886_), .C1(KEYINPUT60), .C2(new_n368_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n882_), .A2(new_n666_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n368_), .ZN(G1341gat));
  NAND3_X1  g688(.A1(new_n877_), .A2(new_n362_), .A3(new_n624_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n882_), .A2(new_n624_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n362_), .ZN(G1342gat));
  NAND3_X1  g691(.A1(new_n877_), .A2(new_n364_), .A3(new_n534_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n882_), .A2(new_n712_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n364_), .ZN(G1343gat));
  AOI21_X1  g694(.A(new_n694_), .B1(new_n865_), .B2(new_n873_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n669_), .A2(new_n299_), .A3(new_n355_), .ZN(new_n897_));
  AOI21_X1  g696(.A(KEYINPUT124), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n871_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n899_));
  AOI211_X1 g698(.A(KEYINPUT122), .B(new_n864_), .C1(new_n869_), .C2(new_n623_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n455_), .B(new_n897_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n651_), .B1(new_n898_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G141gat), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n301_), .B(new_n651_), .C1(new_n898_), .C2(new_n903_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1344gat));
  OAI21_X1  g706(.A(new_n666_), .B1(new_n898_), .B2(new_n903_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G148gat), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n302_), .B(new_n666_), .C1(new_n898_), .C2(new_n903_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1345gat));
  OAI21_X1  g710(.A(new_n624_), .B1(new_n898_), .B2(new_n903_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT61), .B(G155gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n913_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n624_), .B(new_n915_), .C1(new_n898_), .C2(new_n903_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1346gat));
  INV_X1    g716(.A(G162gat), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n918_), .B(new_n534_), .C1(new_n898_), .C2(new_n903_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n896_), .A2(KEYINPUT124), .A3(new_n897_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n901_), .A2(new_n902_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n664_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n919_), .B1(new_n922_), .B2(new_n918_), .ZN(G1347gat));
  NOR3_X1   g722(.A1(new_n760_), .A2(new_n455_), .A3(new_n300_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n879_), .A2(new_n354_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT125), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n926_), .A2(KEYINPUT125), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n651_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n926_), .A2(new_n651_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(G169gat), .ZN(new_n934_));
  AOI211_X1 g733(.A(KEYINPUT62), .B(new_n211_), .C1(new_n926_), .C2(new_n651_), .ZN(new_n935_));
  OAI22_X1  g734(.A1(new_n930_), .A2(new_n931_), .B1(new_n934_), .B2(new_n935_), .ZN(G1348gat));
  OAI21_X1  g735(.A(new_n666_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n354_), .B1(new_n865_), .B2(new_n873_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n925_), .A2(new_n590_), .A3(new_n213_), .ZN(new_n939_));
  AOI22_X1  g738(.A1(new_n937_), .A2(new_n213_), .B1(new_n938_), .B2(new_n939_), .ZN(G1349gat));
  OR2_X1    g739(.A1(new_n926_), .A2(KEYINPUT125), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n927_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n623_), .A2(new_n240_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n938_), .A2(new_n624_), .A3(new_n924_), .ZN(new_n944_));
  AOI22_X1  g743(.A1(new_n942_), .A2(new_n943_), .B1(new_n225_), .B2(new_n944_), .ZN(G1350gat));
  AOI21_X1  g744(.A(new_n664_), .B1(new_n941_), .B2(new_n927_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n534_), .A2(new_n241_), .ZN(new_n947_));
  OAI22_X1  g746(.A1(new_n946_), .A2(new_n226_), .B1(new_n930_), .B2(new_n947_), .ZN(G1351gat));
  AND2_X1   g747(.A1(new_n299_), .A2(new_n449_), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n455_), .B(new_n949_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n950_), .A2(new_n650_), .ZN(new_n951_));
  XOR2_X1   g750(.A(new_n951_), .B(G197gat), .Z(G1352gat));
  NAND3_X1  g751(.A1(new_n896_), .A2(new_n666_), .A3(new_n949_), .ZN(new_n953_));
  INV_X1    g752(.A(G204gat), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(KEYINPUT126), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n954_), .A2(KEYINPUT126), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n953_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n957_), .B1(new_n953_), .B2(new_n955_), .ZN(G1353gat));
  NAND3_X1  g757(.A1(new_n896_), .A2(new_n624_), .A3(new_n949_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  AND2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n959_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n962_), .B1(new_n959_), .B2(new_n960_), .ZN(G1354gat));
  OAI21_X1  g762(.A(G218gat), .B1(new_n950_), .B2(new_n664_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n661_), .A2(G218gat), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n896_), .A2(new_n949_), .A3(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n964_), .A2(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n967_), .A2(KEYINPUT127), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n964_), .A2(new_n969_), .A3(new_n966_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n970_), .ZN(G1355gat));
endmodule


