//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_;
  XNOR2_X1  g000(.A(KEYINPUT94), .B(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT81), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT24), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n206_), .B1(G169gat), .B2(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT26), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT25), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G183gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(G183gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(KEYINPUT26), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n208_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT82), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT23), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n218_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n220_), .B1(new_n224_), .B2(new_n219_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n204_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(KEYINPUT24), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT90), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT90), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n225_), .B(new_n229_), .C1(KEYINPUT24), .C2(new_n226_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n216_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G197gat), .B(G204gat), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G197gat), .B(G204gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT21), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G211gat), .B(G218gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n234_), .A2(new_n237_), .A3(new_n235_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G169gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n243_), .B1(new_n224_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OR3_X1    g045(.A1(new_n231_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT19), .ZN(new_n249_));
  INV_X1    g048(.A(new_n244_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n225_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n243_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT79), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n253_), .A2(new_n212_), .B1(new_n214_), .B2(KEYINPUT80), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(KEYINPUT80), .B2(new_n214_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n210_), .B(new_n213_), .C1(new_n253_), .C2(new_n212_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n208_), .B(new_n223_), .C1(KEYINPUT24), .C2(new_n205_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n252_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n249_), .B1(new_n259_), .B2(new_n241_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n247_), .A2(KEYINPUT20), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n249_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT20), .ZN(new_n263_));
  INV_X1    g062(.A(new_n259_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n240_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n241_), .B1(new_n231_), .B2(new_n246_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n262_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G8gat), .B(G36gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT18), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G64gat), .B(G92gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n261_), .A2(new_n267_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n267_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n247_), .A2(KEYINPUT20), .A3(new_n260_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n271_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n203_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT95), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n272_), .B1(new_n261_), .B2(new_n267_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(new_n271_), .A3(new_n275_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT95), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(new_n203_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT93), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n247_), .A2(new_n284_), .A3(KEYINPUT20), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n259_), .A2(new_n241_), .ZN(new_n286_));
  NOR3_X1   g085(.A1(new_n231_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT93), .B1(new_n287_), .B2(new_n263_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n289_), .A2(new_n249_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n265_), .A2(new_n266_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(new_n249_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n272_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n280_), .A2(KEYINPUT27), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n278_), .A2(new_n283_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G113gat), .B(G120gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT87), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n307_), .B(KEYINPUT3), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n309_), .B(KEYINPUT2), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n300_), .A2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n310_), .A2(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n298_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n298_), .B(KEYINPUT85), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(new_n317_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT4), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(KEYINPUT4), .B2(new_n319_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n321_), .B(KEYINPUT91), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n322_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G1gat), .B(G29gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G85gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT0), .B(G57gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n322_), .B(new_n333_), .C1(new_n326_), .C2(new_n328_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n240_), .B1(new_n315_), .B2(KEYINPUT29), .ZN(new_n338_));
  AND2_X1   g137(.A1(G228gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n338_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G22gat), .B(G50gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n317_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT28), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n315_), .A2(KEYINPUT29), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n344_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n338_), .A2(new_n340_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n338_), .A2(new_n340_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n342_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n353_), .A2(KEYINPUT88), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n347_), .A2(new_n350_), .A3(new_n344_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n343_), .A2(new_n352_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT88), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT89), .B1(new_n358_), .B2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n355_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n357_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n351_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n361_), .A4(new_n356_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n343_), .A2(new_n359_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(new_n365_), .B2(new_n351_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n337_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n271_), .A2(KEYINPUT32), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n274_), .A2(new_n373_), .A3(new_n275_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n337_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n292_), .B1(new_n289_), .B2(new_n249_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(new_n373_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n333_), .B1(new_n320_), .B2(new_n327_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n378_), .A2(KEYINPUT92), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n324_), .A2(KEYINPUT4), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n320_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n321_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(KEYINPUT92), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n379_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT33), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n336_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n327_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n388_), .A2(KEYINPUT33), .A3(new_n322_), .A4(new_n333_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  OAI22_X1  g189(.A1(new_n375_), .A2(new_n377_), .B1(new_n390_), .B2(new_n281_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n369_), .A2(new_n371_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n295_), .A2(new_n372_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n259_), .B(KEYINPUT30), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT86), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n395_), .A2(new_n396_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n394_), .A2(KEYINPUT84), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  INV_X1    g201(.A(G71gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G99gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G15gat), .B(G43gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT83), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n406_), .B(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n401_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n398_), .A2(new_n400_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n323_), .B(KEYINPUT31), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n410_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n412_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n398_), .A2(new_n400_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n410_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n413_), .B1(new_n419_), .B2(new_n411_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT96), .B1(new_n393_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n293_), .A2(new_n294_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n282_), .B1(new_n281_), .B2(new_n203_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n283_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n392_), .B(new_n423_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n337_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n372_), .B(new_n423_), .C1(new_n425_), .C2(new_n424_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n391_), .A2(new_n392_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT96), .ZN(new_n434_));
  INV_X1    g233(.A(new_n421_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n422_), .A2(new_n430_), .A3(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G15gat), .B(G22gat), .ZN(new_n438_));
  INV_X1    g237(.A(G1gat), .ZN(new_n439_));
  INV_X1    g238(.A(G8gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT14), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G1gat), .B(G8gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G29gat), .B(G36gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G43gat), .B(G50gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n444_), .B(new_n447_), .Z(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n447_), .B(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n444_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n454_), .B2(new_n447_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n451_), .B1(new_n449_), .B2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G113gat), .B(G141gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(G169gat), .B(G197gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n457_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G232gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT34), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT69), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G99gat), .A3(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT66), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n472_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT66), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n405_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(KEYINPUT67), .A3(new_n473_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n471_), .A2(new_n476_), .A3(new_n477_), .A4(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT68), .ZN(new_n483_));
  XOR2_X1   g282(.A(G85gat), .B(G92gat), .Z(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT8), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n483_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n464_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n482_), .A2(new_n484_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT68), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n490_), .A2(KEYINPUT69), .A3(KEYINPUT8), .A4(new_n485_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n469_), .A2(new_n480_), .A3(new_n473_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT65), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT8), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n484_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n488_), .A2(new_n491_), .A3(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(KEYINPUT10), .B(G99gat), .Z(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT64), .B(G106gat), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n484_), .A2(KEYINPUT9), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT9), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(G85gat), .A3(G92gat), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n501_), .A2(new_n502_), .A3(new_n504_), .A4(new_n469_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n498_), .A2(new_n505_), .A3(new_n447_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n453_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n508_));
  OAI211_X1 g307(.A(KEYINPUT35), .B(new_n463_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n463_), .A2(KEYINPUT35), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n463_), .A2(KEYINPUT35), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .A4(new_n506_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT72), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G190gat), .B(G218gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G134gat), .B(G162gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT36), .Z(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(new_n515_), .A3(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n518_), .A2(KEYINPUT36), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n509_), .A2(new_n513_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n515_), .B1(new_n514_), .B2(new_n519_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n514_), .A2(new_n519_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n522_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n525_), .A2(new_n526_), .B1(KEYINPUT37), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n530_), .A2(KEYINPUT70), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(KEYINPUT70), .ZN(new_n532_));
  OR3_X1    g331(.A1(new_n531_), .A2(new_n532_), .A3(KEYINPUT11), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT11), .B1(new_n531_), .B2(new_n532_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G71gat), .B(G78gat), .Z(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n534_), .A2(new_n535_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G231gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n536_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT74), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT74), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n444_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G127gat), .B(G155gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G183gat), .B(G211gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n543_), .A2(new_n546_), .A3(new_n454_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n548_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT76), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n548_), .A2(KEYINPUT76), .A3(new_n555_), .A4(new_n556_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n553_), .B(new_n554_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n548_), .B2(new_n556_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT77), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT77), .ZN(new_n566_));
  AOI211_X1 g365(.A(new_n566_), .B(new_n563_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n529_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT78), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT13), .ZN(new_n572_));
  INV_X1    g371(.A(G230gat), .ZN(new_n573_));
  INV_X1    g372(.A(G233gat), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n505_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n490_), .A2(KEYINPUT8), .A3(new_n485_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n496_), .B1(new_n577_), .B2(new_n464_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n576_), .B1(new_n578_), .B2(new_n491_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n536_), .A2(new_n537_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n575_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n498_), .A2(new_n505_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n580_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  AOI211_X1 g384(.A(KEYINPUT12), .B(new_n580_), .C1(new_n498_), .C2(new_n505_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n581_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n583_), .A2(new_n584_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n580_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n575_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G120gat), .B(G148gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT5), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(new_n590_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n587_), .B2(new_n590_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n572_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n598_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(KEYINPUT13), .A3(new_n596_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n570_), .A2(new_n571_), .A3(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n437_), .A2(new_n461_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n570_), .A2(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT78), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n439_), .A3(new_n337_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610_));
  OR3_X1    g409(.A1(new_n609_), .A2(KEYINPUT97), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n527_), .A2(KEYINPUT72), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n614_), .A2(KEYINPUT98), .A3(new_n522_), .A4(new_n520_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n421_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n429_), .B1(new_n617_), .B2(new_n434_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n616_), .B1(new_n618_), .B2(new_n422_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n561_), .A2(new_n564_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n461_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n602_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n439_), .B1(new_n623_), .B2(new_n337_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n609_), .B1(new_n610_), .B2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT97), .B1(new_n609_), .B2(new_n610_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n611_), .A2(new_n625_), .A3(new_n626_), .ZN(G1324gat));
  OAI21_X1  g426(.A(new_n423_), .B1(new_n425_), .B2(new_n424_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n616_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n437_), .A2(new_n628_), .A3(new_n629_), .A4(new_n622_), .ZN(new_n630_));
  XOR2_X1   g429(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n631_));
  AND3_X1   g430(.A1(new_n630_), .A2(G8gat), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n630_), .B2(G8gat), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n295_), .A2(G8gat), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n605_), .A2(new_n635_), .A3(new_n607_), .A4(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n621_), .B1(new_n618_), .B2(new_n422_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n638_), .A2(new_n607_), .A3(new_n604_), .A4(new_n636_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT99), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n634_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n634_), .B2(new_n641_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n643_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n634_), .A2(new_n641_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT102), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n634_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n645_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n647_), .A2(new_n651_), .ZN(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n623_), .B2(new_n421_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT41), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n608_), .A2(new_n653_), .A3(new_n421_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1326gat));
  INV_X1    g456(.A(new_n392_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n623_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G22gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT103), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n662_), .A3(G22gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(KEYINPUT42), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n608_), .A2(new_n665_), .A3(new_n658_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT42), .B1(new_n661_), .B2(new_n663_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1327gat));
  NAND3_X1  g468(.A1(new_n569_), .A2(new_n603_), .A3(new_n461_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT104), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n529_), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT43), .B(new_n673_), .C1(new_n618_), .C2(new_n422_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n437_), .B2(new_n529_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n672_), .B(KEYINPUT44), .C1(new_n674_), .C2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(G29gat), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n427_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n437_), .A2(new_n529_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT43), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n437_), .A2(new_n675_), .A3(new_n529_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n671_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n677_), .B(new_n679_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n629_), .A2(new_n568_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(new_n602_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n638_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n678_), .B1(new_n689_), .B2(new_n427_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n685_), .A2(new_n690_), .ZN(G1328gat));
  OR2_X1    g490(.A1(new_n628_), .A2(KEYINPUT106), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n628_), .A2(KEYINPUT106), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(G36gat), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT107), .B1(new_n689_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n638_), .A2(new_n688_), .A3(new_n699_), .A4(new_n696_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n698_), .A2(KEYINPUT45), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT45), .B1(new_n698_), .B2(new_n700_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n677_), .B(new_n628_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G36gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(new_n705_), .A3(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  OAI21_X1  g509(.A(new_n677_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n421_), .A2(G43gat), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n689_), .A2(new_n435_), .ZN(new_n713_));
  OAI22_X1  g512(.A1(new_n711_), .A2(new_n712_), .B1(G43gat), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g514(.A1(new_n689_), .A2(G50gat), .A3(new_n392_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n677_), .B(new_n658_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G50gat), .B1(new_n717_), .B2(new_n718_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1331gat));
  NAND2_X1  g520(.A1(new_n620_), .A2(new_n566_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n561_), .A2(KEYINPUT77), .A3(new_n564_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n621_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n603_), .A2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n619_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n427_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n461_), .B1(new_n618_), .B2(new_n422_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n729_), .A2(new_n602_), .A3(new_n570_), .ZN(new_n730_));
  INV_X1    g529(.A(G57gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n337_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n732_), .ZN(G1332gat));
  INV_X1    g532(.A(G64gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n726_), .B2(new_n694_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT48), .Z(new_n736_));
  NAND3_X1  g535(.A1(new_n730_), .A2(new_n734_), .A3(new_n694_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1333gat));
  AOI21_X1  g537(.A(new_n403_), .B1(new_n726_), .B2(new_n421_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT49), .Z(new_n740_));
  NAND2_X1  g539(.A1(new_n421_), .A2(new_n403_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT109), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n730_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(G1334gat));
  OAI21_X1  g543(.A(G78gat), .B1(new_n727_), .B2(new_n392_), .ZN(new_n745_));
  XOR2_X1   g544(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n392_), .A2(G78gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT111), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n730_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(G1335gat));
  NOR2_X1   g550(.A1(new_n687_), .A2(new_n603_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n729_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(G85gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(new_n337_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n603_), .A2(new_n568_), .A3(new_n461_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT112), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n757_), .C1(new_n674_), .C2(new_n676_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n427_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n756_), .B1(new_n762_), .B2(new_n755_), .ZN(G1336gat));
  INV_X1    g562(.A(G92gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n754_), .A2(new_n764_), .A3(new_n628_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n695_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n764_), .ZN(G1337gat));
  NAND2_X1  g566(.A1(new_n421_), .A2(new_n499_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n753_), .A2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT113), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n435_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n405_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT51), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n770_), .C1(new_n771_), .C2(new_n405_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n754_), .A2(new_n500_), .A3(new_n658_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n658_), .B(new_n757_), .C1(new_n674_), .C2(new_n676_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(G106gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G106gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n596_), .A2(KEYINPUT116), .A3(new_n461_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT116), .B1(new_n596_), .B2(new_n461_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI22_X1  g586(.A1(new_n585_), .A2(new_n586_), .B1(new_n584_), .B2(new_n583_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n575_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n587_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n581_), .B(KEYINPUT55), .C1(new_n585_), .C2(new_n586_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n594_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n793_), .B2(new_n594_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n787_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n456_), .A2(KEYINPUT117), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n456_), .A2(KEYINPUT117), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n450_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n460_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n457_), .A2(new_n460_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n600_), .B2(new_n596_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n616_), .B1(new_n796_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n784_), .B1(new_n806_), .B2(KEYINPUT57), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n793_), .A2(new_n594_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n594_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n804_), .B1(new_n813_), .B2(new_n787_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT118), .B(new_n808_), .C1(new_n814_), .C2(new_n616_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n806_), .A2(KEYINPUT57), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n597_), .A2(new_n803_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n813_), .A2(KEYINPUT58), .A3(new_n817_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n529_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n807_), .A2(new_n815_), .A3(new_n816_), .A4(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n620_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n724_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n568_), .A2(KEYINPUT114), .A3(new_n621_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n603_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n826_), .B1(new_n830_), .B2(new_n529_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT114), .B1(new_n568_), .B2(new_n621_), .ZN(new_n832_));
  NOR4_X1   g631(.A1(new_n565_), .A2(new_n567_), .A3(new_n827_), .A4(new_n461_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(new_n603_), .A3(new_n673_), .A4(new_n825_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n824_), .A2(new_n837_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n435_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n808_), .B1(new_n814_), .B2(new_n616_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n816_), .A3(new_n822_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n836_), .B1(new_n843_), .B2(new_n569_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n841_), .ZN(new_n845_));
  OAI22_X1  g644(.A1(new_n840_), .A2(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(G113gat), .B1(new_n846_), .B2(new_n621_), .ZN(new_n847_));
  INV_X1    g646(.A(G113gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n840_), .A2(new_n848_), .A3(new_n461_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1340gat));
  OAI21_X1  g649(.A(G120gat), .B1(new_n846_), .B2(new_n603_), .ZN(new_n851_));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n603_), .B2(KEYINPUT60), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n840_), .B(new_n853_), .C1(KEYINPUT60), .C2(new_n852_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n846_), .B2(new_n620_), .ZN(new_n856_));
  INV_X1    g655(.A(G127gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n840_), .A2(new_n857_), .A3(new_n568_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1342gat));
  OAI21_X1  g658(.A(G134gat), .B1(new_n846_), .B2(new_n673_), .ZN(new_n860_));
  INV_X1    g659(.A(G134gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n840_), .A2(new_n861_), .A3(new_n616_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1343gat));
  AOI21_X1  g662(.A(new_n836_), .B1(new_n823_), .B2(new_n620_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n695_), .A2(new_n435_), .A3(new_n658_), .A4(new_n337_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n461_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n602_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT119), .B(G148gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1345gat));
  OR2_X1    g670(.A1(new_n864_), .A2(new_n865_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT120), .B1(new_n872_), .B2(new_n569_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n866_), .A2(new_n874_), .A3(new_n568_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n873_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1346gat));
  OR3_X1    g678(.A1(new_n872_), .A2(G162gat), .A3(new_n629_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G162gat), .B1(new_n872_), .B2(new_n673_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1347gat));
  OR3_X1    g681(.A1(new_n695_), .A2(KEYINPUT121), .A3(new_n428_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT121), .B1(new_n695_), .B2(new_n428_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n392_), .A3(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n844_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT22), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n461_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n889_));
  INV_X1    g688(.A(G169gat), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n844_), .A2(new_n885_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n621_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n888_), .A2(KEYINPUT62), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n889_), .B1(new_n894_), .B2(new_n895_), .ZN(G1348gat));
  NOR2_X1   g695(.A1(new_n864_), .A2(new_n885_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n602_), .A2(G176gat), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n897_), .A2(KEYINPUT122), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT122), .B1(new_n897_), .B2(new_n898_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G176gat), .B1(new_n886_), .B2(new_n602_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(G1349gat));
  AOI21_X1  g701(.A(G183gat), .B1(new_n897_), .B2(new_n568_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n620_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n886_), .B2(new_n904_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n891_), .B2(new_n673_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n616_), .A2(new_n210_), .A3(new_n214_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n891_), .B2(new_n907_), .ZN(G1351gat));
  NOR2_X1   g707(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(KEYINPUT125), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n694_), .A2(new_n435_), .A3(new_n372_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n838_), .B2(new_n913_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n864_), .A2(KEYINPUT123), .A3(new_n912_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n461_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n910_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n838_), .A2(new_n911_), .A3(new_n913_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT123), .B1(new_n864_), .B2(new_n912_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n621_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n917_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n910_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n918_), .A2(new_n924_), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n919_), .A2(new_n920_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n603_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  OR2_X1    g727(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1353gat));
  INV_X1    g729(.A(new_n620_), .ZN(new_n931_));
  AOI211_X1 g730(.A(KEYINPUT63), .B(G211gat), .C1(new_n926_), .C2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n914_), .A2(new_n915_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT63), .B(G211gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n933_), .A2(new_n620_), .A3(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n932_), .A2(new_n935_), .ZN(G1354gat));
  OAI21_X1  g735(.A(G218gat), .B1(new_n933_), .B2(new_n673_), .ZN(new_n937_));
  INV_X1    g736(.A(G218gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n926_), .A2(new_n938_), .A3(new_n616_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(G1355gat));
endmodule


