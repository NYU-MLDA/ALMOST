//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G29gat), .B(G36gat), .Z(new_n204_));
  XOR2_X1   g003(.A(G43gat), .B(G50gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208_));
  INV_X1    g007(.A(G1gat), .ZN(new_n209_));
  INV_X1    g008(.A(G8gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G1gat), .B(G8gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n207_), .A2(new_n214_), .A3(KEYINPUT75), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT75), .B1(new_n207_), .B2(new_n214_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n206_), .B(KEYINPUT15), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n214_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n203_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n215_), .A2(new_n216_), .B1(new_n214_), .B2(new_n207_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n203_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G141gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G169gat), .B(G197gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n225_), .B(new_n226_), .Z(new_n227_));
  XNOR2_X1  g026(.A(new_n224_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT79), .B1(new_n229_), .B2(G190gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT26), .B(G190gat), .Z(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(KEYINPUT79), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT76), .B(G183gat), .Z(new_n233_));
  INV_X1    g032(.A(KEYINPUT77), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(KEYINPUT25), .ZN(new_n235_));
  INV_X1    g034(.A(G183gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n236_), .B1(KEYINPUT78), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(KEYINPUT78), .B2(new_n237_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT76), .B(G183gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT77), .B1(new_n240_), .B2(new_n237_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n232_), .A2(new_n235_), .A3(new_n239_), .A4(new_n241_), .ZN(new_n242_));
  OR3_X1    g041(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n243_));
  INV_X1    g042(.A(G169gat), .ZN(new_n244_));
  INV_X1    g043(.A(G176gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n243_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT23), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n249_), .B1(G183gat), .B2(G190gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(G183gat), .A3(G190gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n248_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(G169gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(KEYINPUT80), .A3(new_n252_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n252_), .A2(KEYINPUT80), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n250_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n240_), .A2(G190gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n256_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n254_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G71gat), .B(G99gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G43gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n263_), .B(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G227gat), .A2(G233gat), .ZN(new_n267_));
  INV_X1    g066(.A(G15gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT30), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n266_), .B(new_n270_), .Z(new_n271_));
  INV_X1    g070(.A(KEYINPUT81), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT84), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT82), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G127gat), .B(G134gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G113gat), .B(G120gat), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G113gat), .B(G120gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n276_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT82), .B1(new_n278_), .B2(new_n279_), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n283_), .A2(KEYINPUT83), .A3(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT83), .B1(new_n283_), .B2(new_n284_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT31), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n275_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(KEYINPUT84), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(KEYINPUT81), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n291_), .A2(new_n271_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293_));
  INV_X1    g092(.A(G141gat), .ZN(new_n294_));
  INV_X1    g093(.A(G148gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n296_), .A2(new_n298_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT87), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT87), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n301_), .A2(new_n308_), .A3(new_n305_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT86), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT85), .B1(new_n302_), .B2(KEYINPUT1), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n304_), .B1(new_n303_), .B2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n302_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G141gat), .B(G148gat), .Z(new_n318_));
  AOI21_X1  g117(.A(new_n311_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n304_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n316_), .B(new_n320_), .C1(KEYINPUT1), .C2(new_n302_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n311_), .B(new_n318_), .C1(new_n321_), .C2(new_n312_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n310_), .B1(new_n319_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n318_), .B1(new_n321_), .B2(new_n312_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT86), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n327_), .A2(new_n322_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n280_), .A2(new_n282_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT97), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n325_), .A2(KEYINPUT4), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n324_), .A2(new_n285_), .A3(new_n336_), .A4(new_n286_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n325_), .A2(new_n334_), .A3(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(G85gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT0), .B(G57gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n344_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n338_), .A2(new_n339_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n289_), .A2(new_n292_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n324_), .A2(KEYINPUT29), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G197gat), .B(G204gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT91), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G211gat), .B(G218gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(G197gat), .A2(G204gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G197gat), .A2(G204gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(KEYINPUT91), .A3(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n354_), .A2(new_n356_), .A3(KEYINPUT21), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n352_), .A2(KEYINPUT21), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT21), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n357_), .A2(new_n362_), .A3(new_n358_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n356_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n360_), .B1(new_n364_), .B2(KEYINPUT90), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT90), .ZN(new_n366_));
  AOI211_X1 g165(.A(new_n366_), .B(new_n356_), .C1(new_n361_), .C2(new_n363_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT92), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n363_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n362_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n355_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n366_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n364_), .A2(KEYINPUT90), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT92), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .A4(new_n360_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G228gat), .A2(G233gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n376_), .B(KEYINPUT89), .Z(new_n377_));
  NAND4_X1  g176(.A1(new_n351_), .A2(new_n368_), .A3(new_n375_), .A4(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n372_), .A2(new_n373_), .A3(new_n360_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n379_), .B1(new_n328_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT93), .ZN(new_n382_));
  INV_X1    g181(.A(new_n376_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n378_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(new_n378_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n328_), .A2(new_n380_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G22gat), .B(G50gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n391_), .B(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n388_), .A2(KEYINPUT94), .A3(new_n390_), .A4(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT94), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n390_), .A2(new_n398_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n399_), .A2(new_n395_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT19), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n263_), .B1(new_n368_), .B2(new_n375_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n365_), .A2(new_n367_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n257_), .A2(new_n259_), .ZN(new_n406_));
  XOR2_X1   g205(.A(KEYINPUT25), .B(G183gat), .Z(new_n407_));
  NOR2_X1   g206(.A1(new_n231_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(new_n248_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n251_), .A2(new_n252_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(G183gat), .B2(G190gat), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n406_), .A2(new_n409_), .B1(new_n411_), .B2(new_n256_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT20), .B1(new_n405_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n403_), .B1(new_n404_), .B2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G8gat), .B(G36gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n368_), .A2(new_n263_), .A3(new_n375_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n405_), .B2(new_n412_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n403_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n414_), .A2(new_n420_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n420_), .B1(new_n414_), .B2(new_n425_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n427_), .A2(new_n428_), .A3(KEYINPUT27), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n404_), .A2(new_n413_), .A3(new_n403_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n424_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n419_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT99), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT99), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n434_), .B(new_n419_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n426_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n429_), .B1(new_n436_), .B2(KEYINPUT27), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT100), .B1(new_n401_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n399_), .A2(new_n395_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n388_), .A2(new_n390_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n396_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n421_), .A2(new_n423_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n403_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n368_), .A2(new_n375_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n263_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n412_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n422_), .B1(new_n448_), .B2(new_n379_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n424_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n420_), .B1(new_n444_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n426_), .B1(new_n451_), .B2(new_n434_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n435_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT27), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n429_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT100), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n442_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n350_), .B1(new_n438_), .B2(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n289_), .A2(new_n292_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT32), .B(new_n420_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n420_), .A2(KEYINPUT32), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n414_), .A2(new_n462_), .A3(new_n425_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n348_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n424_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n419_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n467_), .A2(KEYINPUT96), .A3(new_n426_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT96), .B1(new_n467_), .B2(new_n426_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n325_), .A2(new_n335_), .A3(new_n332_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n344_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n333_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT98), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n333_), .A2(KEYINPUT98), .A3(new_n334_), .A4(new_n337_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n347_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n338_), .A2(KEYINPUT33), .A3(new_n339_), .A4(new_n346_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n464_), .B1(new_n470_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n442_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n456_), .A2(new_n349_), .A3(new_n396_), .A4(new_n441_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n460_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n228_), .B1(new_n459_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G57gat), .B(G64gat), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n490_));
  XOR2_X1   g289(.A(G71gat), .B(G78gat), .Z(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n490_), .A2(new_n491_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(new_n214_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G231gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G127gat), .B(G155gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT16), .ZN(new_n499_));
  XOR2_X1   g298(.A(G183gat), .B(G211gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n501_), .A2(new_n502_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n497_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(new_n503_), .B2(new_n497_), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT74), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G190gat), .B(G218gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G134gat), .B(G162gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT34), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT35), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n521_), .B2(KEYINPUT9), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT9), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n520_), .A2(KEYINPUT65), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT65), .B1(new_n520_), .B2(new_n523_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n522_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT6), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(G99gat), .A3(G106gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT10), .B(G99gat), .Z(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT64), .B(G106gat), .Z(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n526_), .B(new_n531_), .C1(new_n533_), .C2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT8), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n529_), .B1(G99gat), .B2(G106gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n527_), .A2(KEYINPUT6), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n528_), .A2(new_n530_), .A3(KEYINPUT68), .ZN(new_n542_));
  NOR2_X1   g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT66), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT67), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n543_), .B(new_n544_), .C1(new_n545_), .C2(KEYINPUT7), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI22_X1  g346(.A1(new_n544_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT7), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT66), .B1(new_n549_), .B2(KEYINPUT67), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n541_), .B(new_n542_), .C1(new_n547_), .C2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n521_), .A2(new_n519_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n537_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n537_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n548_), .B(new_n550_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n556_), .B2(new_n531_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n536_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT69), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n560_), .B(new_n536_), .C1(new_n554_), .C2(new_n557_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n218_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT72), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n559_), .A2(KEYINPUT72), .A3(new_n218_), .A4(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI22_X1  g365(.A1(new_n558_), .A2(new_n207_), .B1(KEYINPUT35), .B2(new_n514_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n518_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  AOI211_X1 g368(.A(new_n517_), .B(new_n567_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT36), .B(new_n512_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT73), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n569_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n512_), .A2(KEYINPUT36), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n571_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n566_), .A2(new_n568_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n517_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n566_), .A2(new_n518_), .A3(new_n568_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(KEYINPUT73), .A3(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(new_n574_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n509_), .B1(new_n576_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n573_), .A2(new_n575_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n574_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(KEYINPUT37), .A4(new_n571_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n508_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n494_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT12), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n559_), .A2(new_n561_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n558_), .A2(new_n587_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT12), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n536_), .B(new_n494_), .C1(new_n554_), .C2(new_n557_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n594_), .A2(KEYINPUT70), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT70), .B1(new_n594_), .B2(new_n595_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n590_), .B(new_n593_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT71), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n594_), .A2(new_n595_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT70), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n594_), .A2(KEYINPUT70), .A3(new_n595_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(KEYINPUT71), .A3(new_n590_), .A4(new_n593_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n591_), .A2(new_n594_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n595_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT5), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n614_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n600_), .A2(new_n606_), .A3(new_n609_), .A4(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n615_), .A2(KEYINPUT13), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT13), .B1(new_n615_), .B2(new_n617_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n487_), .A2(KEYINPUT101), .A3(new_n586_), .A4(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n586_), .A2(new_n620_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n622_), .B1(new_n486_), .B2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n348_), .A2(KEYINPUT102), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n348_), .A2(KEYINPUT102), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(G1gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n621_), .A2(new_n624_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n459_), .A2(new_n485_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n583_), .A2(new_n584_), .A3(new_n571_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n620_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n228_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n635_), .A2(new_n507_), .A3(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n639_), .A2(new_n349_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n632_), .B1(G1gat), .B2(new_n640_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n630_), .A2(KEYINPUT103), .A3(new_n631_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT103), .B1(new_n630_), .B2(new_n631_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT104), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n641_), .B(new_n646_), .C1(new_n643_), .C2(new_n642_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1324gat));
  NAND4_X1  g447(.A1(new_n621_), .A2(new_n210_), .A3(new_n437_), .A4(new_n624_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT105), .Z(new_n650_));
  OAI21_X1  g449(.A(G8gat), .B1(new_n639_), .B2(new_n456_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT39), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n650_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  NAND2_X1  g455(.A1(new_n289_), .A2(new_n292_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G15gat), .B1(new_n639_), .B2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT41), .Z(new_n659_));
  NAND2_X1  g458(.A1(new_n621_), .A2(new_n624_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n460_), .A2(new_n268_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n660_), .B2(new_n661_), .ZN(G1326gat));
  OAI21_X1  g461(.A(G22gat), .B1(new_n639_), .B2(new_n442_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT42), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n442_), .A2(G22gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n660_), .B2(new_n665_), .ZN(G1327gat));
  NAND2_X1  g465(.A1(new_n634_), .A2(new_n508_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT109), .Z(new_n668_));
  AND3_X1   g467(.A1(new_n668_), .A2(new_n487_), .A3(new_n620_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n348_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n638_), .A2(new_n508_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n582_), .A2(new_n585_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n350_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n401_), .A2(new_n437_), .A3(KEYINPUT100), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n457_), .B1(new_n442_), .B2(new_n456_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n442_), .A2(new_n437_), .A3(new_n348_), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n476_), .A2(new_n475_), .B1(new_n347_), .B2(new_n478_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(new_n480_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n681_), .A2(new_n464_), .B1(new_n396_), .B2(new_n441_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n657_), .B1(new_n679_), .B2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n674_), .B1(new_n678_), .B2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n673_), .B1(new_n684_), .B2(KEYINPUT107), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n582_), .A2(new_n585_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n485_), .B2(new_n459_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(KEYINPUT43), .ZN(new_n689_));
  AOI211_X1 g488(.A(new_n671_), .B(new_n672_), .C1(new_n685_), .C2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n672_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n684_), .A2(KEYINPUT107), .A3(new_n673_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT43), .B1(new_n687_), .B2(new_n688_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n671_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n672_), .B1(new_n685_), .B2(new_n689_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT108), .B1(new_n697_), .B2(KEYINPUT44), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n690_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n627_), .A2(G29gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n670_), .B1(new_n699_), .B2(new_n700_), .ZN(G1328gat));
  INV_X1    g500(.A(G36gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n669_), .A2(new_n702_), .A3(new_n437_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT45), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT44), .B(new_n691_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n437_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n698_), .B2(new_n696_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n707_), .B2(new_n702_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n704_), .B(KEYINPUT46), .C1(new_n707_), .C2(new_n702_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1329gat));
  AOI21_X1  g511(.A(G43gat), .B1(new_n669_), .B2(new_n460_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n460_), .A2(G43gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n713_), .B1(new_n699_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI211_X1 g517(.A(new_n690_), .B(new_n714_), .C1(new_n696_), .C2(new_n698_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT47), .B1(new_n719_), .B2(new_n713_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1330gat));
  INV_X1    g520(.A(G50gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n401_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT110), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n669_), .A2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n699_), .A2(new_n401_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n722_), .ZN(G1331gat));
  NAND3_X1  g526(.A1(new_n636_), .A2(new_n637_), .A3(new_n507_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n633_), .A2(new_n634_), .A3(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(G57gat), .A3(new_n348_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT112), .ZN(new_n731_));
  INV_X1    g530(.A(G57gat), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n633_), .A2(new_n228_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n586_), .A3(new_n636_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n628_), .B1(new_n734_), .B2(KEYINPUT111), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(KEYINPUT111), .B2(new_n734_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n731_), .B1(new_n732_), .B2(new_n736_), .ZN(G1332gat));
  INV_X1    g536(.A(new_n729_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G64gat), .B1(new_n738_), .B2(new_n456_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT48), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n456_), .A2(G64gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT113), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n734_), .B2(new_n742_), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n738_), .B2(new_n657_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT49), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n657_), .A2(G71gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n734_), .B2(new_n746_), .ZN(G1334gat));
  OAI21_X1  g546(.A(G78gat), .B1(new_n738_), .B2(new_n442_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT50), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n442_), .A2(G78gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n734_), .B2(new_n750_), .ZN(G1335gat));
  NAND3_X1  g550(.A1(new_n636_), .A2(new_n637_), .A3(new_n508_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n685_), .B2(new_n689_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(new_n348_), .ZN(new_n754_));
  INV_X1    g553(.A(G85gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n733_), .A2(new_n668_), .A3(new_n636_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n627_), .A2(new_n755_), .ZN(new_n757_));
  OAI22_X1  g556(.A1(new_n754_), .A2(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(G1336gat));
  NOR3_X1   g557(.A1(new_n756_), .A2(G92gat), .A3(new_n456_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n753_), .A2(new_n437_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(G92gat), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT114), .Z(G1337gat));
  NOR3_X1   g561(.A1(new_n756_), .A2(new_n657_), .A3(new_n533_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n753_), .A2(new_n460_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(G99gat), .ZN(new_n765_));
  NAND2_X1  g564(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(G1338gat));
  INV_X1    g566(.A(new_n752_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n401_), .B(new_n768_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G106gat), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(KEYINPUT116), .A3(G106gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(KEYINPUT52), .A3(new_n773_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n756_), .A2(new_n442_), .A3(new_n535_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT116), .B1(new_n769_), .B2(G106gat), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n774_), .A2(new_n781_), .A3(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT59), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n674_), .A2(new_n637_), .A3(new_n507_), .A4(new_n620_), .ZN(new_n785_));
  XOR2_X1   g584(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n586_), .A2(new_n637_), .A3(new_n620_), .A4(new_n786_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n228_), .A2(new_n617_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n598_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n590_), .A2(new_n594_), .A3(new_n593_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n792_), .A2(KEYINPUT55), .B1(new_n608_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n600_), .A2(new_n606_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n616_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(KEYINPUT56), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n799_), .B(new_n616_), .C1(new_n794_), .C2(new_n796_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n791_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n615_), .A2(new_n617_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n224_), .A2(new_n227_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804_));
  INV_X1    g603(.A(new_n227_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n222_), .B2(new_n203_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n217_), .A2(new_n203_), .A3(new_n219_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n803_), .A2(new_n804_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n805_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n806_), .A2(new_n808_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT118), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n802_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n634_), .B1(new_n801_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT57), .B1(new_n816_), .B2(KEYINPUT119), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  INV_X1    g618(.A(new_n815_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n600_), .A2(new_n795_), .A3(new_n606_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n793_), .A2(new_n608_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n795_), .B2(new_n598_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n614_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n799_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n797_), .A2(KEYINPUT56), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n820_), .B1(new_n827_), .B2(new_n791_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n818_), .B(new_n819_), .C1(new_n828_), .C2(new_n634_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n814_), .A2(new_n617_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(KEYINPUT58), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n686_), .A2(new_n831_), .A3(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n817_), .A2(new_n829_), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n790_), .B1(new_n508_), .B2(new_n836_), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n657_), .B(new_n628_), .C1(new_n458_), .C2(new_n438_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n784_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n508_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n788_), .A2(new_n789_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(KEYINPUT59), .A3(new_n838_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n840_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845_), .B2(new_n637_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n837_), .A2(new_n839_), .ZN(new_n847_));
  INV_X1    g646(.A(G113gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n228_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(G1340gat));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n620_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n847_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n851_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n620_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n851_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT120), .B(new_n853_), .C1(new_n854_), .C2(new_n851_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1341gat));
  OAI21_X1  g658(.A(G127gat), .B1(new_n845_), .B2(new_n508_), .ZN(new_n860_));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n847_), .A2(new_n861_), .A3(new_n507_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1342gat));
  OAI21_X1  g662(.A(G134gat), .B1(new_n845_), .B2(new_n674_), .ZN(new_n864_));
  INV_X1    g663(.A(G134gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n847_), .A2(new_n865_), .A3(new_n634_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1343gat));
  NOR4_X1   g666(.A1(new_n628_), .A2(new_n460_), .A3(new_n442_), .A4(new_n437_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n843_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n637_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT121), .B(G141gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n869_), .A2(new_n620_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n295_), .ZN(G1345gat));
  NOR2_X1   g673(.A1(new_n869_), .A2(new_n508_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT61), .B(G155gat), .Z(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1346gat));
  OAI21_X1  g676(.A(G162gat), .B1(new_n869_), .B2(new_n674_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n634_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n879_), .A2(G162gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n869_), .B2(new_n880_), .ZN(G1347gat));
  NOR4_X1   g680(.A1(new_n657_), .A2(new_n627_), .A3(new_n401_), .A4(new_n456_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n843_), .A2(new_n228_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n244_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n843_), .A2(KEYINPUT122), .A3(new_n228_), .A4(new_n882_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n885_), .A2(new_n886_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT22), .B(G169gat), .Z(new_n890_));
  OAI22_X1  g689(.A1(new_n888_), .A2(new_n889_), .B1(new_n883_), .B2(new_n890_), .ZN(G1348gat));
  AND2_X1   g690(.A1(new_n843_), .A2(new_n882_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n636_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n407_), .A3(new_n507_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n843_), .A2(new_n507_), .A3(new_n882_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n233_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1350gat));
  NOR2_X1   g699(.A1(new_n879_), .A2(new_n231_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n892_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(G190gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n892_), .B2(new_n686_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n904_), .A2(KEYINPUT124), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(KEYINPUT124), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n902_), .B1(new_n905_), .B2(new_n906_), .ZN(G1351gat));
  NOR4_X1   g706(.A1(new_n460_), .A2(new_n456_), .A3(new_n442_), .A4(new_n348_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n843_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n228_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g711(.A1(new_n909_), .A2(new_n620_), .ZN(new_n913_));
  INV_X1    g712(.A(G204gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(KEYINPUT125), .B2(new_n914_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT125), .B(G204gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n913_), .B2(new_n916_), .ZN(G1353gat));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n508_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n910_), .A2(new_n922_), .ZN(new_n923_));
  MUX2_X1   g722(.A(new_n919_), .B(new_n921_), .S(new_n923_), .Z(G1354gat));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n910_), .A2(new_n925_), .A3(new_n634_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n909_), .A2(new_n674_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n925_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n926_), .B(KEYINPUT127), .C1(new_n925_), .C2(new_n927_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1355gat));
endmodule


