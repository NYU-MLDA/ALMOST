//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_;
  XOR2_X1   g000(.A(G64gat), .B(G92gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT25), .B(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT77), .B1(new_n209_), .B2(KEYINPUT26), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(KEYINPUT26), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT26), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(G190gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .A4(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n219_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n217_), .A2(new_n218_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n215_), .A2(new_n224_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT78), .ZN(new_n229_));
  OR2_X1    g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n222_), .A2(new_n230_), .A3(new_n223_), .ZN(new_n231_));
  OR2_X1    g030(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n226_), .B(new_n231_), .C1(new_n234_), .C2(G176gat), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n228_), .A2(new_n229_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n229_), .B1(new_n228_), .B2(new_n235_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT83), .ZN(new_n239_));
  INV_X1    g038(.A(G204gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(G197gat), .ZN(new_n241_));
  INV_X1    g040(.A(G197gat), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT83), .B1(new_n242_), .B2(G204gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(G204gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n241_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G211gat), .ZN(new_n246_));
  INV_X1    g045(.A(G218gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G211gat), .A2(G218gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n245_), .A2(new_n251_), .A3(KEYINPUT21), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT84), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT21), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n255_), .B(new_n241_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n250_), .B1(new_n258_), .B2(new_n255_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n254_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n240_), .A2(G197gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n242_), .A2(G204gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n263_), .A2(KEYINPUT21), .B1(new_n248_), .B2(new_n249_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(KEYINPUT84), .A3(new_n256_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n253_), .B1(new_n260_), .B2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n238_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT19), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT88), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n232_), .A2(new_n271_), .A3(new_n233_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n218_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275_));
  AND3_X1   g074(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n275_), .B1(new_n278_), .B2(new_n230_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT87), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n219_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n275_), .A2(new_n283_), .A3(new_n216_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n213_), .A2(G190gat), .ZN(new_n286_));
  AND2_X1   g085(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n286_), .B(new_n211_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n281_), .B1(new_n285_), .B2(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n289_), .A2(new_n278_), .A3(new_n227_), .A4(new_n219_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(KEYINPUT87), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n280_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n263_), .A2(KEYINPUT21), .ZN(new_n294_));
  AND4_X1   g093(.A1(KEYINPUT84), .A2(new_n256_), .A3(new_n294_), .A4(new_n250_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT84), .B1(new_n264_), .B2(new_n256_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n252_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(KEYINPUT20), .B(new_n270_), .C1(new_n293_), .C2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n267_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT20), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n228_), .A2(new_n235_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT78), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n228_), .A2(new_n229_), .A3(new_n235_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n266_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n270_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n207_), .B1(new_n299_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n305_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n269_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n291_), .A2(KEYINPUT87), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n224_), .A2(new_n281_), .A3(new_n227_), .A4(new_n289_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n310_), .A2(new_n311_), .B1(new_n274_), .B2(new_n279_), .ZN(new_n312_));
  AOI211_X1 g111(.A(new_n300_), .B(new_n269_), .C1(new_n266_), .C2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n303_), .A2(new_n304_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n297_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n309_), .A2(new_n316_), .A3(new_n206_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n307_), .A2(new_n317_), .A3(KEYINPUT90), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n308_), .A2(new_n269_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT90), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n206_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n293_), .A2(new_n297_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n305_), .A2(new_n324_), .A3(KEYINPUT20), .A4(new_n270_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT93), .B(KEYINPUT20), .Z(new_n326_));
  AOI22_X1  g125(.A1(new_n274_), .A2(new_n279_), .B1(new_n285_), .B2(new_n289_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n327_), .B(new_n252_), .C1(new_n296_), .C2(new_n295_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n326_), .B(new_n328_), .C1(new_n238_), .C2(new_n266_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(KEYINPUT94), .A2(new_n325_), .B1(new_n329_), .B2(new_n269_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n329_), .A2(KEYINPUT94), .A3(new_n269_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n207_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT95), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n319_), .B1(new_n320_), .B2(new_n206_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n333_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n323_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT81), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342_));
  AND3_X1   g141(.A1(KEYINPUT80), .A2(G141gat), .A3(G148gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT80), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n346_));
  INV_X1    g145(.A(G141gat), .ZN(new_n347_));
  INV_X1    g146(.A(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(KEYINPUT3), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n347_), .B(new_n348_), .C1(new_n352_), .C2(KEYINPUT82), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n345_), .A2(new_n346_), .A3(new_n351_), .A4(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n350_), .A2(KEYINPUT3), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n340_), .B(new_n341_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n341_), .B(KEYINPUT1), .ZN(new_n358_));
  OAI221_X1 g157(.A(new_n349_), .B1(new_n344_), .B2(new_n343_), .C1(new_n339_), .C2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G78gat), .B(G106gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT86), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n360_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n356_), .A2(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT29), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n297_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G22gat), .B(G50gat), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n357_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT28), .B1(new_n369_), .B2(new_n266_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n368_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n373_));
  OAI211_X1 g172(.A(G228gat), .B(G233gat), .C1(new_n266_), .C2(KEYINPUT85), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n372_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n368_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n366_), .B1(new_n365_), .B2(new_n297_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n369_), .A2(new_n266_), .A3(KEYINPUT28), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n374_), .B1(new_n380_), .B2(new_n371_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n363_), .B1(new_n376_), .B2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G127gat), .B(G134gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G113gat), .B(G120gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n356_), .A2(new_n359_), .A3(new_n385_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(KEYINPUT4), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT91), .B(KEYINPUT0), .Z(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G57gat), .B(G85gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n388_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(new_n386_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(new_n394_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n395_), .A2(new_n401_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n393_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n400_), .B1(new_n407_), .B2(new_n404_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n375_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n363_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n380_), .A2(new_n371_), .A3(new_n374_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n382_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT96), .B1(new_n337_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n318_), .A2(new_n322_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n400_), .B1(new_n403_), .B2(new_n394_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n418_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n419_), .B(new_n420_), .C1(new_n394_), .C2(new_n392_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n408_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT33), .B(new_n400_), .C1(new_n407_), .C2(new_n404_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n416_), .A2(new_n421_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n406_), .A2(new_n408_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n320_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n426_), .B(new_n428_), .C1(new_n427_), .C2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n382_), .A2(new_n413_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n382_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n325_), .A2(KEYINPUT94), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n329_), .A2(new_n269_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n329_), .A2(KEYINPUT94), .A3(new_n269_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n206_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n317_), .A2(KEYINPUT27), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT95), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT96), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n434_), .A2(new_n443_), .A3(new_n444_), .A4(new_n323_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n415_), .A2(new_n433_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT79), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(G71gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT30), .B(G99gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n238_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n314_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n451_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G15gat), .B(G43gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(new_n455_), .A3(new_n451_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n458_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n447_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n458_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n459_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n465_), .B2(new_n456_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n460_), .A2(new_n466_), .A3(KEYINPUT79), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n385_), .B(KEYINPUT31), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n463_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n447_), .B(new_n470_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n446_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n469_), .A2(new_n409_), .A3(new_n471_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n432_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n474_), .A2(new_n337_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT76), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G229gat), .A2(G233gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT71), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(G1gat), .B2(G8gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT72), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G1gat), .B(G8gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n489_), .A2(new_n492_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n481_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n489_), .A2(new_n492_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G43gat), .B(G50gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(new_n490_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT15), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n492_), .A2(KEYINPUT15), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n496_), .B(new_n480_), .C1(new_n489_), .C2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT75), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n495_), .A2(new_n504_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n495_), .B2(new_n504_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n479_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n495_), .A2(new_n504_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n508_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n495_), .A2(new_n504_), .A3(new_n509_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(KEYINPUT76), .A3(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518_));
  INV_X1    g317(.A(G99gat), .ZN(new_n519_));
  INV_X1    g318(.A(G106gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT6), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n521_), .A2(new_n524_), .A3(new_n525_), .A4(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G85gat), .B(G92gat), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT8), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT8), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT10), .B(G99gat), .Z(new_n533_));
  INV_X1    g332(.A(KEYINPUT64), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT10), .B(G99gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT64), .ZN(new_n537_));
  AOI21_X1  g336(.A(G106gat), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n524_), .A2(new_n525_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G85gat), .A2(G92gat), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(KEYINPUT9), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n528_), .A2(KEYINPUT9), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  OAI22_X1  g343(.A1(new_n530_), .A2(new_n532_), .B1(new_n538_), .B2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G71gat), .B(G78gat), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G57gat), .B(G64gat), .Z(new_n548_));
  INV_X1    g347(.A(KEYINPUT11), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G57gat), .B(G64gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT11), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n547_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n546_), .B1(KEYINPUT11), .B2(new_n551_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n545_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n529_), .B(KEYINPUT8), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n536_), .B(new_n534_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n542_), .B(new_n543_), .C1(new_n558_), .C2(G106gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n553_), .A2(new_n554_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n556_), .A2(new_n561_), .A3(KEYINPUT12), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n545_), .A2(new_n555_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n556_), .A2(new_n561_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n566_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT66), .ZN(new_n573_));
  XOR2_X1   g372(.A(G176gat), .B(G204gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT65), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n571_), .A2(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT13), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n585_), .B(new_n586_), .Z(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n502_), .A2(new_n545_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n557_), .A2(new_n492_), .A3(new_n559_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n590_), .A2(new_n591_), .A3(new_n594_), .A4(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT67), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n590_), .A2(new_n591_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n594_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  AOI211_X1 g400(.A(KEYINPUT67), .B(new_n594_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n589_), .B(new_n597_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n597_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT68), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n587_), .B(KEYINPUT36), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n584_), .B(new_n603_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT69), .ZN(new_n611_));
  INV_X1    g410(.A(new_n597_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n599_), .A2(new_n600_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT67), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n599_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n608_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n603_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n611_), .B1(new_n618_), .B2(KEYINPUT37), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n610_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(KEYINPUT68), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n622_), .A2(new_n611_), .A3(new_n584_), .A4(new_n603_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT70), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n620_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n489_), .B(KEYINPUT73), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n560_), .B(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n627_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(new_n246_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT16), .B(G183gat), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(KEYINPUT17), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(KEYINPUT17), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n630_), .A2(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT74), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n634_), .A2(KEYINPUT17), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n638_), .B(KEYINPUT74), .C1(new_n640_), .C2(new_n630_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n625_), .A2(new_n626_), .A3(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n478_), .A2(new_n517_), .A3(new_n583_), .A4(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n426_), .B(KEYINPUT97), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n645_), .A2(G1gat), .A3(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT98), .Z(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n649_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n476_), .B1(new_n446_), .B2(new_n472_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n583_), .A2(new_n517_), .A3(new_n642_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n622_), .A2(new_n603_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G1gat), .B1(new_n660_), .B2(new_n409_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n650_), .A2(new_n651_), .A3(new_n661_), .ZN(G1324gat));
  INV_X1    g461(.A(new_n655_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n478_), .A2(new_n663_), .A3(new_n337_), .A4(new_n659_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT100), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n656_), .A2(new_n666_), .A3(new_n337_), .A4(new_n659_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(G8gat), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT39), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT101), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n665_), .A2(new_n667_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT39), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n671_), .A2(KEYINPUT102), .A3(new_n672_), .A4(G8gat), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT101), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n668_), .A2(new_n674_), .A3(KEYINPUT39), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n668_), .B2(KEYINPUT39), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n670_), .A2(new_n673_), .A3(new_n675_), .A4(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n337_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n645_), .A2(G8gat), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n678_), .A2(KEYINPUT40), .A3(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1325gat));
  OAI21_X1  g484(.A(G15gat), .B1(new_n660_), .B2(new_n472_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT41), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n645_), .A2(G15gat), .A3(new_n472_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1326gat));
  OAI21_X1  g488(.A(G22gat), .B1(new_n660_), .B2(new_n432_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT42), .Z(new_n691_));
  NOR3_X1   g490(.A1(new_n645_), .A2(G22gat), .A3(new_n432_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT103), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n583_), .A2(new_n517_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(new_n642_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n625_), .A2(new_n626_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n478_), .B2(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n652_), .A2(KEYINPUT43), .A3(new_n698_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n696_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT44), .B(new_n696_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n646_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n643_), .A2(new_n658_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n652_), .A2(new_n695_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(G29gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n426_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(G1328gat));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n709_), .A2(new_n713_), .A3(new_n337_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n714_), .B(new_n715_), .Z(new_n716_));
  NOR2_X1   g515(.A1(new_n706_), .A2(new_n679_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n713_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(G1329gat));
  INV_X1    g519(.A(new_n472_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G43gat), .B1(new_n709_), .B2(new_n721_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT106), .Z(new_n723_));
  NAND4_X1  g522(.A1(new_n704_), .A2(G43gat), .A3(new_n721_), .A4(new_n705_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n724_), .A2(new_n725_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT107), .B(KEYINPUT108), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT47), .Z(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n723_), .B(new_n730_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1330gat));
  OAI21_X1  g533(.A(G50gat), .B1(new_n706_), .B2(new_n432_), .ZN(new_n735_));
  INV_X1    g534(.A(G50gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n709_), .A2(new_n736_), .A3(new_n475_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1331gat));
  NOR3_X1   g537(.A1(new_n652_), .A2(new_n517_), .A3(new_n583_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(new_n642_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n698_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n646_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(KEYINPUT109), .A3(new_n698_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747_));
  INV_X1    g546(.A(G57gat), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n746_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n739_), .A2(new_n642_), .A3(new_n657_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(G57gat), .A3(new_n426_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT111), .Z(new_n753_));
  NOR3_X1   g552(.A1(new_n749_), .A2(new_n750_), .A3(new_n753_), .ZN(G1332gat));
  INV_X1    g553(.A(G64gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n751_), .B2(new_n337_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT48), .Z(new_n757_));
  AND2_X1   g556(.A1(new_n743_), .A2(new_n745_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n755_), .A3(new_n337_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1333gat));
  AOI21_X1  g559(.A(new_n449_), .B1(new_n751_), .B2(new_n721_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT49), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(new_n449_), .A3(new_n721_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n751_), .A2(new_n475_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G78gat), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT112), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT112), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n769_));
  OR3_X1    g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(G78gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n758_), .A2(new_n771_), .A3(new_n475_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n769_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n772_), .A3(new_n773_), .ZN(G1335gat));
  INV_X1    g573(.A(new_n708_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n739_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(G85gat), .B1(new_n777_), .B2(new_n744_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n583_), .A2(new_n517_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n643_), .B(new_n779_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(new_n409_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n778_), .B1(new_n781_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g581(.A(G92gat), .B1(new_n777_), .B2(new_n337_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT113), .ZN(new_n784_));
  INV_X1    g583(.A(new_n780_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n337_), .A2(G92gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(G1337gat));
  NOR3_X1   g586(.A1(new_n776_), .A2(new_n558_), .A3(new_n472_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n721_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(G99gat), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT51), .Z(G1338gat));
  OAI21_X1  g590(.A(G106gat), .B1(new_n780_), .B2(new_n432_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT114), .B(G106gat), .C1(new_n780_), .C2(new_n432_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(KEYINPUT52), .A3(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n777_), .A2(new_n520_), .A3(new_n475_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n792_), .A2(new_n793_), .A3(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n797_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n796_), .A2(new_n802_), .A3(new_n797_), .A4(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1339gat));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n512_), .A2(new_n516_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n567_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT116), .B1(new_n565_), .B2(new_n566_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n562_), .A2(new_n810_), .A3(new_n569_), .A4(new_n564_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n565_), .A2(KEYINPUT55), .A3(new_n566_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n808_), .A2(new_n809_), .A3(new_n811_), .A4(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT117), .B1(new_n813_), .B2(new_n578_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n806_), .B1(KEYINPUT56), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n578_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n579_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n480_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n496_), .B1(new_n489_), .B2(new_n503_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n821_), .B(new_n508_), .C1(new_n480_), .C2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n515_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n815_), .A2(new_n820_), .B1(new_n582_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n805_), .B1(new_n826_), .B2(new_n658_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n813_), .A2(new_n578_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n824_), .B1(new_n828_), .B2(new_n819_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n579_), .B1(new_n816_), .B2(KEYINPUT56), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(KEYINPUT58), .A3(new_n830_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n833_), .B(new_n834_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n582_), .A2(new_n825_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n517_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n580_), .B1(new_n814_), .B2(KEYINPUT56), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT57), .A3(new_n657_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n827_), .A2(new_n835_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n643_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n644_), .A2(new_n806_), .A3(new_n583_), .A4(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n843_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n620_), .A2(new_n623_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT70), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n620_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n847_), .A2(new_n806_), .A3(new_n848_), .A4(new_n642_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n583_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n845_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n844_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n842_), .A2(new_n852_), .ZN(new_n853_));
  NOR4_X1   g652(.A1(new_n472_), .A2(new_n337_), .A3(new_n646_), .A4(new_n475_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT118), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G113gat), .B1(new_n857_), .B2(new_n517_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n842_), .A2(KEYINPUT120), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n841_), .A2(new_n860_), .A3(new_n643_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n852_), .A3(new_n861_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n855_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n856_), .A2(KEYINPUT59), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n867_), .A2(G113gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n858_), .B1(new_n868_), .B2(new_n517_), .ZN(G1340gat));
  OAI21_X1  g668(.A(G120gat), .B1(new_n866_), .B2(new_n583_), .ZN(new_n870_));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n583_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n857_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n871_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(G1341gat));
  INV_X1    g673(.A(G127gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n856_), .B2(new_n643_), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(KEYINPUT121), .Z(new_n877_));
  NOR3_X1   g676(.A1(new_n866_), .A2(new_n875_), .A3(new_n643_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1342gat));
  AOI21_X1  g678(.A(G134gat), .B1(new_n857_), .B2(new_n658_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT122), .B(G134gat), .Z(new_n881_));
  NOR2_X1   g680(.A1(new_n698_), .A2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n867_), .B2(new_n882_), .ZN(G1343gat));
  AOI211_X1 g682(.A(new_n721_), .B(new_n432_), .C1(new_n842_), .C2(new_n852_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n679_), .A2(new_n744_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n806_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n347_), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n583_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n348_), .ZN(G1345gat));
  OR3_X1    g690(.A1(new_n887_), .A2(KEYINPUT123), .A3(new_n643_), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT123), .B1(new_n887_), .B2(new_n643_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1346gat));
  INV_X1    g696(.A(new_n887_), .ZN(new_n898_));
  AOI21_X1  g697(.A(G162gat), .B1(new_n898_), .B2(new_n658_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n887_), .A2(new_n698_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(G162gat), .B2(new_n900_), .ZN(G1347gat));
  NOR4_X1   g700(.A1(new_n679_), .A2(new_n744_), .A3(new_n472_), .A4(new_n475_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n862_), .A2(new_n517_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(G169gat), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n904_), .A2(KEYINPUT62), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(KEYINPUT62), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n841_), .A2(new_n860_), .A3(new_n643_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n860_), .B1(new_n841_), .B2(new_n643_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n844_), .A2(new_n851_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n902_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT124), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n862_), .A2(new_n913_), .A3(new_n902_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n517_), .B1(new_n273_), .B2(new_n272_), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT125), .Z(new_n918_));
  OAI22_X1  g717(.A1(new_n905_), .A2(new_n906_), .B1(new_n916_), .B2(new_n918_), .ZN(G1348gat));
  AOI21_X1  g718(.A(new_n911_), .B1(new_n842_), .B2(new_n852_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(G176gat), .A3(new_n850_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT126), .Z(new_n922_));
  NAND2_X1  g721(.A1(new_n915_), .A2(new_n850_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n218_), .ZN(G1349gat));
  NOR3_X1   g723(.A1(new_n916_), .A2(new_n643_), .A3(new_n208_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G183gat), .B1(new_n920_), .B2(new_n642_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1350gat));
  NAND4_X1  g726(.A1(new_n915_), .A2(new_n286_), .A3(new_n211_), .A4(new_n658_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n698_), .B1(new_n912_), .B2(new_n914_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n929_), .A2(new_n930_), .A3(new_n209_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n862_), .A2(new_n913_), .A3(new_n902_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n913_), .B1(new_n862_), .B2(new_n902_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n699_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(KEYINPUT127), .B1(new_n934_), .B2(G190gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n928_), .B1(new_n931_), .B2(new_n935_), .ZN(G1351gat));
  NOR2_X1   g735(.A1(new_n679_), .A2(new_n426_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n884_), .A2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n806_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(new_n242_), .ZN(G1352gat));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n583_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(new_n240_), .ZN(G1353gat));
  NOR2_X1   g741(.A1(new_n938_), .A2(new_n643_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n943_), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n946_), .B1(new_n943_), .B2(new_n944_), .ZN(G1354gat));
  NOR3_X1   g746(.A1(new_n938_), .A2(new_n247_), .A3(new_n698_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n884_), .A2(new_n658_), .A3(new_n937_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n948_), .B1(new_n247_), .B2(new_n949_), .ZN(G1355gat));
endmodule


