//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(G113gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G120gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT3), .Z(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n212_), .B(KEYINPUT2), .Z(new_n213_));
  OAI21_X1  g012(.A(new_n209_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n210_), .B1(new_n209_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(new_n212_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n206_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n204_), .B(G120gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n219_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n223_), .A3(KEYINPUT4), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G225gat), .A2(G233gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT100), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n224_), .B(new_n226_), .C1(KEYINPUT4), .C2(new_n223_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n221_), .A2(new_n223_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n226_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G1gat), .B(G29gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G85gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n227_), .A2(new_n230_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT104), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G99gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G15gat), .B(G43gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G169gat), .B(G176gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT25), .B(G183gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT26), .B(G190gat), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n251_), .A2(KEYINPUT24), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT23), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OR3_X1    g058(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n254_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT22), .B(G169gat), .ZN(new_n262_));
  INV_X1    g061(.A(G176gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(KEYINPUT87), .A3(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n257_), .B(new_n258_), .C1(G183gat), .C2(G190gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n266_));
  OAI21_X1  g065(.A(G169gat), .B1(new_n266_), .B2(G176gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n206_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n269_), .B(KEYINPUT30), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n222_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n250_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(new_n274_), .A3(new_n250_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n246_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n246_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n279_), .A2(new_n275_), .A3(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n243_), .B1(new_n278_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G197gat), .B(G204gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT21), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n284_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n288_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n285_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n292_), .B1(new_n220_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G78gat), .B(G106gat), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G228gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT92), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT91), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n292_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(new_n295_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n296_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n300_), .B1(new_n296_), .B2(new_n301_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT93), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n294_), .B(new_n295_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n300_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT93), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n302_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G22gat), .B(G50gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n305_), .A2(new_n310_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n317_), .A2(new_n309_), .A3(new_n302_), .A4(new_n308_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n276_), .A2(new_n246_), .A3(new_n277_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n280_), .B1(new_n279_), .B2(new_n275_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(KEYINPUT89), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n282_), .A2(new_n316_), .A3(new_n318_), .A4(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(new_n318_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n320_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n242_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT94), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n259_), .A2(new_n327_), .A3(new_n260_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n260_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT94), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n254_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT95), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n254_), .A2(new_n328_), .A3(new_n330_), .A4(KEYINPUT95), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n262_), .B(KEYINPUT96), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n335_), .B(new_n265_), .C1(new_n336_), .C2(G176gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n292_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n290_), .B(new_n286_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(new_n261_), .A3(new_n268_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(KEYINPUT20), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT97), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT19), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n340_), .A2(new_n337_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n347_), .A2(KEYINPUT98), .A3(new_n333_), .A4(new_n334_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n345_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT98), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n340_), .A2(new_n337_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n333_), .A2(new_n334_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n269_), .B2(new_n292_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n348_), .A2(new_n349_), .A3(new_n353_), .A4(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT20), .B1(new_n269_), .B2(new_n292_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(new_n292_), .B2(new_n338_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT97), .B1(new_n358_), .B2(new_n349_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n346_), .A2(new_n356_), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT18), .B(G64gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G92gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n346_), .A2(new_n356_), .A3(new_n359_), .A4(new_n364_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(KEYINPUT99), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT99), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n360_), .A2(new_n369_), .A3(new_n365_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n371_), .A2(KEYINPUT27), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n347_), .A2(new_n331_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n355_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n345_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n345_), .B2(new_n342_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n365_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(KEYINPUT27), .A3(new_n367_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n326_), .A2(new_n372_), .A3(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n227_), .A2(KEYINPUT33), .A3(new_n230_), .A4(new_n238_), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n380_), .B(KEYINPUT102), .Z(new_n381_));
  NAND2_X1  g180(.A1(new_n228_), .A2(new_n226_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n224_), .B1(KEYINPUT4), .B2(new_n223_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n236_), .B(new_n382_), .C1(new_n383_), .C2(new_n226_), .ZN(new_n384_));
  XOR2_X1   g183(.A(KEYINPUT103), .B(KEYINPUT33), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n239_), .A2(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n371_), .A2(new_n381_), .A3(new_n384_), .A4(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n376_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n240_), .B(new_n389_), .C1(new_n388_), .C2(new_n360_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n282_), .A2(new_n321_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n323_), .A3(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n379_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G57gat), .ZN(new_n396_));
  INV_X1    g195(.A(G64gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT11), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G57gat), .A2(G64gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G71gat), .A2(G78gat), .ZN(new_n402_));
  INV_X1    g201(.A(G71gat), .ZN(new_n403_));
  INV_X1    g202(.A(G78gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n401_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT67), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT67), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n401_), .A2(new_n408_), .A3(new_n402_), .A4(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n398_), .A2(new_n400_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n411_), .A2(new_n399_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n407_), .A2(new_n412_), .A3(new_n409_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G231gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G1gat), .B(G8gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT79), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G15gat), .B(G22gat), .ZN(new_n421_));
  INV_X1    g220(.A(G1gat), .ZN(new_n422_));
  INV_X1    g221(.A(G8gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT14), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n419_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n425_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n418_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G127gat), .B(G155gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G183gat), .B(G211gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT17), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n432_), .A2(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n440_), .B(KEYINPUT81), .Z(new_n441_));
  XNOR2_X1  g240(.A(new_n432_), .B(KEYINPUT82), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n438_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n439_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT66), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT8), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT7), .ZN(new_n448_));
  INV_X1    g247(.A(G99gat), .ZN(new_n449_));
  INV_X1    g248(.A(G106gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT65), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(KEYINPUT6), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n457_), .A2(KEYINPUT65), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n454_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(KEYINPUT65), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(KEYINPUT6), .ZN(new_n461_));
  AND2_X1   g260(.A1(G99gat), .A2(G106gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n453_), .B1(new_n459_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G85gat), .B(G92gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n446_), .B(new_n447_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(KEYINPUT9), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(KEYINPUT64), .ZN(new_n469_));
  XOR2_X1   g268(.A(KEYINPUT10), .B(G99gat), .Z(new_n470_));
  AOI22_X1  g269(.A1(new_n467_), .A2(new_n469_), .B1(new_n470_), .B2(new_n450_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n459_), .A2(new_n463_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n451_), .A2(new_n452_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n462_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n465_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n446_), .A2(new_n447_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .A4(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G50gat), .ZN(new_n483_));
  INV_X1    g282(.A(G43gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT73), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT73), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G43gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n483_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(new_n487_), .A3(new_n483_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G29gat), .B(G36gat), .Z(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n491_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n490_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n493_), .B1(new_n494_), .B2(new_n488_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n466_), .A2(new_n474_), .A3(new_n482_), .A4(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT72), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT34), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT35), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n500_), .A2(new_n501_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n466_), .A2(new_n474_), .A3(new_n482_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n492_), .A2(new_n495_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT15), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n496_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n504_), .A2(new_n506_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT74), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n497_), .A2(new_n515_), .A3(new_n502_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n512_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n497_), .B2(new_n502_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n505_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT75), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT75), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n521_), .B(new_n505_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n514_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G190gat), .B(G218gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G134gat), .ZN(new_n525_));
  INV_X1    g324(.A(G162gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT36), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT77), .B1(new_n523_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n522_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n503_), .A2(KEYINPUT74), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(new_n516_), .A3(new_n512_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n521_), .B1(new_n533_), .B2(new_n505_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n513_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT77), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n528_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n530_), .A2(new_n537_), .A3(KEYINPUT37), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT36), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n527_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n541_), .B(new_n513_), .C1(new_n531_), .C2(new_n534_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT76), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT76), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n523_), .A2(new_n544_), .A3(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n538_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n535_), .A2(KEYINPUT78), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT78), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n523_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n528_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT37), .B1(new_n551_), .B2(new_n542_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n395_), .A2(new_n445_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT13), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n466_), .A2(new_n474_), .A3(new_n482_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT68), .B1(new_n558_), .B2(new_n416_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT12), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n407_), .A2(new_n412_), .A3(new_n409_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n412_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(new_n507_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n507_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(KEYINPUT68), .A3(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n560_), .A2(new_n561_), .A3(new_n566_), .A4(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n567_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n561_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  INV_X1    g374(.A(G204gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT5), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n263_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(G176gat), .A3(new_n580_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n582_), .A2(new_n583_), .A3(KEYINPUT69), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT69), .B1(new_n582_), .B2(new_n583_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT70), .B1(new_n574_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT70), .ZN(new_n589_));
  AOI211_X1 g388(.A(new_n589_), .B(new_n586_), .C1(new_n570_), .C2(new_n573_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n582_), .A2(new_n583_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n570_), .A2(new_n573_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n557_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  NOR4_X1   g394(.A1(new_n588_), .A2(new_n590_), .A3(new_n595_), .A4(KEYINPUT71), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n556_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n574_), .A2(new_n587_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n589_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n574_), .A2(KEYINPUT70), .A3(new_n587_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n593_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT71), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n591_), .A2(new_n557_), .A3(new_n593_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(KEYINPUT13), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G169gat), .B(G197gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(G141gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT84), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(new_n203_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n431_), .A2(new_n508_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n496_), .A2(new_n430_), .A3(new_n426_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT83), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n609_), .A2(KEYINPUT83), .A3(new_n610_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n509_), .A2(new_n511_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n431_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n614_), .B(new_n610_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n608_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n620_), .A3(new_n608_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT85), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT86), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n622_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT86), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n621_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n597_), .A2(new_n604_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n555_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n422_), .A3(new_n242_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT105), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n635_), .A2(KEYINPUT106), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n634_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n551_), .A2(new_n542_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n445_), .B(new_n647_), .C1(new_n379_), .C2(new_n394_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n242_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n640_), .A2(new_n641_), .A3(new_n652_), .ZN(G1324gat));
  NAND2_X1  g452(.A1(new_n372_), .A2(new_n378_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n648_), .A2(new_n654_), .A3(new_n644_), .A4(new_n642_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G8gat), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT107), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(KEYINPUT107), .A3(G8gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(KEYINPUT39), .A3(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n636_), .A2(new_n423_), .A3(new_n654_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n656_), .A2(new_n657_), .A3(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT108), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n660_), .A2(new_n666_), .A3(new_n661_), .A4(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(KEYINPUT40), .A3(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  INV_X1    g471(.A(G15gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n649_), .B2(new_n392_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT41), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n636_), .A2(new_n673_), .A3(new_n392_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1326gat));
  INV_X1    g476(.A(G22gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n323_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n649_), .B2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT42), .Z(new_n681_));
  NAND3_X1  g480(.A1(new_n636_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1327gat));
  AND2_X1   g482(.A1(new_n441_), .A2(new_n444_), .ZN(new_n684_));
  NOR4_X1   g483(.A1(new_n395_), .A2(new_n634_), .A3(new_n684_), .A4(new_n646_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G29gat), .B1(new_n685_), .B2(new_n242_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n395_), .A2(new_n553_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n554_), .A2(KEYINPUT109), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT43), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT43), .B(new_n688_), .C1(new_n395_), .C2(new_n553_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n445_), .A3(new_n645_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(G29gat), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n692_), .A2(KEYINPUT44), .A3(new_n445_), .A4(new_n645_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(new_n242_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n686_), .B1(new_n696_), .B2(new_n698_), .ZN(G1328gat));
  INV_X1    g498(.A(G36gat), .ZN(new_n700_));
  INV_X1    g499(.A(new_n654_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n700_), .B1(new_n702_), .B2(new_n697_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n685_), .A2(new_n700_), .A3(new_n654_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  OR3_X1    g506(.A1(new_n703_), .A2(new_n704_), .A3(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n703_), .B2(new_n707_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  NAND4_X1  g509(.A1(new_n695_), .A2(G43gat), .A3(new_n324_), .A4(new_n697_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n685_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n484_), .B1(new_n712_), .B2(new_n393_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g514(.A1(new_n685_), .A2(new_n483_), .A3(new_n679_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n695_), .A2(new_n679_), .A3(new_n697_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(KEYINPUT111), .A3(G50gat), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT111), .B1(new_n717_), .B2(G50gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1331gat));
  AND2_X1   g520(.A1(new_n597_), .A2(new_n604_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(new_n633_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n648_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(G57gat), .A3(new_n242_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT112), .Z(new_n726_));
  NAND2_X1  g525(.A1(new_n555_), .A2(new_n723_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n242_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n726_), .A2(new_n729_), .ZN(G1332gat));
  AOI21_X1  g529(.A(new_n397_), .B1(new_n724_), .B2(new_n654_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT113), .Z(new_n732_));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n733_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n728_), .A2(new_n397_), .A3(new_n654_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(G1333gat));
  AOI21_X1  g536(.A(new_n403_), .B1(new_n724_), .B2(new_n392_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT49), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n728_), .A2(new_n403_), .A3(new_n392_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1334gat));
  AOI21_X1  g540(.A(new_n404_), .B1(new_n724_), .B2(new_n679_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT50), .Z(new_n743_));
  NAND2_X1  g542(.A1(new_n679_), .A2(new_n404_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT114), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n727_), .B2(new_n745_), .ZN(G1335gat));
  INV_X1    g545(.A(G85gat), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n395_), .A2(new_n646_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n722_), .A2(new_n633_), .A3(new_n684_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n750_), .B2(new_n651_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT115), .Z(new_n752_));
  INV_X1    g551(.A(new_n749_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n755_), .A2(new_n747_), .A3(new_n651_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n752_), .A2(new_n756_), .ZN(G1336gat));
  INV_X1    g556(.A(new_n750_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G92gat), .B1(new_n758_), .B2(new_n654_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n654_), .A2(G92gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n754_), .B2(new_n760_), .ZN(G1337gat));
  NAND3_X1  g560(.A1(new_n758_), .A2(new_n470_), .A3(new_n324_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT116), .Z(new_n763_));
  AOI21_X1  g562(.A(new_n449_), .B1(new_n754_), .B2(new_n392_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n764_), .A2(KEYINPUT117), .ZN(new_n765_));
  OR3_X1    g564(.A1(new_n763_), .A2(new_n765_), .A3(KEYINPUT51), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT51), .B1(new_n763_), .B2(new_n765_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1338gat));
  NAND3_X1  g567(.A1(new_n758_), .A2(new_n450_), .A3(new_n679_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n754_), .A2(new_n679_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G106gat), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT52), .B(new_n450_), .C1(new_n754_), .C2(new_n679_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g574(.A1(new_n597_), .A2(new_n684_), .A3(new_n604_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n538_), .A2(new_n546_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT37), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n646_), .A2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n628_), .A2(new_n632_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  OR3_X1    g580(.A1(new_n776_), .A2(new_n781_), .A3(KEYINPUT118), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n547_), .A2(new_n552_), .A3(new_n633_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n784_), .A2(new_n604_), .A3(new_n597_), .A4(new_n684_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n785_), .B2(KEYINPUT118), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT118), .B(new_n783_), .C1(new_n776_), .C2(new_n781_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n782_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n608_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n615_), .B(new_n610_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n623_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n568_), .B1(new_n567_), .B2(KEYINPUT68), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT68), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n799_), .B(KEYINPUT12), .C1(new_n564_), .C2(new_n507_), .ZN(new_n800_));
  NOR4_X1   g599(.A1(new_n798_), .A2(new_n800_), .A3(new_n572_), .A4(new_n565_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n560_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n572_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(KEYINPUT55), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n802_), .A2(new_n805_), .A3(new_n572_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n587_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n797_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT56), .B(new_n587_), .C1(new_n804_), .C2(new_n806_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n780_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n593_), .B1(new_n810_), .B2(KEYINPUT119), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n796_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n790_), .B1(new_n814_), .B2(new_n647_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n798_), .A2(new_n800_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n561_), .B1(new_n816_), .B2(new_n566_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n570_), .B1(new_n817_), .B2(new_n805_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n806_), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n808_), .B(new_n586_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n595_), .B1(new_n820_), .B2(KEYINPUT120), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n807_), .A2(new_n808_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n810_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n795_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n821_), .A2(new_n824_), .A3(KEYINPUT58), .A4(new_n825_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n554_), .A3(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n825_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n586_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT119), .B1(new_n832_), .B2(KEYINPUT56), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n633_), .B1(new_n833_), .B2(new_n820_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n831_), .B1(new_n834_), .B2(new_n812_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(KEYINPUT57), .A3(new_n646_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n815_), .A2(new_n830_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n445_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n679_), .B1(new_n789_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n701_), .A2(new_n324_), .A3(new_n242_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n203_), .B1(new_n842_), .B2(new_n780_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n843_), .A2(KEYINPUT121), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(KEYINPUT121), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n789_), .A2(new_n838_), .ZN(new_n846_));
  AND4_X1   g645(.A1(KEYINPUT59), .A2(new_n846_), .A3(new_n323_), .A4(new_n841_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT59), .B1(new_n839_), .B2(new_n841_), .ZN(new_n848_));
  OAI211_X1 g647(.A(G113gat), .B(new_n633_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n844_), .A2(new_n845_), .A3(new_n849_), .ZN(G1340gat));
  INV_X1    g649(.A(new_n722_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT122), .B(new_n851_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(G120gat), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n842_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n205_), .B1(new_n722_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n857_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n205_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n859_), .ZN(G1341gat));
  AOI21_X1  g659(.A(G127gat), .B1(new_n857_), .B2(new_n684_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n847_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n848_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n445_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n864_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g664(.A(G134gat), .B1(new_n857_), .B2(new_n647_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n553_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g667(.A1(new_n654_), .A2(new_n651_), .A3(new_n322_), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n869_), .B(KEYINPUT123), .Z(new_n870_));
  NAND2_X1  g669(.A1(new_n846_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n633_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n851_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g675(.A1(new_n871_), .A2(new_n445_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT61), .B(G155gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  NOR3_X1   g678(.A1(new_n871_), .A2(new_n526_), .A3(new_n553_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n872_), .A2(new_n647_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n526_), .B2(new_n881_), .ZN(G1347gat));
  NOR3_X1   g681(.A1(new_n701_), .A2(new_n393_), .A3(new_n242_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n846_), .A2(new_n633_), .A3(new_n323_), .A4(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G169gat), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n884_), .A2(new_n336_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n884_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n887_), .A2(new_n888_), .A3(KEYINPUT124), .A4(new_n889_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1348gat));
  NAND2_X1  g693(.A1(new_n839_), .A2(new_n883_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n722_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n263_), .ZN(G1349gat));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n445_), .ZN(new_n898_));
  MUX2_X1   g697(.A(G183gat), .B(new_n252_), .S(new_n898_), .Z(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n895_), .B2(new_n553_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n839_), .A2(new_n253_), .A3(new_n883_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n646_), .B2(new_n901_), .ZN(G1351gat));
  NOR2_X1   g701(.A1(new_n322_), .A2(new_n242_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n701_), .B1(new_n903_), .B2(KEYINPUT125), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n903_), .A2(KEYINPUT125), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n846_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n633_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g707(.A1(new_n846_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n722_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n576_), .ZN(G1353gat));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n912_));
  INV_X1    g711(.A(G211gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n906_), .A2(new_n684_), .A3(new_n914_), .A4(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n912_), .B(new_n913_), .C1(new_n909_), .C2(new_n445_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1354gat));
  AOI21_X1  g719(.A(G218gat), .B1(new_n906_), .B2(new_n647_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n909_), .A2(new_n553_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(G218gat), .B2(new_n922_), .ZN(G1355gat));
endmodule


