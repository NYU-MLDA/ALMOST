//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  INV_X1    g005(.A(G92gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G85gat), .B(G92gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT9), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT64), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(KEYINPUT9), .B2(new_n207_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n213_), .B(new_n214_), .C1(KEYINPUT9), .C2(new_n210_), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT6), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT6), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT10), .B(G99gat), .Z(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n217_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n212_), .A2(new_n215_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(KEYINPUT65), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT7), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n218_), .A2(new_n220_), .A3(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n225_), .B1(new_n231_), .B2(new_n206_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n221_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n225_), .A3(new_n206_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n224_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G29gat), .B(G36gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G43gat), .B(G50gat), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT15), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT7), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n227_), .B(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n229_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n210_), .B1(new_n247_), .B2(new_n230_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n234_), .B1(new_n248_), .B2(new_n225_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n241_), .A3(new_n224_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G232gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT34), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT35), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n243_), .A2(new_n250_), .A3(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n253_), .A2(new_n254_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n257_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n205_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(KEYINPUT72), .A3(new_n259_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n258_), .A2(KEYINPUT72), .A3(new_n259_), .A4(new_n262_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n260_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT37), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(KEYINPUT73), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(KEYINPUT73), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n266_), .A2(KEYINPUT73), .A3(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G127gat), .B(G155gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT16), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G183gat), .B(G211gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT17), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT75), .ZN(new_n280_));
  XOR2_X1   g079(.A(G71gat), .B(G78gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(G57gat), .B(G64gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n281_), .B1(KEYINPUT11), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n284_), .A3(KEYINPUT11), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n282_), .B2(KEYINPUT11), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n283_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n282_), .A2(KEYINPUT11), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT66), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n282_), .A2(KEYINPUT11), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n281_), .A4(new_n285_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  INV_X1    g093(.A(G1gat), .ZN(new_n295_));
  INV_X1    g094(.A(G8gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G8gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n293_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G231gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n280_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT17), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n278_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(KEYINPUT74), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n306_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n304_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n274_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n236_), .A2(KEYINPUT12), .A3(new_n293_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n293_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n249_), .A2(new_n315_), .A3(new_n224_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n315_), .B1(new_n249_), .B2(new_n224_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT68), .B1(new_n318_), .B2(KEYINPUT12), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT12), .B1(new_n236_), .B2(new_n293_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n317_), .A2(new_n319_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n236_), .A2(new_n293_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT67), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n316_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n323_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n327_), .B(new_n328_), .C1(new_n326_), .C2(new_n325_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G176gat), .B(G204gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT70), .ZN(new_n331_));
  XOR2_X1   g130(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G120gat), .B(G148gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n324_), .A2(new_n329_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n324_), .B2(new_n329_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(new_n340_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT13), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT13), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n313_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT76), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G227gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(G15gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G71gat), .ZN(new_n352_));
  INV_X1    g151(.A(G15gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n350_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G71gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n352_), .A2(new_n356_), .A3(G99gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(G99gat), .B1(new_n352_), .B2(new_n356_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT24), .ZN(new_n362_));
  INV_X1    g161(.A(G169gat), .ZN(new_n363_));
  INV_X1    g162(.A(G176gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  MUX2_X1   g164(.A(KEYINPUT24), .B(new_n362_), .S(new_n365_), .Z(new_n366_));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT23), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT26), .B(G190gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n369_), .A2(KEYINPUT78), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT25), .B(G183gat), .ZN(new_n371_));
  INV_X1    g170(.A(G190gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT78), .B1(new_n372_), .B2(KEYINPUT26), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n366_), .B(new_n368_), .C1(new_n370_), .C2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G183gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n372_), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n368_), .A2(new_n377_), .B1(G169gat), .B2(G176gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n363_), .B1(KEYINPUT79), .B2(KEYINPUT22), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(KEYINPUT80), .B2(KEYINPUT22), .ZN(new_n380_));
  NAND2_X1  g179(.A1(KEYINPUT80), .A2(G169gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(KEYINPUT79), .A3(KEYINPUT22), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n382_), .A3(new_n364_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n375_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT30), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n375_), .A2(new_n384_), .A3(KEYINPUT30), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n360_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G127gat), .B(G134gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G113gat), .B(G120gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n387_), .A2(new_n360_), .A3(new_n388_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n393_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n394_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n396_), .B1(new_n397_), .B2(new_n389_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT81), .B(G43gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT31), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n395_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT98), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT96), .B(G85gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT0), .B(G57gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT95), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT1), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT82), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT83), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n419_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n417_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G141gat), .ZN(new_n426_));
  INV_X1    g225(.A(G148gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G141gat), .A2(G148gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n422_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n420_), .A2(KEYINPUT83), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n418_), .A2(KEYINPUT82), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n419_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n429_), .A2(KEYINPUT84), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT2), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n442_));
  OAI22_X1  g241(.A1(new_n442_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n439_), .A2(new_n441_), .A3(new_n443_), .A4(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n437_), .A2(new_n415_), .A3(new_n445_), .ZN(new_n446_));
  AOI211_X1 g245(.A(new_n414_), .B(new_n393_), .C1(new_n431_), .C2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n431_), .A2(new_n446_), .A3(new_n393_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT4), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n431_), .A2(new_n446_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n451_), .A2(KEYINPUT95), .A3(new_n452_), .A4(new_n396_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n413_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n448_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n393_), .B1(new_n431_), .B2(new_n446_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n412_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n411_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n415_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n445_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n430_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n463_), .B1(new_n437_), .B2(new_n417_), .ZN(new_n464_));
  OAI211_X1 g263(.A(KEYINPUT95), .B(new_n396_), .C1(new_n462_), .C2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(KEYINPUT4), .A3(new_n448_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n412_), .B1(new_n466_), .B2(new_n453_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n458_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n467_), .A2(new_n410_), .A3(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n405_), .B1(new_n459_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n455_), .A2(new_n411_), .A3(new_n458_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n410_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(KEYINPUT98), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n404_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G8gat), .B(G36gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT18), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT21), .ZN(new_n481_));
  INV_X1    g280(.A(G197gat), .ZN(new_n482_));
  INV_X1    g281(.A(G204gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT87), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G204gat), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n482_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(G197gat), .A2(G204gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n481_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G218gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G211gat), .ZN(new_n491_));
  INV_X1    g290(.A(G211gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G218gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n484_), .A2(new_n486_), .A3(new_n482_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n481_), .B1(G197gat), .B2(G204gat), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n489_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n488_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT87), .B(G204gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n499_), .B1(new_n500_), .B2(new_n482_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(KEYINPUT21), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n484_), .A2(new_n486_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n488_), .B1(new_n505_), .B2(G197gat), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n481_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT88), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n498_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT89), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n503_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n506_), .A2(KEYINPUT88), .A3(new_n507_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n512_), .A2(new_n513_), .B1(new_n489_), .B2(new_n497_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT89), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n511_), .A2(new_n515_), .A3(new_n385_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G226gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT19), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT20), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT22), .B(G169gat), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n521_), .A2(KEYINPUT93), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(KEYINPUT93), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n364_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n369_), .A2(new_n371_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n525_), .A2(new_n368_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n524_), .A2(new_n378_), .B1(new_n526_), .B2(new_n366_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n520_), .B1(new_n527_), .B2(new_n514_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n516_), .A2(new_n519_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n385_), .ZN(new_n530_));
  AOI221_X4 g329(.A(new_n510_), .B1(new_n489_), .B2(new_n497_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n512_), .A2(new_n513_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT89), .B1(new_n532_), .B2(new_n498_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n530_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n527_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n520_), .B1(new_n535_), .B2(new_n509_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n519_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n480_), .B1(new_n529_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n516_), .A2(new_n519_), .A3(new_n528_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT20), .B1(new_n527_), .B2(new_n514_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n511_), .A2(new_n515_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n530_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n479_), .B(new_n540_), .C1(new_n543_), .C2(new_n519_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n538_), .A2(new_n539_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT27), .ZN(new_n546_));
  INV_X1    g345(.A(new_n537_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n547_), .A2(KEYINPUT94), .A3(new_n479_), .A4(new_n540_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n545_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n544_), .A2(KEYINPUT27), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n534_), .A2(new_n519_), .A3(new_n536_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n519_), .B1(new_n516_), .B2(new_n528_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  AOI211_X1 g353(.A(KEYINPUT97), .B(new_n519_), .C1(new_n516_), .C2(new_n528_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n480_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT29), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n431_), .B2(new_n446_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G228gat), .A2(G233gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT86), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n560_), .B2(new_n514_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G78gat), .B(G106gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT90), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(new_n569_), .A3(new_n566_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n451_), .B2(KEYINPUT29), .ZN(new_n576_));
  XOR2_X1   g375(.A(G22gat), .B(G50gat), .Z(new_n577_));
  INV_X1    g376(.A(new_n575_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n431_), .A2(new_n446_), .A3(new_n559_), .A4(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n576_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n577_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n565_), .A2(KEYINPUT91), .A3(new_n569_), .A4(new_n566_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n574_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n451_), .A2(KEYINPUT29), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n562_), .B1(new_n587_), .B2(new_n509_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n531_), .A2(new_n533_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n589_), .B2(new_n564_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n586_), .B1(new_n590_), .B2(new_n569_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n567_), .A2(KEYINPUT92), .A3(new_n570_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n582_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .A4(new_n573_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n585_), .A2(new_n594_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n475_), .A2(new_n558_), .A3(new_n595_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n549_), .A2(new_n595_), .A3(new_n557_), .A4(new_n474_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n594_), .A2(new_n585_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n600_), .A2(KEYINPUT99), .A3(new_n549_), .A4(new_n557_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n595_), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT32), .B(new_n479_), .C1(new_n554_), .C2(new_n555_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n471_), .A2(new_n472_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n479_), .A2(KEYINPUT32), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n547_), .A2(new_n540_), .A3(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  OAI211_X1 g406(.A(KEYINPUT33), .B(new_n410_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n456_), .A2(new_n457_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n410_), .B1(new_n610_), .B2(new_n413_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n466_), .A2(new_n412_), .A3(new_n453_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n608_), .B1(new_n459_), .B2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n602_), .B1(new_n607_), .B2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n599_), .A2(new_n601_), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n596_), .B1(new_n617_), .B2(new_n403_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n241_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n619_), .A2(new_n300_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G229gat), .A2(G233gat), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n242_), .A2(new_n300_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n619_), .B(new_n300_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n621_), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n622_), .A2(new_n623_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G169gat), .B(G197gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT77), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n626_), .A2(new_n629_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n618_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n349_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n474_), .A2(G1gat), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT100), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n640_), .A3(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n347_), .A2(new_n633_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n312_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n266_), .B(KEYINPUT101), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n618_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT102), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n474_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n639_), .A2(KEYINPUT38), .A3(new_n641_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n644_), .A2(new_n653_), .A3(new_n654_), .ZN(G1324gat));
  NAND3_X1  g454(.A1(new_n636_), .A2(new_n296_), .A3(new_n558_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n650_), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT39), .B(new_n296_), .C1(new_n657_), .C2(new_n558_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n558_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(G8gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n656_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g462(.A1(new_n636_), .A2(new_n353_), .A3(new_n404_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n651_), .A2(new_n404_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n665_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT41), .B1(new_n665_), .B2(G15gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n664_), .B1(new_n666_), .B2(new_n667_), .ZN(G1326gat));
  INV_X1    g467(.A(G22gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n636_), .A2(new_n669_), .A3(new_n595_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G22gat), .B1(new_n652_), .B2(new_n602_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(KEYINPUT42), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(KEYINPUT42), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(G1327gat));
  INV_X1    g473(.A(new_n347_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n267_), .A2(new_n312_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n635_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n474_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n273_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n271_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n266_), .A2(new_n269_), .A3(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n617_), .A2(new_n403_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n596_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT104), .B(KEYINPUT43), .C1(new_n688_), .C2(KEYINPUT103), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n645_), .A2(new_n311_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n545_), .A2(new_n548_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n614_), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n694_), .A2(new_n602_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n404_), .B1(new_n695_), .B2(new_n601_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n274_), .B1(new_n696_), .B2(new_n596_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n691_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n691_), .B1(new_n618_), .B2(new_n685_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n689_), .B(new_n690_), .C1(new_n699_), .C2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT104), .B1(new_n688_), .B2(KEYINPUT103), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n701_), .A3(new_n700_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n707_), .A2(KEYINPUT44), .A3(new_n689_), .A4(new_n690_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n680_), .A2(G29gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n681_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  NAND3_X1  g511(.A1(new_n705_), .A2(new_n558_), .A3(new_n708_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G36gat), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n558_), .A2(KEYINPUT105), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n558_), .A2(KEYINPUT105), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n678_), .A2(G36gat), .A3(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT45), .Z(new_n720_));
  NAND2_X1  g519(.A1(new_n714_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n714_), .A2(KEYINPUT46), .A3(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  XOR2_X1   g524(.A(KEYINPUT106), .B(G43gat), .Z(new_n726_));
  OAI21_X1  g525(.A(new_n726_), .B1(new_n678_), .B2(new_n403_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n404_), .A2(G43gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n709_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g529(.A(G50gat), .B1(new_n679_), .B2(new_n595_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n595_), .A2(G50gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n710_), .B2(new_n732_), .ZN(G1331gat));
  NAND2_X1  g532(.A1(new_n675_), .A2(new_n634_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n734_), .A2(new_n618_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(new_n313_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G57gat), .B1(new_n736_), .B2(new_n680_), .ZN(new_n737_));
  NOR4_X1   g536(.A1(new_n734_), .A2(new_n618_), .A3(new_n312_), .A4(new_n648_), .ZN(new_n738_));
  INV_X1    g537(.A(G57gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n680_), .B2(KEYINPUT107), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(KEYINPUT107), .B2(new_n739_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n737_), .B1(new_n738_), .B2(new_n741_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  INV_X1    g542(.A(new_n718_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n738_), .B2(new_n744_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT48), .Z(new_n746_));
  NAND3_X1  g545(.A1(new_n736_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1333gat));
  NAND3_X1  g547(.A1(new_n736_), .A2(new_n355_), .A3(new_n404_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n738_), .A2(new_n404_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(G71gat), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT49), .B(new_n355_), .C1(new_n738_), .C2(new_n404_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT108), .Z(G1334gat));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n738_), .B2(new_n595_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT50), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n736_), .A2(new_n756_), .A3(new_n595_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n734_), .A2(new_n311_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n689_), .C1(new_n699_), .C2(new_n702_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n707_), .A2(KEYINPUT110), .A3(new_n689_), .A4(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n680_), .A2(G85gat), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT111), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(G85gat), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n734_), .A2(new_n618_), .A3(new_n676_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT109), .Z(new_n772_));
  OAI21_X1  g571(.A(new_n770_), .B1(new_n772_), .B2(new_n474_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n769_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n769_), .A2(new_n773_), .A3(KEYINPUT112), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1336gat));
  AOI21_X1  g577(.A(new_n718_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n558_), .A2(new_n207_), .ZN(new_n780_));
  OAI22_X1  g579(.A1(new_n779_), .A2(new_n207_), .B1(new_n772_), .B2(new_n780_), .ZN(G1337gat));
  AOI21_X1  g580(.A(new_n403_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n404_), .A2(new_n222_), .ZN(new_n783_));
  OAI22_X1  g582(.A1(new_n782_), .A2(new_n216_), .B1(new_n772_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  OAI221_X1 g586(.A(new_n785_), .B1(new_n772_), .B2(new_n783_), .C1(new_n782_), .C2(new_n216_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1338gat));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n790_), .B(G106gat), .C1(new_n762_), .C2(new_n602_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n707_), .A2(new_n595_), .A3(new_n689_), .A4(new_n761_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n790_), .B1(new_n793_), .B2(G106gat), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n595_), .A2(new_n217_), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n792_), .A2(new_n794_), .B1(new_n772_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  OAI221_X1 g598(.A(new_n797_), .B1(new_n772_), .B2(new_n795_), .C1(new_n792_), .C2(new_n794_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1339gat));
  INV_X1    g600(.A(new_n558_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n602_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n404_), .A2(new_n680_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n633_), .A2(new_n337_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n314_), .B(new_n316_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n318_), .A2(KEYINPUT68), .A3(KEYINPUT12), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n328_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT115), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n324_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT12), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n321_), .B1(new_n325_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n314_), .A2(new_n316_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n818_), .A2(KEYINPUT55), .A3(new_n323_), .A4(new_n322_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n328_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n812_), .A2(new_n814_), .A3(new_n819_), .A4(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(KEYINPUT56), .A3(new_n335_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n822_), .B2(new_n335_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(KEYINPUT116), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n826_), .B(KEYINPUT56), .C1(new_n822_), .C2(new_n335_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n808_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n623_), .A2(new_n620_), .A3(new_n625_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n629_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n624_), .A2(new_n621_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT117), .Z(new_n833_));
  AND2_X1   g632(.A1(new_n631_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n343_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n267_), .B1(new_n828_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT57), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n834_), .A2(new_n337_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n823_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n838_), .B(KEYINPUT58), .C1(new_n839_), .C2(new_n824_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n840_), .A2(KEYINPUT119), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n838_), .B1(new_n839_), .B2(new_n824_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n685_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n840_), .A2(KEYINPUT119), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n837_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n836_), .A2(KEYINPUT57), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n312_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n347_), .A2(new_n311_), .A3(new_n685_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n634_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n348_), .A2(KEYINPUT54), .A3(new_n633_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n807_), .B1(new_n849_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n852_), .A2(new_n853_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n836_), .B2(KEYINPUT57), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860_));
  INV_X1    g659(.A(new_n821_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n317_), .A2(new_n322_), .A3(new_n319_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n820_), .B1(new_n862_), .B2(new_n328_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n814_), .A2(new_n819_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n336_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n826_), .B1(new_n866_), .B2(KEYINPUT56), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n824_), .A2(KEYINPUT116), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n823_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n869_), .A2(new_n808_), .B1(new_n343_), .B2(new_n834_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT118), .B(new_n860_), .C1(new_n870_), .C2(new_n267_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n859_), .A2(new_n871_), .A3(new_n837_), .A4(new_n846_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n857_), .B1(new_n872_), .B2(new_n312_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n805_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n856_), .B(new_n633_), .C1(new_n875_), .C2(new_n806_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G113gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n872_), .A2(new_n312_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n854_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n805_), .ZN(new_n880_));
  OR3_X1    g679(.A1(new_n880_), .A2(G113gat), .A3(new_n634_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n881_), .ZN(G1340gat));
  OAI211_X1 g681(.A(new_n856_), .B(new_n675_), .C1(new_n875_), .C2(new_n806_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G120gat), .ZN(new_n884_));
  INV_X1    g683(.A(G120gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n347_), .B2(KEYINPUT60), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n875_), .B(new_n886_), .C1(KEYINPUT60), .C2(new_n885_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n887_), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT120), .B(new_n889_), .C1(new_n880_), .C2(new_n312_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n873_), .A2(new_n312_), .A3(new_n874_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(G127gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n855_), .B1(new_n880_), .B2(KEYINPUT59), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n312_), .A2(new_n889_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n890_), .A2(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1342gat));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897_));
  INV_X1    g696(.A(G134gat), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n897_), .B(new_n898_), .C1(new_n880_), .C2(new_n647_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n873_), .A2(new_n647_), .A3(new_n874_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT121), .B1(new_n900_), .B2(G134gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n685_), .A2(new_n898_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT122), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n899_), .A2(new_n901_), .B1(new_n894_), .B2(new_n903_), .ZN(G1343gat));
  NAND4_X1  g703(.A1(new_n718_), .A2(new_n595_), .A3(new_n680_), .A4(new_n403_), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(KEYINPUT123), .Z(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(new_n878_), .B2(new_n854_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n633_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT124), .B(G141gat), .Z(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1344gat));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n675_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g711(.A1(new_n907_), .A2(new_n311_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT61), .B(G155gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1346gat));
  INV_X1    g714(.A(G162gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n907_), .B2(new_n274_), .ZN(new_n917_));
  NOR4_X1   g716(.A1(new_n873_), .A2(G162gat), .A3(new_n647_), .A4(new_n906_), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT125), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n907_), .A2(new_n916_), .A3(new_n648_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n873_), .A2(new_n685_), .A3(new_n906_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n920_), .B(new_n921_), .C1(new_n922_), .C2(new_n916_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n919_), .A2(new_n923_), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n718_), .A2(new_n475_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n602_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n849_), .B2(new_n854_), .ZN(new_n927_));
  AOI211_X1 g726(.A(KEYINPUT62), .B(new_n363_), .C1(new_n927_), .C2(new_n633_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n633_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(G169gat), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n927_), .B(new_n633_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n928_), .B1(new_n931_), .B2(new_n932_), .ZN(G1348gat));
  AOI21_X1  g732(.A(G176gat), .B1(new_n927_), .B2(new_n675_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n675_), .A2(new_n925_), .A3(G176gat), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n873_), .A2(new_n595_), .A3(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n935_), .A2(new_n936_), .A3(new_n939_), .ZN(new_n940_));
  OAI21_X1  g739(.A(KEYINPUT126), .B1(new_n934_), .B2(new_n938_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1349gat));
  INV_X1    g741(.A(new_n927_), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n943_), .A2(new_n371_), .A3(new_n312_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n879_), .A2(new_n602_), .A3(new_n311_), .A4(new_n925_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n945_), .B2(new_n376_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n943_), .B2(new_n685_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n927_), .A2(new_n369_), .A3(new_n648_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1351gat));
  NOR4_X1   g748(.A1(new_n718_), .A2(new_n602_), .A3(new_n680_), .A4(new_n404_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n879_), .A2(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(G197gat), .B1(new_n952_), .B2(new_n633_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n951_), .A2(new_n482_), .A3(new_n634_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1352gat));
  NOR3_X1   g754(.A1(new_n951_), .A2(new_n500_), .A3(new_n347_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n952_), .A2(new_n675_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n956_), .B1(new_n483_), .B2(new_n957_), .ZN(G1353gat));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n959_));
  AND3_X1   g758(.A1(new_n959_), .A2(new_n492_), .A3(KEYINPUT127), .ZN(new_n960_));
  AOI211_X1 g759(.A(new_n960_), .B(new_n312_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n879_), .A2(new_n950_), .A3(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(KEYINPUT127), .B1(new_n959_), .B2(new_n492_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n962_), .B(new_n963_), .ZN(G1354gat));
  OAI21_X1  g763(.A(G218gat), .B1(new_n951_), .B2(new_n685_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n648_), .A2(new_n490_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n951_), .B2(new_n966_), .ZN(G1355gat));
endmodule


