//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n207_), .A2(new_n210_), .A3(new_n211_), .A4(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT8), .B1(new_n217_), .B2(KEYINPUT65), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n213_), .B(new_n217_), .C1(KEYINPUT65), .C2(KEYINPUT8), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT10), .B(G99gat), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n210_), .B(new_n211_), .C1(new_n223_), .C2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT9), .ZN(new_n225_));
  OR2_X1    g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(new_n226_), .B2(new_n214_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n214_), .A2(new_n225_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT64), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT9), .B1(new_n215_), .B2(new_n216_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n228_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n224_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT66), .B1(new_n222_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n224_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n227_), .A2(KEYINPUT64), .A3(new_n229_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n232_), .B1(new_n231_), .B2(new_n228_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT67), .B(G71gat), .ZN(new_n242_));
  INV_X1    g041(.A(G78gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(G71gat), .ZN(new_n246_));
  INV_X1    g045(.A(G71gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(KEYINPUT67), .ZN(new_n248_));
  OAI21_X1  g047(.A(G78gat), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G57gat), .B(G64gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(KEYINPUT11), .A3(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G57gat), .B(G64gat), .Z(new_n253_));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(KEYINPUT11), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n255_), .A2(new_n249_), .A3(new_n256_), .A4(new_n244_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n252_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n235_), .A2(new_n241_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n262_));
  OAI211_X1 g061(.A(KEYINPUT68), .B(new_n203_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n235_), .A2(new_n241_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n220_), .A2(new_n221_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n258_), .B1(new_n266_), .B2(new_n239_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n265_), .A2(new_n258_), .B1(new_n267_), .B2(KEYINPUT12), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n260_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n202_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT68), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n203_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n264_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G120gat), .B(G148gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(G176gat), .B(G204gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n274_), .B(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n282_));
  NOR2_X1   g081(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n281_), .A2(new_n282_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT15), .ZN(new_n290_));
  INV_X1    g089(.A(G29gat), .ZN(new_n291_));
  INV_X1    g090(.A(G36gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G29gat), .A2(G36gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G43gat), .ZN(new_n296_));
  INV_X1    g095(.A(G43gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n297_), .A3(new_n294_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(G50gat), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(G50gat), .B1(new_n296_), .B2(new_n298_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n290_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(KEYINPUT15), .A3(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G1gat), .B(G8gat), .Z(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G15gat), .B(G22gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n309_));
  INV_X1    g108(.A(G1gat), .ZN(new_n310_));
  INV_X1    g109(.A(G8gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT14), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(new_n309_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n309_), .B1(new_n308_), .B2(new_n312_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n307_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n306_), .A3(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n305_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G229gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n300_), .A2(new_n301_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n319_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n323_), .B1(new_n319_), .B2(new_n324_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n321_), .B(new_n322_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n319_), .A2(new_n324_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n319_), .A2(new_n324_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT77), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n331_), .B2(new_n325_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n328_), .B1(new_n332_), .B2(new_n322_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G113gat), .B(G141gat), .ZN(new_n336_));
  INV_X1    g135(.A(G169gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(G197gat), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n333_), .A2(new_n334_), .A3(new_n339_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n265_), .A2(new_n324_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n305_), .B1(new_n234_), .B2(new_n222_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G232gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT34), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(KEYINPUT35), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(KEYINPUT35), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n349_), .A2(KEYINPUT35), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n345_), .A2(new_n351_), .A3(new_n352_), .A4(new_n346_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT72), .B(G190gat), .ZN(new_n355_));
  INV_X1    g154(.A(G218gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G134gat), .B(G162gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(KEYINPUT36), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(KEYINPUT36), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n354_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n350_), .A2(new_n361_), .A3(new_n353_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(KEYINPUT74), .ZN(new_n370_));
  INV_X1    g169(.A(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT73), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n354_), .A2(new_n373_), .A3(new_n362_), .A4(new_n363_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n370_), .A2(new_n372_), .A3(new_n374_), .A4(new_n368_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n369_), .B1(new_n375_), .B2(KEYINPUT37), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n289_), .A2(new_n344_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G113gat), .ZN(new_n382_));
  INV_X1    g181(.A(G120gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n381_), .A2(G113gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(G113gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(G120gat), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(G141gat), .A2(G148gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT3), .Z(new_n394_));
  NAND2_X1  g193(.A1(G141gat), .A2(G148gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n395_), .B(KEYINPUT2), .Z(new_n396_));
  OAI21_X1  g195(.A(new_n392_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n392_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n390_), .A2(KEYINPUT1), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n395_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n389_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT95), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n388_), .A2(new_n405_), .A3(new_n402_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n380_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n406_), .A2(new_n380_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n379_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n403_), .B(new_n388_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n378_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G1gat), .B(G29gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G57gat), .B(G85gat), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n416_), .B(new_n417_), .Z(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT97), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n412_), .B2(new_n418_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n413_), .A2(new_n421_), .A3(new_n419_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G22gat), .B(G50gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G211gat), .B(G218gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(G197gat), .B(G204gat), .Z(new_n430_));
  OAI21_X1  g229(.A(new_n429_), .B1(new_n430_), .B2(KEYINPUT21), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(KEYINPUT21), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n434_), .B1(new_n403_), .B2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT86), .B(G233gat), .Z(new_n437_));
  AND2_X1   g236(.A1(new_n437_), .A2(G228gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G78gat), .B(G106gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n434_), .B(new_n440_), .C1(new_n403_), .C2(new_n435_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n402_), .A2(KEYINPUT29), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n446_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .A4(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT87), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n447_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n428_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n455_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(new_n427_), .A3(new_n453_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT80), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(G169gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n337_), .A2(KEYINPUT80), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT22), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT81), .ZN(new_n467_));
  AOI21_X1  g266(.A(G176gat), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  OAI221_X1 g267(.A(new_n468_), .B1(new_n467_), .B2(new_n466_), .C1(KEYINPUT22), .C2(new_n337_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G169gat), .A2(G176gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT82), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G183gat), .A2(G190gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT23), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT79), .B(G183gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n474_), .B1(G190gat), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n469_), .A2(new_n477_), .A3(new_n470_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n472_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n480_));
  INV_X1    g279(.A(G176gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n337_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(KEYINPUT24), .A3(new_n470_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n474_), .B(new_n483_), .C1(KEYINPUT24), .C2(new_n482_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT26), .B(G190gat), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n475_), .A2(KEYINPUT25), .ZN(new_n486_));
  OR2_X1    g285(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n479_), .A2(new_n480_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n480_), .B1(new_n479_), .B2(new_n489_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n462_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n479_), .A2(new_n489_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT30), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(new_n490_), .A3(new_n461_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G15gat), .B(G43gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G227gat), .A2(G233gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n493_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G71gat), .B(G99gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n388_), .B(new_n504_), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n502_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n493_), .A2(new_n496_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n499_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n505_), .B1(new_n509_), .B2(new_n501_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n460_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n506_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n509_), .A2(new_n505_), .A3(new_n501_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n459_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n426_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT27), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT22), .B(G169gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT91), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n481_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n474_), .B1(G183gat), .B2(G190gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n470_), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT25), .B(G183gat), .Z(new_n524_));
  NOR2_X1   g323(.A1(new_n485_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n484_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n434_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(KEYINPUT20), .B(new_n527_), .C1(new_n494_), .C2(new_n434_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT89), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G226gat), .A2(G233gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(new_n531_), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT90), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G8gat), .B(G36gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(G64gat), .B(G92gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n494_), .A2(new_n434_), .ZN(new_n541_));
  OR3_X1    g340(.A1(new_n523_), .A2(new_n434_), .A3(new_n526_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(KEYINPUT20), .A4(new_n532_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n534_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n540_), .B1(new_n534_), .B2(new_n543_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n516_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n526_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n521_), .A2(new_n433_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n494_), .B2(new_n434_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n532_), .B1(new_n549_), .B2(KEYINPUT20), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n528_), .A2(new_n533_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n539_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n534_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(KEYINPUT27), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n534_), .A2(new_n543_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n539_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(KEYINPUT94), .A3(new_n553_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n378_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n410_), .A2(new_n379_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n418_), .A3(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n420_), .B(KEYINPUT33), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n558_), .A2(new_n561_), .A3(new_n564_), .A4(new_n565_), .ZN(new_n566_));
  OAI211_X1 g365(.A(KEYINPUT32), .B(new_n540_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n540_), .A2(KEYINPUT32), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n534_), .A2(new_n569_), .A3(new_n543_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n423_), .A2(new_n570_), .A3(new_n424_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT98), .B1(new_n568_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n426_), .A2(new_n573_), .A3(new_n567_), .A4(new_n570_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n566_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n507_), .A2(new_n510_), .A3(new_n459_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n515_), .A2(new_n556_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n258_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(new_n319_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G127gat), .B(G155gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(G183gat), .B(G211gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n580_), .A2(KEYINPUT17), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n585_), .B(KEYINPUT17), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n587_), .B1(new_n580_), .B2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n577_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n377_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT99), .Z(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(new_n310_), .A3(new_n426_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT38), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n365_), .A2(new_n371_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n577_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n590_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n287_), .A2(new_n344_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G1gat), .B1(new_n602_), .B2(new_n425_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n594_), .A2(new_n595_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n596_), .A2(new_n603_), .A3(new_n604_), .ZN(G1324gat));
  NAND3_X1  g404(.A1(new_n593_), .A2(new_n311_), .A3(new_n555_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G8gat), .B1(new_n602_), .B2(new_n556_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(KEYINPUT39), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(KEYINPUT39), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n606_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT40), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n606_), .B(new_n612_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1325gat));
  INV_X1    g415(.A(G15gat), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n507_), .A2(new_n510_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n601_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT41), .ZN(new_n621_));
  INV_X1    g420(.A(new_n592_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(G1326gat));
  NAND2_X1  g423(.A1(new_n601_), .A2(new_n459_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT42), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n625_), .A2(new_n626_), .A3(G22gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n625_), .B2(G22gat), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n460_), .A2(G22gat), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT102), .Z(new_n630_));
  OAI22_X1  g429(.A1(new_n627_), .A2(new_n628_), .B1(new_n592_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1327gat));
  NAND2_X1  g432(.A1(new_n600_), .A2(new_n590_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n597_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n577_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n291_), .A3(new_n426_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n376_), .B2(KEYINPUT104), .ZN(new_n640_));
  INV_X1    g439(.A(new_n376_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(new_n577_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n575_), .A2(new_n576_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n514_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n459_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n556_), .B(new_n425_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n640_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(new_n376_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n634_), .B1(new_n642_), .B2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n638_), .B1(new_n650_), .B2(KEYINPUT105), .ZN(new_n651_));
  INV_X1    g450(.A(new_n634_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n577_), .A2(new_n641_), .A3(new_n640_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n648_), .B1(new_n647_), .B2(new_n376_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n652_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(KEYINPUT44), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n425_), .B1(new_n651_), .B2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n637_), .B1(new_n658_), .B2(new_n291_), .ZN(G1328gat));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT107), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n636_), .A2(new_n292_), .A3(new_n555_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT45), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n556_), .B1(new_n651_), .B2(new_n657_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n661_), .B(new_n663_), .C1(new_n664_), .C2(new_n292_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT107), .B1(new_n660_), .B2(KEYINPUT106), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT108), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n665_), .B(new_n667_), .ZN(G1329gat));
  INV_X1    g467(.A(KEYINPUT47), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT44), .B1(new_n655_), .B2(new_n656_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n650_), .A2(KEYINPUT105), .A3(new_n638_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n619_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G43gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n636_), .A2(new_n297_), .A3(new_n619_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n669_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n618_), .B1(new_n651_), .B2(new_n657_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n669_), .B(new_n674_), .C1(new_n676_), .C2(new_n297_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n675_), .A2(new_n678_), .ZN(G1330gat));
  OAI21_X1  g478(.A(new_n459_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT109), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n459_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n681_), .A2(G50gat), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n636_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n460_), .A2(G50gat), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT110), .Z(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(new_n685_), .B2(new_n687_), .ZN(G1331gat));
  OR2_X1    g487(.A1(new_n285_), .A2(new_n286_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n343_), .A2(new_n590_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n641_), .A2(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n577_), .A2(new_n689_), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G57gat), .B1(new_n692_), .B2(new_n426_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n598_), .A2(new_n289_), .A3(new_n690_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(G57gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n695_), .B2(new_n426_), .ZN(G1332gat));
  INV_X1    g495(.A(G64gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n694_), .B2(new_n555_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT48), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n692_), .A2(new_n697_), .A3(new_n555_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1333gat));
  NAND3_X1  g500(.A1(new_n692_), .A2(new_n247_), .A3(new_n619_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n694_), .A2(new_n619_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G71gat), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(KEYINPUT49), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(KEYINPUT49), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT111), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n709_), .B(new_n702_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1334gat));
  AOI21_X1  g510(.A(new_n243_), .B1(new_n694_), .B2(new_n459_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT50), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n692_), .A2(new_n243_), .A3(new_n459_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n599_), .A2(new_n343_), .ZN(new_n716_));
  AND4_X1   g515(.A1(new_n597_), .A2(new_n647_), .A3(new_n289_), .A4(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G85gat), .B1(new_n717_), .B2(new_n426_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n642_), .A2(new_n649_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n287_), .A2(new_n716_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT112), .Z(new_n721_));
  AND3_X1   g520(.A1(new_n719_), .A2(G85gat), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n718_), .B1(new_n722_), .B2(new_n426_), .ZN(G1336gat));
  AOI21_X1  g522(.A(G92gat), .B1(new_n717_), .B2(new_n555_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n719_), .A2(new_n555_), .A3(new_n721_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(G92gat), .ZN(G1337gat));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n719_), .A2(new_n619_), .A3(new_n721_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n618_), .A2(new_n223_), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n728_), .A2(G99gat), .B1(new_n717_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n731_));
  AND4_X1   g530(.A1(new_n727_), .A2(new_n730_), .A3(new_n731_), .A4(KEYINPUT51), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT51), .B1(new_n730_), .B2(new_n731_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n730_), .A2(new_n727_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(G1338gat));
  NAND3_X1  g534(.A1(new_n717_), .A2(new_n206_), .A3(new_n459_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n719_), .A2(new_n459_), .A3(new_n721_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(G106gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G106gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g541(.A1(new_n555_), .A2(new_n425_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n645_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n202_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n271_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n268_), .A2(KEYINPUT55), .A3(new_n202_), .A4(new_n270_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n280_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT56), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n274_), .A2(new_n280_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n321_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(G229gat), .A3(G233gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n332_), .A2(new_n322_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  MUX2_X1   g554(.A(new_n333_), .B(new_n755_), .S(new_n339_), .Z(new_n756_));
  NOR2_X1   g555(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n750_), .A2(new_n751_), .A3(new_n756_), .A4(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n747_), .A2(new_n748_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT56), .B1(new_n760_), .B2(new_n279_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n762_), .B(new_n280_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n751_), .B(new_n756_), .C1(new_n761_), .C2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n757_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n759_), .A2(new_n765_), .A3(new_n376_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT57), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n274_), .A2(new_n280_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n274_), .A2(new_n280_), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n279_), .B(new_n264_), .C1(new_n273_), .C2(new_n272_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n756_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n769_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n767_), .B1(new_n773_), .B2(new_n635_), .ZN(new_n774_));
  AOI211_X1 g573(.A(KEYINPUT57), .B(new_n597_), .C1(new_n769_), .C2(new_n772_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n766_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n766_), .B(KEYINPUT116), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n590_), .A3(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n691_), .A2(new_n287_), .A3(KEYINPUT54), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n376_), .A2(new_n590_), .A3(new_n343_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n689_), .B2(new_n783_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n781_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n744_), .B1(new_n780_), .B2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(G113gat), .B1(new_n786_), .B2(new_n343_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n780_), .A2(new_n785_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n744_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(KEYINPUT117), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n744_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT59), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n776_), .A2(new_n590_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n781_), .A2(new_n784_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n791_), .A2(new_n343_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n787_), .B1(new_n800_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n791_), .A2(new_n802_), .A3(new_n289_), .A4(new_n798_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT59), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n289_), .B(new_n798_), .C1(new_n786_), .C2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT118), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n803_), .A2(G120gat), .A3(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n383_), .B1(new_n689_), .B2(KEYINPUT60), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n786_), .B(new_n808_), .C1(KEYINPUT60), .C2(new_n383_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n807_), .A2(KEYINPUT119), .A3(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1341gat));
  AOI21_X1  g613(.A(G127gat), .B1(new_n786_), .B2(new_n599_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n791_), .A2(G127gat), .A3(new_n798_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n817_), .B2(new_n599_), .ZN(G1342gat));
  AOI21_X1  g617(.A(G134gat), .B1(new_n786_), .B2(new_n597_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n791_), .A2(G134gat), .A3(new_n798_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n821_), .B2(new_n376_), .ZN(G1343gat));
  AOI21_X1  g621(.A(new_n514_), .B1(new_n780_), .B2(new_n785_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n743_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT120), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(new_n826_), .A3(new_n743_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n343_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n289_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n599_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT61), .B(G155gat), .Z(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT121), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n833_), .B(new_n835_), .ZN(G1346gat));
  AOI21_X1  g635(.A(G162gat), .B1(new_n828_), .B2(new_n597_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n828_), .A2(G162gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n376_), .B2(new_n838_), .ZN(G1347gat));
  NOR2_X1   g638(.A1(new_n556_), .A2(new_n426_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n619_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n460_), .B(new_n842_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n843_));
  OAI21_X1  g642(.A(G169gat), .B1(new_n843_), .B2(new_n344_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n843_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n518_), .A3(new_n343_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1348gat));
  NAND2_X1  g648(.A1(new_n788_), .A2(new_n460_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AND4_X1   g650(.A1(G176gat), .A2(new_n851_), .A3(new_n289_), .A4(new_n842_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n481_), .B1(new_n843_), .B2(new_n689_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n854_), .A2(KEYINPUT123), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(KEYINPUT123), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n852_), .B1(new_n855_), .B2(new_n856_), .ZN(G1349gat));
  NAND3_X1  g656(.A1(new_n851_), .A2(new_n599_), .A3(new_n842_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n475_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n599_), .A2(new_n524_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n858_), .A2(new_n859_), .B1(new_n847_), .B2(new_n860_), .ZN(G1350gat));
  NOR3_X1   g660(.A1(new_n843_), .A2(new_n635_), .A3(new_n485_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n847_), .A2(new_n376_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(G190gat), .B2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT124), .ZN(G1351gat));
  NAND2_X1  g664(.A1(new_n823_), .A2(new_n840_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n343_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n289_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(G204gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT125), .B(G204gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n870_), .B2(new_n873_), .ZN(G1353gat));
  AOI21_X1  g673(.A(new_n590_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n866_), .A2(KEYINPUT126), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT126), .B1(new_n866_), .B2(new_n876_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1354gat));
  NAND3_X1  g680(.A1(new_n867_), .A2(KEYINPUT127), .A3(new_n597_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT127), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n866_), .B2(new_n635_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n882_), .A2(new_n356_), .A3(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n867_), .A2(G218gat), .A3(new_n376_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1355gat));
endmodule


