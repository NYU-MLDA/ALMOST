//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n977_,
    new_n978_, new_n979_, new_n981_, new_n982_, new_n984_, new_n985_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1001_, new_n1002_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G78gat), .Z(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n204_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209_));
  INV_X1    g008(.A(G1gat), .ZN(new_n210_));
  INV_X1    g009(.A(G8gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n208_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G231gat), .A2(G233gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G127gat), .B(G155gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT16), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(G211gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n223_), .B(new_n224_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT80), .ZN(new_n228_));
  OAI211_X1 g027(.A(KEYINPUT79), .B(new_n226_), .C1(new_n228_), .C2(new_n218_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n226_), .A2(KEYINPUT79), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT10), .B(G99gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(G106gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G85gat), .A2(G92gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n235_), .A2(KEYINPUT9), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT6), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT6), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(G99gat), .A3(G106gat), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n236_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n242_));
  INV_X1    g041(.A(G85gat), .ZN(new_n243_));
  INV_X1    g042(.A(G92gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n242_), .A2(new_n245_), .A3(new_n235_), .A4(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n234_), .A2(new_n241_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT8), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G85gat), .B(G92gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT65), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n245_), .A2(new_n252_), .A3(new_n235_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n238_), .A2(new_n240_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G99gat), .A2(G106gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT7), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n256_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n249_), .B1(new_n254_), .B2(new_n260_), .ZN(new_n261_));
  AND4_X1   g060(.A1(new_n249_), .A2(new_n260_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n248_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(G29gat), .A2(G36gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G29gat), .A2(G36gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(G43gat), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G29gat), .ZN(new_n267_));
  INV_X1    g066(.A(G36gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G43gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G29gat), .A2(G36gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n266_), .A2(new_n272_), .A3(G50gat), .ZN(new_n273_));
  AOI21_X1  g072(.A(G50gat), .B1(new_n266_), .B2(new_n272_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT71), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G50gat), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n264_), .A2(new_n265_), .A3(G43gat), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n270_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n266_), .A2(new_n272_), .A3(G50gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n275_), .A2(KEYINPUT15), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT15), .B1(new_n275_), .B2(new_n282_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n263_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n248_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n260_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n251_), .A2(new_n253_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT8), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n254_), .A2(new_n249_), .A3(new_n260_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n286_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n273_), .A2(new_n274_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G232gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT34), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT35), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n295_), .A2(KEYINPUT35), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n285_), .A2(new_n293_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n285_), .A2(KEYINPUT72), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT15), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT71), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n280_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n275_), .A2(new_n282_), .A3(KEYINPUT15), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(new_n263_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n309_), .A3(new_n293_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n300_), .B1(new_n310_), .B2(new_n297_), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n312_));
  XNOR2_X1  g111(.A(G190gat), .B(G218gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT73), .ZN(new_n314_));
  INV_X1    g113(.A(G134gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G162gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n311_), .A2(new_n312_), .A3(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(KEYINPUT36), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n291_), .B1(new_n306_), .B2(new_n305_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n321_), .A2(new_n308_), .B1(new_n292_), .B2(new_n291_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n296_), .B1(new_n322_), .B2(new_n301_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n320_), .B1(new_n323_), .B2(new_n300_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT37), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n319_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n319_), .A2(new_n324_), .A3(KEYINPUT77), .A4(new_n325_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT36), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n318_), .B(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n311_), .B2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n320_), .B(KEYINPUT75), .C1(new_n323_), .C2(new_n300_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n319_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n336_), .A2(KEYINPUT76), .A3(KEYINPUT37), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT76), .B1(new_n336_), .B2(KEYINPUT37), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n330_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(KEYINPUT78), .B(new_n330_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n232_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(G127gat), .A2(G134gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G127gat), .A2(G134gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(G113gat), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G127gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n315_), .ZN(new_n351_));
  INV_X1    g150(.A(G113gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G127gat), .A2(G134gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n349_), .A2(new_n354_), .A3(G120gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(G120gat), .B1(new_n349_), .B2(new_n354_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT89), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G120gat), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n347_), .A2(new_n348_), .A3(G113gat), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n352_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n359_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n349_), .A2(new_n354_), .A3(G120gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT89), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT93), .B(KEYINPUT2), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT94), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G141gat), .ZN(new_n370_));
  INV_X1    g169(.A(G148gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(KEYINPUT3), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n372_), .A2(new_n374_), .B1(new_n368_), .B2(KEYINPUT2), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT94), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT2), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n377_), .A2(KEYINPUT93), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(KEYINPUT93), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n376_), .B(new_n367_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n369_), .A2(new_n375_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n382_));
  INV_X1    g181(.A(G155gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n317_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT91), .B1(G155gat), .B2(G162gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT92), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(KEYINPUT1), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(G155gat), .A3(G162gat), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n386_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G141gat), .B(G148gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n390_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  AOI211_X1 g197(.A(KEYINPUT92), .B(new_n396_), .C1(new_n394_), .C2(new_n386_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n389_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT4), .B1(new_n365_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT98), .ZN(new_n403_));
  INV_X1    g202(.A(new_n385_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(KEYINPUT91), .A2(G155gat), .A3(G162gat), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n391_), .A2(new_n393_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n397_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT92), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n395_), .A2(new_n390_), .A3(new_n397_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n355_), .A2(new_n356_), .ZN(new_n412_));
  AND4_X1   g211(.A1(new_n403_), .A2(new_n411_), .A3(new_n389_), .A4(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n389_), .A3(new_n412_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n409_), .A2(new_n410_), .B1(new_n388_), .B2(new_n381_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n357_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n362_), .A2(KEYINPUT89), .A3(new_n363_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n403_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n413_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n346_), .B(new_n402_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n414_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n415_), .A2(new_n403_), .A3(new_n412_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n346_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G85gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT0), .ZN(new_n430_));
  INV_X1    g229(.A(G57gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n432_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT104), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT18), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(G64gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(G92gat), .ZN(new_n441_));
  INV_X1    g240(.A(G64gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n439_), .B(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n244_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G226gat), .A2(G233gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n447_), .B(KEYINPUT97), .Z(new_n448_));
  XOR2_X1   g247(.A(new_n448_), .B(KEYINPUT19), .Z(new_n449_));
  AND2_X1   g248(.A1(KEYINPUT95), .A2(G197gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(KEYINPUT95), .A2(G197gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(G204gat), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT96), .B(G204gat), .ZN(new_n453_));
  INV_X1    g252(.A(G197gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G211gat), .B(G218gat), .Z(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(KEYINPUT21), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT21), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n452_), .B(new_n458_), .C1(new_n454_), .C2(new_n453_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n456_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n450_), .A2(new_n451_), .ZN(new_n462_));
  INV_X1    g261(.A(G204gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n453_), .A2(new_n454_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n458_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n457_), .B1(new_n461_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT22), .B(G169gat), .ZN(new_n468_));
  INV_X1    g267(.A(G176gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G169gat), .A2(G176gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G183gat), .A2(G190gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(KEYINPUT23), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(new_n474_), .B2(new_n472_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G183gat), .A2(G190gat), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n470_), .B(new_n471_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n472_), .A2(KEYINPUT23), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n474_), .B2(new_n472_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n471_), .A2(KEYINPUT24), .ZN(new_n481_));
  INV_X1    g280(.A(G169gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n469_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n480_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT25), .B(G183gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT26), .B(G190gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n479_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n477_), .A2(new_n488_), .ZN(new_n489_));
  OAI211_X1 g288(.A(KEYINPUT100), .B(KEYINPUT20), .C1(new_n467_), .C2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n476_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n479_), .A2(new_n491_), .B1(G169gat), .B2(G176gat), .ZN(new_n492_));
  AND2_X1   g291(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n493_));
  NOR2_X1   g292(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n494_));
  OAI21_X1  g293(.A(G169gat), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n482_), .A2(KEYINPUT22), .ZN(new_n498_));
  OAI211_X1 g297(.A(KEYINPUT86), .B(G169gat), .C1(new_n493_), .C2(new_n494_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n497_), .A2(new_n469_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n492_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT25), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT83), .B1(new_n502_), .B2(G183gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT83), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n504_), .B(new_n486_), .C1(new_n485_), .C2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n474_), .A2(new_n472_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n506_), .B(new_n484_), .C1(new_n507_), .C2(new_n473_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n467_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n490_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n463_), .A2(KEYINPUT96), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT96), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(G204gat), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n512_), .A2(new_n514_), .A3(new_n454_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n450_), .A2(new_n451_), .A3(G204gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT21), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n518_), .A2(new_n457_), .A3(new_n477_), .A4(new_n488_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT100), .B1(new_n519_), .B2(KEYINPUT20), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n449_), .B1(new_n511_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n522_));
  INV_X1    g321(.A(new_n467_), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT25), .B(G183gat), .Z(new_n524_));
  AOI21_X1  g323(.A(new_n503_), .B1(new_n524_), .B2(KEYINPUT83), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n475_), .B1(new_n525_), .B2(new_n486_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n526_), .A2(new_n484_), .B1(new_n492_), .B2(new_n500_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n522_), .B1(new_n523_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n449_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n467_), .A2(new_n489_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n446_), .B1(new_n521_), .B2(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n530_), .B(KEYINPUT20), .C1(new_n467_), .C2(new_n509_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n449_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n510_), .A2(KEYINPUT20), .A3(new_n529_), .A4(new_n519_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n534_), .A2(new_n446_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT27), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n532_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n539_));
  INV_X1    g338(.A(new_n535_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n529_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n445_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n534_), .A2(new_n446_), .A3(new_n535_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n539_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n437_), .B1(new_n538_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n521_), .A2(new_n531_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n445_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(KEYINPUT27), .A3(new_n543_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n539_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n446_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(new_n536_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(KEYINPUT104), .A3(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n436_), .A2(new_n545_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n365_), .B(KEYINPUT31), .ZN(new_n554_));
  XOR2_X1   g353(.A(G71gat), .B(G99gat), .Z(new_n555_));
  NAND2_X1  g354(.A1(G227gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G15gat), .B(G43gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n501_), .A2(new_n561_), .A3(new_n508_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n501_), .B2(new_n508_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n509_), .A2(KEYINPUT30), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n501_), .A2(new_n561_), .A3(new_n508_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n560_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT90), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n564_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n567_), .A2(new_n568_), .A3(new_n566_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n559_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n570_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n554_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n570_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n554_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n400_), .A2(KEYINPUT29), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n467_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(G50gat), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n276_), .A3(new_n467_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G78gat), .B(G106gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n589_), .A3(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G228gat), .A2(G233gat), .ZN(new_n592_));
  INV_X1    g391(.A(G22gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n400_), .A2(KEYINPUT29), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT28), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n595_), .A2(new_n596_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n594_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n594_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n591_), .A2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n588_), .A2(new_n603_), .A3(new_n600_), .A4(new_n590_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n581_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT105), .B1(new_n553_), .B2(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n538_), .A2(new_n437_), .A3(new_n544_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT104), .B1(new_n548_), .B2(new_n551_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT105), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n577_), .A2(new_n580_), .B1(new_n606_), .B2(new_n605_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n436_), .A4(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n617_));
  OAI21_X1  g416(.A(KEYINPUT33), .B1(new_n435_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT98), .B1(new_n365_), .B2(new_n400_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n414_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n424_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n401_), .B1(new_n622_), .B2(KEYINPUT4), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n425_), .B1(new_n623_), .B2(new_n346_), .ZN(new_n624_));
  OAI211_X1 g423(.A(KEYINPUT99), .B(new_n619_), .C1(new_n624_), .C2(new_n434_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n542_), .A2(new_n543_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n402_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n432_), .B1(new_n627_), .B2(new_n345_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n420_), .A2(new_n346_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n626_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n618_), .A2(new_n625_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n441_), .A2(new_n444_), .A3(KEYINPUT32), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n546_), .B2(new_n634_), .ZN(new_n635_));
  AOI211_X1 g434(.A(KEYINPUT101), .B(new_n633_), .C1(new_n521_), .C2(new_n531_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n534_), .A2(new_n535_), .A3(new_n633_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n637_), .B(new_n638_), .C1(new_n433_), .C2(new_n435_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n631_), .A2(new_n639_), .A3(new_n607_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n624_), .A2(new_n434_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n427_), .A2(new_n432_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n548_), .A4(new_n551_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n605_), .A2(new_n606_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n581_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n640_), .A2(KEYINPUT103), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT103), .B1(new_n640_), .B2(new_n645_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n616_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT70), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT5), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(G176gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(G204gat), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT68), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n291_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT66), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT66), .B1(new_n291_), .B2(new_n656_), .ZN(new_n660_));
  OAI22_X1  g459(.A1(new_n659_), .A2(new_n660_), .B1(new_n291_), .B2(new_n656_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT12), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n665_), .B1(new_n291_), .B2(new_n656_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n263_), .A2(KEYINPUT12), .A3(new_n208_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT67), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n263_), .A2(new_n208_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(new_n663_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n657_), .A2(KEYINPUT67), .A3(new_n662_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n668_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n655_), .B1(new_n664_), .B2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n671_), .A2(new_n672_), .ZN(new_n675_));
  AOI22_X1  g474(.A1(new_n675_), .A2(new_n668_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT69), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n653_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n664_), .A2(new_n673_), .A3(new_n653_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT69), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n674_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT13), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT13), .B(new_n674_), .C1(new_n678_), .C2(new_n680_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n649_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n674_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n677_), .B1(new_n676_), .B2(new_n653_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n679_), .A2(KEYINPUT69), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT13), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n681_), .A2(new_n682_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(KEYINPUT70), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n307_), .A2(new_n215_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(G229gat), .A2(G233gat), .ZN(new_n694_));
  INV_X1    g493(.A(new_n215_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n292_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n215_), .B(new_n292_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(KEYINPUT81), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(KEYINPUT81), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n701_), .B2(new_n694_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(G113gat), .B(G141gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(new_n482_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(new_n454_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT82), .ZN(new_n707_));
  INV_X1    g506(.A(new_n705_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n697_), .B(new_n708_), .C1(new_n701_), .C2(new_n694_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n706_), .A2(new_n707_), .A3(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n702_), .A2(KEYINPUT82), .A3(new_n705_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n685_), .A2(new_n692_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n648_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n344_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n436_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n210_), .A3(new_n717_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT38), .Z(new_n719_));
  NAND2_X1  g518(.A1(new_n319_), .A2(new_n324_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n232_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n715_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n210_), .B1(new_n724_), .B2(new_n717_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n719_), .A2(new_n725_), .ZN(G1324gat));
  INV_X1    g525(.A(new_n612_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n211_), .B1(new_n724_), .B2(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT39), .Z(new_n729_));
  NAND3_X1  g528(.A1(new_n716_), .A2(new_n211_), .A3(new_n727_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g531(.A(G15gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n724_), .B2(new_n581_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT41), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n716_), .A2(new_n733_), .A3(new_n581_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1326gat));
  AOI21_X1  g536(.A(new_n593_), .B1(new_n724_), .B2(new_n644_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT42), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n716_), .A2(new_n593_), .A3(new_n644_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1327gat));
  NOR2_X1   g540(.A1(new_n231_), .A2(new_n720_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n648_), .A2(new_n714_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT108), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n648_), .A2(new_n714_), .A3(new_n745_), .A4(new_n742_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n267_), .A3(new_n717_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n714_), .A2(new_n232_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n640_), .A2(new_n645_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT103), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n640_), .A2(KEYINPUT103), .A3(new_n645_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n754_), .A2(new_n755_), .B1(new_n609_), .B2(new_n615_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n341_), .A2(new_n342_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(KEYINPUT43), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n336_), .A2(KEYINPUT37), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT76), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n336_), .A2(KEYINPUT76), .A3(KEYINPUT37), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT78), .B1(new_n764_), .B2(new_n330_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n342_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n759_), .B1(new_n767_), .B2(new_n648_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n751_), .B1(new_n758_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n749_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT43), .B1(new_n756_), .B2(new_n757_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n767_), .A2(new_n759_), .A3(new_n648_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n750_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n771_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n769_), .A2(new_n777_), .A3(new_n770_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT106), .B1(new_n774_), .B2(KEYINPUT44), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n776_), .A2(new_n717_), .A3(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n748_), .B1(new_n781_), .B2(new_n267_), .ZN(G1328gat));
  NAND4_X1  g581(.A1(new_n780_), .A2(new_n727_), .A3(new_n771_), .A4(new_n775_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(G36gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n612_), .B(KEYINPUT109), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n744_), .A2(new_n268_), .A3(new_n746_), .A4(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(KEYINPUT110), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(KEYINPUT110), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n747_), .A2(new_n791_), .A3(new_n268_), .A4(new_n785_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n786_), .A2(KEYINPUT110), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n790_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n784_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n799_));
  AOI211_X1 g598(.A(KEYINPUT111), .B(new_n799_), .C1(new_n784_), .C2(new_n795_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1329gat));
  NAND4_X1  g600(.A1(new_n776_), .A2(G43gat), .A3(new_n581_), .A4(new_n780_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n747_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n581_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n270_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g606(.A1(new_n747_), .A2(new_n276_), .A3(new_n644_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n776_), .A2(new_n644_), .A3(new_n780_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n276_), .ZN(G1331gat));
  AND2_X1   g609(.A1(new_n685_), .A2(new_n692_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(new_n648_), .A3(new_n712_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n723_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n815_), .A2(new_n431_), .A3(new_n436_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n813_), .A2(new_n344_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n817_), .A2(KEYINPUT112), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(KEYINPUT112), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n717_), .A3(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(new_n431_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n821_), .A2(KEYINPUT113), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(KEYINPUT113), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n816_), .B1(new_n822_), .B2(new_n823_), .ZN(G1332gat));
  NAND3_X1  g623(.A1(new_n817_), .A2(new_n442_), .A3(new_n785_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n785_), .ZN(new_n826_));
  OAI21_X1  g625(.A(G64gat), .B1(new_n815_), .B2(new_n826_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n827_), .A2(KEYINPUT114), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(KEYINPUT114), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n828_), .A2(KEYINPUT48), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT48), .B1(new_n828_), .B2(new_n829_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n825_), .B1(new_n830_), .B2(new_n831_), .ZN(G1333gat));
  INV_X1    g631(.A(G71gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n814_), .B2(new_n581_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT49), .Z(new_n835_));
  NAND3_X1  g634(.A1(new_n817_), .A2(new_n833_), .A3(new_n581_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1334gat));
  INV_X1    g636(.A(G78gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n814_), .B2(new_n644_), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT50), .Z(new_n840_));
  NAND3_X1  g639(.A1(new_n817_), .A2(new_n838_), .A3(new_n644_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1335gat));
  NOR3_X1   g641(.A1(new_n813_), .A2(new_n720_), .A3(new_n231_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G85gat), .B1(new_n843_), .B2(new_n717_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n772_), .A2(new_n773_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n845_), .A2(KEYINPUT115), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n811_), .A2(new_n713_), .A3(new_n231_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(KEYINPUT115), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n436_), .A2(new_n243_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n844_), .B1(new_n850_), .B2(new_n851_), .ZN(G1336gat));
  AOI21_X1  g651(.A(G92gat), .B1(new_n843_), .B2(new_n727_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n826_), .A2(new_n244_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n850_), .B2(new_n854_), .ZN(G1337gat));
  OAI21_X1  g654(.A(G99gat), .B1(new_n849_), .B2(new_n804_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n804_), .A2(new_n233_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n843_), .A2(new_n857_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n859_));
  NAND3_X1  g658(.A1(new_n856_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n860_), .A2(KEYINPUT117), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT51), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(KEYINPUT117), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n863_), .A3(new_n864_), .ZN(G1338gat));
  NAND3_X1  g664(.A1(new_n845_), .A2(new_n644_), .A3(new_n847_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G106gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT52), .ZN(new_n868_));
  INV_X1    g667(.A(G106gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n843_), .A2(new_n869_), .A3(new_n644_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n673_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n659_), .A2(new_n660_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n666_), .A2(new_n667_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n663_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n668_), .A2(new_n671_), .A3(KEYINPUT55), .A4(new_n672_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n874_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n655_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n874_), .A2(new_n877_), .A3(KEYINPUT118), .A4(new_n878_), .ZN(new_n883_));
  AND4_X1   g682(.A1(KEYINPUT56), .A2(new_n881_), .A3(new_n882_), .A4(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n712_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT56), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n881_), .A2(KEYINPUT56), .A3(new_n882_), .A4(new_n883_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(KEYINPUT119), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n678_), .A2(new_n680_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n886_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n701_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n694_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n693_), .A2(new_n696_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n897_), .B(new_n705_), .C1(new_n694_), .C2(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n689_), .A2(new_n709_), .A3(new_n899_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n886_), .A2(new_n891_), .A3(KEYINPUT120), .A4(new_n892_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n895_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n720_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n889_), .A2(new_n890_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n906_), .A2(new_n709_), .A3(new_n892_), .A4(new_n899_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT58), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n767_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n902_), .A2(KEYINPUT57), .A3(new_n720_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n905_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n343_), .B(new_n712_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT54), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n912_), .A2(KEYINPUT54), .ZN(new_n914_));
  AOI22_X1  g713(.A1(new_n911_), .A2(new_n232_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n727_), .A2(new_n436_), .A3(new_n608_), .ZN(new_n916_));
  XOR2_X1   g715(.A(new_n916_), .B(KEYINPUT121), .Z(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n915_), .A2(new_n712_), .A3(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT122), .B1(new_n919_), .B2(G113gat), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n911_), .A2(new_n232_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n914_), .A2(new_n913_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n917_), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n921_), .B(new_n352_), .C1(new_n925_), .C2(new_n712_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n920_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928_));
  AOI21_X1  g727(.A(KEYINPUT59), .B1(new_n924_), .B2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n925_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n924_), .B(new_n917_), .C1(new_n928_), .C2(KEYINPUT59), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n712_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n927_), .B1(new_n932_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g732(.A(new_n925_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n811_), .B2(G120gat), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n934_), .B(new_n936_), .C1(new_n935_), .C2(G120gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n811_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n359_), .ZN(G1341gat));
  AOI21_X1  g738(.A(G127gat), .B1(new_n934_), .B2(new_n231_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n232_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g741(.A(G134gat), .B1(new_n934_), .B2(new_n721_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n757_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n944_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g744(.A1(new_n581_), .A2(new_n607_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n924_), .A2(new_n717_), .A3(new_n826_), .A4(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n712_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n370_), .ZN(G1344gat));
  NOR2_X1   g748(.A1(new_n947_), .A2(new_n811_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(new_n371_), .ZN(G1345gat));
  NOR2_X1   g750(.A1(new_n947_), .A2(new_n232_), .ZN(new_n952_));
  XOR2_X1   g751(.A(KEYINPUT61), .B(G155gat), .Z(new_n953_));
  XNOR2_X1  g752(.A(new_n952_), .B(new_n953_), .ZN(G1346gat));
  INV_X1    g753(.A(new_n947_), .ZN(new_n955_));
  AOI21_X1  g754(.A(G162gat), .B1(new_n955_), .B2(new_n721_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n767_), .A2(G162gat), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(KEYINPUT124), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n956_), .B1(new_n955_), .B2(new_n958_), .ZN(G1347gat));
  NOR2_X1   g758(.A1(new_n826_), .A2(new_n717_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n924_), .A2(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(new_n608_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n962_), .A2(new_n713_), .A3(new_n468_), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n924_), .A2(new_n713_), .A3(new_n614_), .A4(new_n960_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(G169gat), .ZN(new_n965_));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n964_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n963_), .A2(new_n967_), .A3(new_n968_), .ZN(G1348gat));
  NOR3_X1   g768(.A1(new_n915_), .A2(new_n717_), .A3(new_n826_), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n970_), .A2(new_n812_), .A3(new_n614_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n972_));
  AND2_X1   g771(.A1(new_n971_), .A2(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n972_), .B1(new_n971_), .B2(new_n974_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n973_), .A2(new_n975_), .ZN(G1349gat));
  NAND2_X1  g775(.A1(new_n970_), .A2(new_n614_), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n977_), .A2(new_n485_), .A3(new_n232_), .ZN(new_n978_));
  AOI21_X1  g777(.A(G183gat), .B1(new_n962_), .B2(new_n231_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n978_), .A2(new_n979_), .ZN(G1350gat));
  OAI21_X1  g779(.A(G190gat), .B1(new_n977_), .B2(new_n757_), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n962_), .A2(new_n486_), .A3(new_n721_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n981_), .A2(new_n982_), .ZN(G1351gat));
  AND3_X1   g782(.A1(new_n924_), .A2(new_n946_), .A3(new_n960_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n984_), .A2(new_n713_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n985_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g785(.A1(new_n924_), .A2(new_n812_), .A3(new_n946_), .A4(new_n960_), .ZN(new_n987_));
  OR3_X1    g786(.A1(new_n987_), .A2(KEYINPUT126), .A3(new_n453_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n987_), .A2(G204gat), .ZN(new_n989_));
  OAI21_X1  g788(.A(KEYINPUT126), .B1(new_n987_), .B2(new_n453_), .ZN(new_n990_));
  NAND3_X1  g789(.A1(new_n988_), .A2(new_n989_), .A3(new_n990_), .ZN(G1353gat));
  NAND4_X1  g790(.A1(new_n924_), .A2(new_n231_), .A3(new_n946_), .A4(new_n960_), .ZN(new_n992_));
  XNOR2_X1  g791(.A(KEYINPUT63), .B(G211gat), .ZN(new_n993_));
  NOR2_X1   g792(.A1(new_n992_), .A2(new_n993_), .ZN(new_n994_));
  INV_X1    g793(.A(KEYINPUT63), .ZN(new_n995_));
  NAND3_X1  g794(.A1(new_n992_), .A2(new_n995_), .A3(new_n222_), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n996_), .A2(KEYINPUT127), .ZN(new_n997_));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998_));
  NAND4_X1  g797(.A1(new_n992_), .A2(new_n998_), .A3(new_n995_), .A4(new_n222_), .ZN(new_n999_));
  AOI21_X1  g798(.A(new_n994_), .B1(new_n997_), .B2(new_n999_), .ZN(G1354gat));
  AOI21_X1  g799(.A(G218gat), .B1(new_n984_), .B2(new_n721_), .ZN(new_n1001_));
  AND2_X1   g800(.A1(new_n767_), .A2(G218gat), .ZN(new_n1002_));
  AOI21_X1  g801(.A(new_n1001_), .B1(new_n984_), .B2(new_n1002_), .ZN(G1355gat));
endmodule


