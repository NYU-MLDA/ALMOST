//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT8), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n205_), .B(new_n206_), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT7), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n208_), .B(new_n209_), .C1(G99gat), .C2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT6), .B1(new_n205_), .B2(new_n206_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  AOI21_X1  g016(.A(new_n204_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n215_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n212_), .A2(KEYINPUT66), .A3(new_n214_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n211_), .A3(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n217_), .A2(new_n204_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n218_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT10), .B(G99gat), .Z(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n206_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(G85gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT9), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(G92gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n220_), .A2(new_n221_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n203_), .B1(new_n224_), .B2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n231_), .A2(new_n232_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n222_), .A2(new_n223_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n235_), .B(KEYINPUT70), .C1(new_n236_), .C2(new_n218_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G78gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(KEYINPUT11), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n241_));
  INV_X1    g040(.A(new_n239_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n240_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT12), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n244_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT71), .B1(new_n249_), .B2(new_n240_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n234_), .A2(new_n237_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n224_), .A2(new_n233_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n253_), .B1(new_n254_), .B2(new_n245_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G230gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT64), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n254_), .B2(new_n245_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n252_), .A2(new_n255_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n254_), .A2(new_n261_), .A3(new_n245_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n235_), .B(new_n245_), .C1(new_n236_), .C2(new_n218_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT68), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n254_), .A2(new_n245_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n262_), .A2(new_n264_), .A3(KEYINPUT69), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n260_), .B1(new_n270_), .B2(new_n257_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G120gat), .B(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT5), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G176gat), .B(G204gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n271_), .A2(new_n276_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n202_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G15gat), .B(G22gat), .ZN(new_n281_));
  INV_X1    g080(.A(G1gat), .ZN(new_n282_));
  INV_X1    g081(.A(G8gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT14), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G1gat), .B(G8gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G29gat), .B(G36gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G43gat), .B(G50gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n287_), .B(new_n290_), .Z(new_n291_));
  NAND2_X1  g090(.A1(G229gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n290_), .B(KEYINPUT15), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n287_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n287_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n290_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n298_), .A3(new_n292_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G113gat), .B(G141gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G169gat), .B(G197gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT77), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n294_), .A2(new_n299_), .A3(KEYINPUT77), .A4(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n294_), .A2(new_n299_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n302_), .B(KEYINPUT76), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n305_), .A2(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n270_), .A2(new_n257_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n259_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n275_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(KEYINPUT13), .A3(new_n277_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G231gat), .A2(G233gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n245_), .B(new_n315_), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n287_), .B(KEYINPUT75), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G127gat), .B(G155gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT16), .ZN(new_n321_));
  XOR2_X1   g120(.A(G183gat), .B(G211gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(new_n246_), .A3(KEYINPUT17), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n319_), .A2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(KEYINPUT17), .B2(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n318_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n280_), .A2(new_n310_), .A3(new_n314_), .A4(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT101), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G1gat), .B(G29gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G85gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT0), .B(G57gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n336_), .B(KEYINPUT96), .Z(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G127gat), .B(G134gat), .Z(new_n339_));
  XOR2_X1   g138(.A(G113gat), .B(G120gat), .Z(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G127gat), .B(G134gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G113gat), .B(G120gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n346_));
  INV_X1    g145(.A(G141gat), .ZN(new_n347_));
  INV_X1    g146(.A(G148gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT3), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n350_), .B1(G141gat), .B2(G148gat), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n346_), .B1(new_n352_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT83), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT83), .A3(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n349_), .A2(new_n351_), .ZN(new_n366_));
  AND3_X1   g165(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n367_), .A2(new_n353_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n368_), .A3(KEYINPUT82), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n357_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n347_), .A2(new_n348_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT1), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n363_), .B1(new_n360_), .B2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n359_), .A2(KEYINPUT1), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n371_), .B(new_n372_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  AOI211_X1 g175(.A(KEYINPUT4), .B(new_n345_), .C1(new_n370_), .C2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT95), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n341_), .A2(new_n378_), .A3(new_n344_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n369_), .A2(new_n365_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT82), .B1(new_n366_), .B2(new_n368_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n379_), .B(new_n376_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n345_), .A2(KEYINPUT95), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n370_), .A2(new_n383_), .A3(new_n379_), .A4(new_n376_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  AOI211_X1 g186(.A(new_n338_), .B(new_n377_), .C1(new_n387_), .C2(KEYINPUT4), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n337_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n335_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n339_), .B(new_n343_), .ZN(new_n391_));
  AOI211_X1 g190(.A(new_n378_), .B(new_n391_), .C1(new_n370_), .C2(new_n376_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n382_), .A2(new_n384_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT4), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n377_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n337_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n389_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n335_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n390_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT29), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n370_), .A2(new_n401_), .A3(new_n376_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT28), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G22gat), .B(G50gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n376_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT29), .ZN(new_n407_));
  INV_X1    g206(.A(G218gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G211gat), .ZN(new_n409_));
  INV_X1    g208(.A(G211gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G218gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n413_));
  INV_X1    g212(.A(G204gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G197gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT21), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(G197gat), .B2(G204gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n412_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n415_), .A2(G197gat), .A3(new_n417_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n416_), .A2(KEYINPUT88), .A3(G204gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT88), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n414_), .B2(G197gat), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n422_), .A2(new_n419_), .A3(new_n423_), .A4(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT89), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n419_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n429_));
  AND2_X1   g228(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n416_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(new_n423_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n428_), .B(new_n429_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n422_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n428_), .B1(new_n436_), .B2(new_n429_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n427_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n407_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(G233gat), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n440_), .A2(KEYINPUT86), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(KEYINPUT86), .ZN(new_n442_));
  OAI21_X1  g241(.A(G228gat), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G78gat), .B(G106gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT85), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n407_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n406_), .A2(KEYINPUT85), .A3(KEYINPUT29), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n429_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT89), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n453_), .A2(new_n434_), .B1(new_n426_), .B2(new_n421_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(new_n444_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n447_), .B1(new_n451_), .B2(new_n455_), .ZN(new_n456_));
  AOI211_X1 g255(.A(new_n448_), .B(new_n401_), .C1(new_n370_), .C2(new_n376_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT85), .B1(new_n406_), .B2(KEYINPUT29), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n447_), .B(new_n455_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n445_), .B(new_n446_), .C1(new_n456_), .C2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT84), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n455_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT90), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n464_), .A2(new_n459_), .B1(new_n444_), .B2(new_n439_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(new_n446_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n405_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n465_), .B2(new_n446_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n405_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n445_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n446_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n469_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n467_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT27), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G226gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT19), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT91), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G183gat), .A2(G190gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT23), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n483_));
  INV_X1    g282(.A(G169gat), .ZN(new_n484_));
  INV_X1    g283(.A(G176gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n482_), .B(new_n483_), .C1(new_n486_), .C2(KEYINPUT24), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n484_), .A2(new_n485_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT25), .B(G183gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT26), .B(G190gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT78), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n493_), .A3(KEYINPUT78), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n491_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G169gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n484_), .A2(KEYINPUT79), .A3(KEYINPUT22), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n485_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT80), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT80), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n500_), .A2(new_n501_), .A3(new_n504_), .A4(new_n485_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n488_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n482_), .B(new_n483_), .C1(G183gat), .C2(G190gat), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n503_), .A2(new_n505_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n498_), .A2(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n479_), .B(KEYINPUT20), .C1(new_n438_), .C2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT26), .B(G190gat), .Z(new_n511_));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n493_), .A2(KEYINPUT92), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n492_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n491_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT22), .B(G169gat), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n488_), .B1(new_n517_), .B2(new_n485_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n507_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n438_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n510_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n453_), .A2(new_n434_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n523_), .A2(new_n427_), .A3(new_n508_), .A4(new_n498_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n479_), .B1(new_n524_), .B2(KEYINPUT20), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n478_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G8gat), .B(G36gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G64gat), .B(G92gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n438_), .A2(new_n520_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT93), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n535_));
  AOI211_X1 g334(.A(new_n535_), .B(new_n478_), .C1(new_n438_), .C2(new_n509_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n438_), .B2(new_n520_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n534_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n526_), .A2(new_n532_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n532_), .B1(new_n526_), .B2(new_n539_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n476_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n478_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n515_), .A2(new_n491_), .B1(new_n507_), .B2(new_n518_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n535_), .B1(new_n454_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT98), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n545_), .A2(new_n546_), .B1(new_n438_), .B2(new_n509_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT98), .B1(new_n533_), .B2(new_n535_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n543_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n522_), .A2(new_n525_), .A3(new_n478_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n531_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n526_), .A2(new_n532_), .A3(new_n539_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(KEYINPUT27), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n542_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G227gat), .A2(G233gat), .ZN(new_n555_));
  INV_X1    g354(.A(G15gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT30), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n509_), .B(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n391_), .A2(KEYINPUT31), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT81), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n391_), .A2(KEYINPUT31), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n559_), .A2(new_n564_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G71gat), .B(G99gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G43gat), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OR3_X1    g368(.A1(new_n565_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n377_), .B1(new_n387_), .B2(KEYINPUT4), .ZN(new_n573_));
  AOI211_X1 g372(.A(new_n389_), .B(new_n335_), .C1(new_n573_), .C2(new_n337_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n398_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n475_), .A2(new_n554_), .A3(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n462_), .A2(new_n466_), .A3(new_n405_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n470_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n540_), .A2(new_n541_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT33), .B1(new_n574_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n399_), .A2(KEYINPUT97), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n573_), .A2(new_n338_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n398_), .B1(new_n387_), .B2(new_n337_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n582_), .A2(new_n584_), .A3(new_n586_), .A4(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n532_), .A2(KEYINPUT32), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n526_), .A2(new_n539_), .A3(new_n591_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT99), .B1(new_n595_), .B2(new_n576_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n400_), .A2(new_n597_), .A3(new_n593_), .A4(new_n594_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n581_), .A2(new_n590_), .A3(new_n596_), .A4(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n542_), .A2(new_n553_), .A3(new_n576_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n572_), .B1(new_n475_), .B2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n578_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT34), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT35), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT72), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n234_), .A2(new_n237_), .A3(new_n295_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT73), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n604_), .A2(KEYINPUT35), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n254_), .B2(new_n290_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n607_), .B(new_n611_), .C1(new_n608_), .C2(new_n606_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT36), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT74), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n618_), .A2(KEYINPUT36), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n613_), .A2(new_n614_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT74), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n615_), .A2(new_n624_), .A3(new_n619_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n621_), .A2(KEYINPUT102), .A3(new_n623_), .A4(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n602_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n331_), .A2(new_n400_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G1gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT103), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT37), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n626_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n620_), .A2(KEYINPUT37), .A3(new_n623_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n329_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n314_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT13), .B1(new_n313_), .B2(new_n277_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT100), .B1(new_n602_), .B2(new_n309_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n572_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n600_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n596_), .A2(new_n474_), .A3(new_n467_), .A4(new_n598_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n590_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n646_), .B(new_n647_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n475_), .A2(new_n554_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n577_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n310_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n644_), .B1(new_n645_), .B2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n282_), .A3(new_n400_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(KEYINPUT38), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n658_), .A2(KEYINPUT38), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n634_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n634_), .B(KEYINPUT104), .C1(new_n659_), .C2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1324gat));
  NAND3_X1  g464(.A1(new_n657_), .A2(new_n283_), .A3(new_n554_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n331_), .A2(new_n554_), .A3(new_n631_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  AND4_X1   g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .A4(G8gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n283_), .B1(KEYINPUT105), .B2(KEYINPUT39), .ZN(new_n671_));
  AOI22_X1  g470(.A1(new_n668_), .A2(new_n671_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n666_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1325gat));
  AND2_X1   g474(.A1(new_n331_), .A2(new_n631_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n556_), .B1(new_n676_), .B2(new_n572_), .ZN(new_n677_));
  XOR2_X1   g476(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n657_), .A2(new_n556_), .A3(new_n572_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n678_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(G1326gat));
  INV_X1    g481(.A(G22gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n657_), .A2(new_n683_), .A3(new_n475_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n676_), .A2(new_n475_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(G22gat), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT42), .B(new_n683_), .C1(new_n676_), .C2(new_n475_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(new_n630_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n329_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n643_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n656_), .B2(new_n645_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n400_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n637_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n626_), .B2(new_n635_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n602_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n654_), .A2(new_n698_), .A3(new_n638_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n643_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n701_), .A2(new_n309_), .A3(new_n329_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n700_), .A2(KEYINPUT44), .A3(new_n702_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n400_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n694_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n706_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n554_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G36gat), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(G36gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n693_), .B2(new_n714_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n693_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n712_), .B(KEYINPUT46), .C1(new_n715_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  XNOR2_X1  g520(.A(KEYINPUT108), .B(G43gat), .ZN(new_n722_));
  INV_X1    g521(.A(new_n693_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n646_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n572_), .A2(G43gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n710_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g526(.A1(new_n723_), .A2(G50gat), .A3(new_n581_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n707_), .A2(new_n475_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n729_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT109), .B1(new_n729_), .B2(G50gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(new_n730_), .B2(new_n731_), .ZN(G1331gat));
  NOR3_X1   g531(.A1(new_n643_), .A2(new_n310_), .A3(new_n639_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n631_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(G57gat), .A3(new_n400_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n602_), .A2(new_n310_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n737_), .A2(new_n701_), .A3(new_n640_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n400_), .ZN(new_n739_));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(KEYINPUT110), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(KEYINPUT110), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n736_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT111), .B(new_n736_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1332gat));
  OAI21_X1  g547(.A(G64gat), .B1(new_n734_), .B2(new_n711_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT48), .ZN(new_n750_));
  INV_X1    g549(.A(G64gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n738_), .A2(new_n751_), .A3(new_n554_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1333gat));
  OAI21_X1  g552(.A(G71gat), .B1(new_n734_), .B2(new_n646_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT49), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n646_), .A2(G71gat), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT112), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n738_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(G1334gat));
  INV_X1    g558(.A(G78gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n738_), .A2(new_n760_), .A3(new_n475_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G78gat), .B1(new_n734_), .B2(new_n581_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(KEYINPUT50), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(KEYINPUT50), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT113), .ZN(G1335gat));
  NAND3_X1  g565(.A1(new_n737_), .A2(new_n701_), .A3(new_n691_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n400_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n309_), .B(new_n639_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT114), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n400_), .A2(new_n228_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1336gat));
  INV_X1    g573(.A(G92gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n768_), .A2(new_n775_), .A3(new_n554_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n772_), .A2(new_n554_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n775_), .ZN(G1337gat));
  AOI21_X1  g577(.A(new_n205_), .B1(new_n772_), .B2(new_n572_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n768_), .A2(new_n572_), .A3(new_n226_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OR3_X1    g580(.A1(new_n779_), .A2(KEYINPUT51), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT51), .B1(new_n779_), .B2(new_n781_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1338gat));
  NAND3_X1  g583(.A1(new_n768_), .A2(new_n206_), .A3(new_n475_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n581_), .B(new_n770_), .C1(new_n697_), .C2(new_n699_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n206_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n771_), .B2(new_n475_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n786_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n770_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n698_), .B1(new_n654_), .B2(new_n638_), .ZN(new_n794_));
  AOI211_X1 g593(.A(KEYINPUT43), .B(new_n696_), .C1(new_n650_), .C2(new_n653_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n475_), .B(new_n793_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G106gat), .B1(new_n796_), .B2(KEYINPUT115), .ZN(new_n797_));
  INV_X1    g596(.A(new_n786_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n797_), .A2(new_n790_), .A3(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n785_), .B1(new_n792_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n785_), .C1(new_n792_), .C2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1339gat));
  NAND3_X1  g603(.A1(new_n640_), .A2(new_n309_), .A3(new_n643_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n805_), .B(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT121), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n252_), .A2(new_n255_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n810_), .A2(new_n811_), .A3(KEYINPUT55), .A4(new_n258_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT119), .B1(new_n259_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n252_), .A2(new_n255_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n257_), .B1(new_n815_), .B2(new_n265_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n259_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n812_), .A2(new_n814_), .A3(new_n816_), .A4(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n275_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n305_), .A2(new_n306_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n302_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n296_), .A2(new_n298_), .A3(new_n293_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n278_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n824_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n824_), .A2(new_n830_), .A3(KEYINPUT58), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n638_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n819_), .B2(new_n275_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n837_), .A2(new_n838_), .A3(KEYINPUT120), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n819_), .A2(KEYINPUT120), .A3(KEYINPUT56), .A4(new_n275_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n309_), .B1(new_n271_), .B2(new_n276_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n313_), .A2(new_n277_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OAI22_X1  g643(.A1(new_n839_), .A2(new_n842_), .B1(new_n844_), .B2(new_n829_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n836_), .B1(new_n845_), .B2(new_n690_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n829_), .B1(new_n313_), .B2(new_n277_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n822_), .A2(new_n848_), .A3(new_n823_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n840_), .A2(new_n841_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n847_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n851_), .A2(KEYINPUT57), .A3(new_n630_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n809_), .B(new_n835_), .C1(new_n846_), .C2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n639_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n845_), .A2(new_n836_), .A3(new_n690_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n851_), .B2(new_n630_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n809_), .B1(new_n857_), .B2(new_n835_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n808_), .B1(new_n854_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n651_), .A2(new_n400_), .A3(new_n572_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(G113gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n310_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865_));
  INV_X1    g664(.A(new_n861_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n859_), .B2(new_n866_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n868_));
  NAND2_X1  g667(.A1(new_n857_), .A2(new_n835_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n639_), .ZN(new_n870_));
  AOI211_X1 g669(.A(new_n861_), .B(new_n868_), .C1(new_n870_), .C2(new_n808_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n867_), .A2(new_n309_), .A3(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n864_), .B1(new_n872_), .B2(new_n863_), .ZN(G1340gat));
  INV_X1    g672(.A(G120gat), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n874_), .A2(KEYINPUT60), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n643_), .B2(KEYINPUT60), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n862_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n867_), .A2(new_n643_), .A3(new_n871_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n874_), .ZN(G1341gat));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n862_), .A2(new_n880_), .A3(new_n329_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n867_), .A2(new_n639_), .A3(new_n871_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n880_), .ZN(G1342gat));
  INV_X1    g682(.A(G134gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n862_), .A2(new_n884_), .A3(new_n630_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n867_), .A2(new_n696_), .A3(new_n871_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n884_), .ZN(G1343gat));
  NOR4_X1   g686(.A1(new_n581_), .A2(new_n576_), .A3(new_n554_), .A4(new_n572_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n859_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n310_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G141gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n889_), .A2(new_n347_), .A3(new_n310_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1344gat));
  XNOR2_X1  g692(.A(KEYINPUT123), .B(G148gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n889_), .B2(new_n701_), .ZN(new_n895_));
  AND4_X1   g694(.A1(new_n701_), .A2(new_n859_), .A3(new_n888_), .A4(new_n894_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1345gat));
  NAND2_X1  g696(.A1(new_n889_), .A2(new_n329_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT61), .B(G155gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n899_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n889_), .A2(new_n329_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1346gat));
  INV_X1    g702(.A(G162gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n889_), .A2(new_n904_), .A3(new_n630_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n889_), .A2(new_n638_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n904_), .ZN(G1347gat));
  NAND2_X1  g706(.A1(new_n652_), .A2(new_n554_), .ZN(new_n908_));
  XOR2_X1   g707(.A(new_n908_), .B(KEYINPUT124), .Z(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  AOI211_X1 g709(.A(new_n475_), .B(new_n910_), .C1(new_n870_), .C2(new_n808_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n517_), .A3(new_n310_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n310_), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT125), .Z(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n475_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n870_), .A2(new_n808_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n484_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n918_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n912_), .B1(new_n919_), .B2(new_n920_), .ZN(G1348gat));
  AOI21_X1  g720(.A(G176gat), .B1(new_n911_), .B2(new_n701_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n860_), .A2(new_n475_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n910_), .A2(new_n485_), .A3(new_n643_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  NAND4_X1  g724(.A1(new_n859_), .A2(new_n581_), .A3(new_n329_), .A4(new_n909_), .ZN(new_n926_));
  INV_X1    g725(.A(G183gat), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n639_), .A2(new_n492_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n926_), .A2(new_n927_), .B1(new_n911_), .B2(new_n928_), .ZN(G1350gat));
  NAND2_X1  g728(.A1(new_n911_), .A2(new_n638_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(G190gat), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n911_), .A2(new_n513_), .A3(new_n514_), .A4(new_n630_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1351gat));
  NAND3_X1  g732(.A1(new_n475_), .A2(new_n576_), .A3(new_n646_), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n934_), .A2(KEYINPUT126), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(KEYINPUT126), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n935_), .A2(new_n554_), .A3(new_n936_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n859_), .A2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938_), .B2(new_n310_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n937_), .ZN(new_n940_));
  NOR4_X1   g739(.A1(new_n860_), .A2(new_n416_), .A3(new_n309_), .A4(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n415_), .A2(new_n417_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n859_), .A2(new_n944_), .A3(new_n701_), .A4(new_n937_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(KEYINPUT127), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n945_), .A2(KEYINPUT127), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n859_), .A2(new_n701_), .A3(new_n937_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(G204gat), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n946_), .B1(new_n947_), .B2(new_n949_), .ZN(G1353gat));
  XNOR2_X1  g749(.A(KEYINPUT63), .B(G211gat), .ZN(new_n951_));
  NOR4_X1   g750(.A1(new_n860_), .A2(new_n639_), .A3(new_n940_), .A4(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n938_), .A2(new_n329_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n952_), .B1(new_n953_), .B2(new_n954_), .ZN(G1354gat));
  NAND3_X1  g754(.A1(new_n938_), .A2(new_n408_), .A3(new_n630_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n860_), .A2(new_n696_), .A3(new_n940_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n957_), .B2(new_n408_), .ZN(G1355gat));
endmodule


