//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n972_, new_n973_, new_n974_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n984_, new_n985_;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT66), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT66), .B1(new_n211_), .B2(new_n213_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n209_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(KEYINPUT8), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT67), .B1(new_n211_), .B2(new_n213_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(new_n208_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT67), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n221_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n223_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT64), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n205_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n212_), .B1(G99gat), .B2(G106gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT66), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n219_), .B1(new_n218_), .B2(KEYINPUT9), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT9), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n217_), .A2(KEYINPUT65), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT65), .B1(new_n217_), .B2(new_n245_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n244_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n237_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT70), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n237_), .A2(new_n243_), .A3(new_n248_), .A4(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n229_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G29gat), .B(G36gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G43gat), .B(G50gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT15), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n202_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G232gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT34), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT35), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT15), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n256_), .B(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n234_), .A2(KEYINPUT64), .A3(new_n235_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n232_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n205_), .A2(new_n269_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n251_), .B1(new_n270_), .B2(new_n248_), .ZN(new_n271_));
  AND4_X1   g070(.A1(new_n251_), .A2(new_n237_), .A3(new_n243_), .A4(new_n248_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n266_), .B1(new_n273_), .B2(new_n229_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n229_), .A2(new_n256_), .A3(new_n249_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI22_X1  g075(.A1(new_n258_), .A2(new_n264_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n261_), .A2(new_n262_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n250_), .A2(new_n252_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(new_n209_), .A3(new_n226_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n220_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n283_), .A2(KEYINPUT8), .B1(new_n216_), .B2(new_n222_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n257_), .B1(new_n279_), .B2(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n285_), .A2(new_n202_), .A3(new_n275_), .A4(new_n263_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n277_), .A2(new_n278_), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G190gat), .B(G218gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G134gat), .B(G162gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n290_), .A2(KEYINPUT36), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n290_), .A2(KEYINPUT36), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n285_), .A2(KEYINPUT73), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n296_), .A2(new_n263_), .B1(new_n285_), .B2(new_n275_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n286_), .A2(new_n278_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n294_), .B(new_n295_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n295_), .B1(new_n287_), .B2(new_n294_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n293_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT37), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT37), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n304_), .B(new_n293_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT75), .B(G8gat), .Z(new_n307_));
  INV_X1    g106(.A(G1gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT14), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G15gat), .B(G22gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G1gat), .B(G8gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G231gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G64gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G57gat), .ZN(new_n320_));
  INV_X1    g119(.A(G57gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(G64gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(KEYINPUT68), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G57gat), .B(G64gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT11), .B1(new_n324_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT69), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n323_), .A2(KEYINPUT68), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n326_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT11), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G71gat), .B(G78gat), .Z(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n331_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT69), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(KEYINPUT11), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n329_), .A2(new_n333_), .A3(new_n334_), .A4(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(new_n334_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n335_), .B2(KEYINPUT11), .ZN(new_n340_));
  AOI211_X1 g139(.A(KEYINPUT69), .B(new_n332_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n318_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT17), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G183gat), .B(G211gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT77), .ZN(new_n347_));
  XOR2_X1   g146(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G127gat), .B(G155gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n344_), .A2(new_n345_), .A3(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(KEYINPUT17), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n344_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n306_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n358_));
  NAND2_X1  g157(.A1(new_n283_), .A2(KEYINPUT8), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n359_), .A2(new_n223_), .B1(new_n248_), .B2(new_n270_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(new_n343_), .B2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(G230gat), .A2(G233gat), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n343_), .B2(new_n360_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n253_), .A2(KEYINPUT12), .A3(new_n338_), .A4(new_n342_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT72), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT72), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n361_), .A2(new_n363_), .A3(new_n364_), .A4(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n343_), .B(new_n360_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n362_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G120gat), .B(G148gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT5), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G176gat), .B(G204gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n369_), .A2(new_n371_), .A3(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n377_), .A2(KEYINPUT13), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT13), .B1(new_n377_), .B2(new_n379_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n357_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G113gat), .B(G141gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G169gat), .B(G197gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n314_), .A2(new_n315_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n256_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n256_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n388_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n389_), .A2(new_n256_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(KEYINPUT78), .A3(new_n390_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G229gat), .A2(G233gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT79), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n395_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n400_));
  INV_X1    g199(.A(new_n397_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n316_), .A2(new_n257_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n390_), .A3(new_n397_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT80), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n387_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n400_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n408_));
  AOI211_X1 g207(.A(KEYINPUT79), .B(new_n397_), .C1(new_n393_), .C2(new_n395_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n406_), .B(new_n387_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT98), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n414_));
  INV_X1    g213(.A(G155gat), .ZN(new_n415_));
  INV_X1    g214(.A(G162gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT1), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .A4(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n418_), .A2(KEYINPUT1), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT85), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G141gat), .A2(G148gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(G141gat), .A2(G148gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n417_), .A2(new_n421_), .A3(new_n418_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT87), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n417_), .A2(new_n435_), .A3(new_n421_), .A4(new_n418_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n428_), .B(KEYINPUT2), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT3), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n430_), .A2(KEYINPUT86), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n430_), .A2(KEYINPUT86), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT3), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n437_), .A2(new_n438_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n438_), .B1(new_n437_), .B2(new_n444_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n432_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G127gat), .B(G134gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT82), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G113gat), .B(G120gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  NAND2_X1  g250(.A1(new_n447_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n449_), .B(new_n450_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n453_), .B(new_n432_), .C1(new_n446_), .C2(new_n445_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n452_), .A2(KEYINPUT4), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n447_), .A2(new_n456_), .A3(new_n451_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G225gat), .A2(G233gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n413_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G1gat), .B(G29gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT97), .B(G85gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT0), .B(G57gat), .ZN(new_n464_));
  XOR2_X1   g263(.A(new_n463_), .B(new_n464_), .Z(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n452_), .A2(new_n454_), .A3(KEYINPUT4), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n467_), .A2(KEYINPUT98), .A3(new_n458_), .A4(new_n457_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n458_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n452_), .A2(new_n454_), .A3(new_n469_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n460_), .A2(new_n466_), .A3(new_n468_), .A4(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n452_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n457_), .A2(new_n469_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n472_), .B(new_n465_), .C1(new_n455_), .C2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(G8gat), .B(G36gat), .Z(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G64gat), .B(G92gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G226gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT19), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT93), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT95), .ZN(new_n485_));
  INV_X1    g284(.A(G197gat), .ZN(new_n486_));
  INV_X1    g285(.A(G204gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G197gat), .A2(G204gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT21), .A3(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G211gat), .B(G218gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT90), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(G218gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G211gat), .ZN(new_n494_));
  INV_X1    g293(.A(G211gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G218gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(G197gat), .A2(G204gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G197gat), .A2(G204gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n497_), .A2(new_n500_), .A3(new_n501_), .A4(KEYINPUT21), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n492_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n497_), .B1(KEYINPUT21), .B2(new_n500_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT21), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G176gat), .ZN(new_n509_));
  INV_X1    g308(.A(G169gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT22), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT22), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G169gat), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n511_), .A2(new_n513_), .A3(KEYINPUT94), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT94), .B1(new_n511_), .B2(new_n513_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n509_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G183gat), .A2(G190gat), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(G183gat), .A2(G190gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G169gat), .A2(G176gat), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n516_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT25), .B(G183gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G190gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT24), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(G169gat), .B2(G176gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n510_), .A2(new_n509_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n526_), .A2(new_n527_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n528_), .A2(new_n510_), .A3(new_n509_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n485_), .B(new_n508_), .C1(new_n525_), .C2(new_n535_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n516_), .A2(new_n524_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n492_), .A2(new_n502_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT95), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT81), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n533_), .A2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n532_), .A2(new_n519_), .A3(KEYINPUT81), .A4(new_n521_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n531_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n512_), .A2(new_n510_), .A3(new_n509_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n522_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT20), .B1(new_n548_), .B2(new_n508_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n484_), .B1(new_n540_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n483_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n548_), .A2(new_n508_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n481_), .B1(new_n551_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n481_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n549_), .B1(new_n539_), .B2(new_n536_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n556_), .B(new_n559_), .C1(new_n560_), .C2(new_n484_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n467_), .A2(new_n469_), .A3(new_n457_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n563_), .A2(KEYINPUT33), .A3(new_n472_), .A4(new_n465_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n471_), .A2(new_n476_), .A3(new_n562_), .A4(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n540_), .A2(new_n484_), .A3(new_n550_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n554_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(KEYINPUT32), .A3(new_n559_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n559_), .A2(KEYINPUT32), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n556_), .B(new_n571_), .C1(new_n560_), .C2(new_n484_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n474_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n465_), .B1(new_n563_), .B2(new_n472_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n570_), .B(new_n572_), .C1(new_n573_), .C2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n565_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT89), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT29), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n432_), .B(new_n578_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT28), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n437_), .A2(new_n444_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT88), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n437_), .A2(new_n438_), .A3(new_n444_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT28), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n578_), .A4(new_n432_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G22gat), .B(G50gat), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n580_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n580_), .B2(new_n586_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n577_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n587_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n431_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n585_), .B1(new_n594_), .B2(new_n578_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n579_), .A2(KEYINPUT28), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n591_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n580_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(KEYINPUT89), .A3(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n508_), .B1(new_n594_), .B2(new_n578_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G228gat), .A2(G233gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n447_), .A2(KEYINPUT29), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n601_), .A3(new_n508_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT91), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G78gat), .B(G106gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n590_), .A2(new_n599_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT91), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n601_), .B1(new_n604_), .B2(new_n508_), .ZN(new_n611_));
  AOI211_X1 g410(.A(new_n602_), .B(new_n538_), .C1(new_n447_), .C2(KEYINPUT29), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n603_), .A2(KEYINPUT91), .A3(new_n605_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n614_), .A3(new_n607_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n607_), .A2(KEYINPUT92), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n611_), .A2(new_n612_), .A3(new_n617_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n597_), .A2(new_n598_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n609_), .A2(new_n615_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n576_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n590_), .A2(new_n599_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n606_), .A2(new_n608_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n615_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n618_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n573_), .A2(new_n574_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT27), .B1(new_n558_), .B2(new_n561_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n567_), .B1(new_n560_), .B2(new_n484_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(new_n559_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n569_), .A2(KEYINPUT99), .A3(new_n481_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n561_), .A2(KEYINPUT27), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n630_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n628_), .A2(new_n629_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n623_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n453_), .B(KEYINPUT83), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G71gat), .B(G99gat), .ZN(new_n641_));
  INV_X1    g440(.A(G43gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n548_), .B(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n640_), .B(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G227gat), .A2(G233gat), .ZN(new_n646_));
  INV_X1    g445(.A(G15gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT30), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT31), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n645_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n639_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n629_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n622_), .B2(new_n637_), .ZN(new_n657_));
  AND4_X1   g456(.A1(new_n656_), .A2(new_n637_), .A3(new_n626_), .A4(new_n627_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n412_), .B1(new_n653_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n384_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n629_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n308_), .A3(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT101), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n666_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n653_), .A2(new_n659_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n287_), .A2(new_n292_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n294_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n295_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(new_n673_), .B2(new_n299_), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT102), .B1(new_n669_), .B2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n356_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n669_), .A2(KEYINPUT102), .A3(new_n674_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n382_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(new_n412_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G1gat), .B1(new_n681_), .B2(new_n629_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n667_), .A2(new_n668_), .A3(new_n682_), .ZN(G1324gat));
  INV_X1    g482(.A(new_n637_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n662_), .A2(new_n307_), .A3(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n676_), .A2(new_n680_), .A3(new_n684_), .A4(new_n677_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT39), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(G8gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G8gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n690_), .B(new_n692_), .ZN(G1325gat));
  NAND4_X1  g492(.A1(new_n676_), .A2(new_n680_), .A3(new_n651_), .A4(new_n677_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G15gat), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(KEYINPUT105), .A3(G15gat), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n661_), .A2(G15gat), .A3(new_n652_), .ZN(new_n702_));
  OR3_X1    g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(G1326gat));
  OR3_X1    g502(.A1(new_n661_), .A2(G22gat), .A3(new_n622_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G22gat), .B1(new_n681_), .B2(new_n622_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(KEYINPUT42), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(KEYINPUT42), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(G1327gat));
  NOR4_X1   g507(.A1(new_n380_), .A2(new_n381_), .A3(new_n674_), .A4(new_n355_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n660_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT109), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n660_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  OR3_X1    g513(.A1(new_n714_), .A2(G29gat), .A3(new_n629_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716_));
  INV_X1    g515(.A(new_n306_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT43), .B(new_n717_), .C1(new_n653_), .C2(new_n659_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n674_), .A2(new_n304_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n305_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n303_), .A2(KEYINPUT106), .A3(new_n305_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n653_), .A2(new_n659_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT107), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n651_), .B1(new_n623_), .B2(new_n638_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n637_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT100), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n622_), .A2(new_n656_), .A3(new_n637_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n654_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n303_), .A2(KEYINPUT106), .A3(new_n305_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT106), .B1(new_n303_), .B2(new_n305_), .ZN(new_n733_));
  OAI22_X1  g532(.A1(new_n727_), .A2(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(KEYINPUT43), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n718_), .B1(new_n726_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n680_), .A2(new_n356_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n716_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n718_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n734_), .A2(new_n735_), .A3(KEYINPUT43), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n735_), .B1(new_n734_), .B2(KEYINPUT43), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n738_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(KEYINPUT44), .A3(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n739_), .A2(new_n745_), .A3(new_n663_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n746_), .A2(KEYINPUT108), .A3(G29gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT108), .B1(new_n746_), .B2(G29gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n715_), .B1(new_n747_), .B2(new_n748_), .ZN(G1328gat));
  NAND3_X1  g548(.A1(new_n739_), .A2(new_n745_), .A3(new_n684_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G36gat), .ZN(new_n751_));
  INV_X1    g550(.A(new_n714_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n637_), .A2(G36gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT45), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n756_), .A3(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n751_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n751_), .A2(new_n758_), .A3(KEYINPUT46), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1329gat));
  NAND4_X1  g562(.A1(new_n739_), .A2(new_n745_), .A3(G43gat), .A4(new_n651_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n642_), .B1(new_n714_), .B2(new_n652_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g566(.A1(new_n739_), .A2(new_n745_), .A3(new_n628_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G50gat), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n622_), .A2(G50gat), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT110), .Z(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n714_), .B2(new_n771_), .ZN(G1331gat));
  NAND2_X1  g571(.A1(new_n403_), .A2(new_n406_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n387_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n410_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n382_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n678_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G57gat), .B1(new_n778_), .B2(new_n629_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n776_), .B1(new_n653_), .B2(new_n659_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n780_), .A2(new_n679_), .A3(new_n357_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n321_), .A3(new_n663_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(G1332gat));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n319_), .A3(new_n684_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT48), .ZN(new_n785_));
  INV_X1    g584(.A(new_n778_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n684_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n787_), .B2(G64gat), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT48), .B(new_n319_), .C1(new_n786_), .C2(new_n684_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n784_), .B1(new_n788_), .B2(new_n789_), .ZN(G1333gat));
  INV_X1    g589(.A(G71gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n781_), .A2(new_n791_), .A3(new_n651_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G71gat), .B1(new_n778_), .B2(new_n652_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(KEYINPUT49), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(KEYINPUT49), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n792_), .B1(new_n794_), .B2(new_n795_), .ZN(G1334gat));
  INV_X1    g595(.A(G78gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n781_), .A2(new_n797_), .A3(new_n628_), .ZN(new_n798_));
  OAI21_X1  g597(.A(G78gat), .B1(new_n778_), .B2(new_n622_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n799_), .A2(new_n800_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(G1335gat));
  NAND2_X1  g602(.A1(new_n777_), .A2(new_n356_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n737_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(G85gat), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n629_), .A2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT112), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n808_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n382_), .A2(new_n674_), .A3(new_n355_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n780_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n806_), .B1(new_n811_), .B2(new_n629_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT113), .Z(G1336gat));
  INV_X1    g613(.A(new_n811_), .ZN(new_n815_));
  AOI21_X1  g614(.A(G92gat), .B1(new_n815_), .B2(new_n684_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n684_), .A2(G92gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT114), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n805_), .B2(new_n818_), .ZN(G1337gat));
  AND3_X1   g618(.A1(new_n815_), .A2(new_n269_), .A3(new_n651_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n805_), .A2(new_n651_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(G99gat), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1338gat));
  NAND3_X1  g623(.A1(new_n815_), .A2(new_n205_), .A3(new_n628_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n804_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n743_), .A2(new_n628_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n827_), .A2(new_n828_), .A3(G106gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n827_), .B2(G106gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n825_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT53), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n833_), .B(new_n825_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1339gat));
  INV_X1    g634(.A(G113gat), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n343_), .A2(new_n360_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n361_), .A2(new_n364_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n362_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n361_), .A2(new_n363_), .A3(new_n364_), .A4(KEYINPUT55), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n366_), .A2(new_n843_), .A3(new_n368_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n366_), .A2(KEYINPUT115), .A3(new_n843_), .A4(new_n368_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n376_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n404_), .A2(new_n390_), .A3(new_n401_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n774_), .B(new_n851_), .C1(new_n396_), .C2(new_n401_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n379_), .A2(new_n410_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n378_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n849_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n837_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n848_), .A2(new_n376_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT56), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n859_), .A2(KEYINPUT118), .A3(new_n850_), .A4(new_n853_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n854_), .A2(new_n856_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n717_), .B1(new_n863_), .B2(KEYINPUT58), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867_));
  AOI211_X1 g666(.A(new_n867_), .B(new_n378_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n849_), .B1(new_n868_), .B2(KEYINPUT117), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n870_), .B2(KEYINPUT56), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n379_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n412_), .B1(new_n858_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n377_), .A2(new_n379_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n410_), .A2(new_n852_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n869_), .A2(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n866_), .B1(new_n876_), .B2(new_n302_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n874_), .A2(new_n875_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n855_), .A2(KEYINPUT116), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT56), .B1(new_n879_), .B2(new_n870_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n872_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n776_), .B1(new_n881_), .B2(new_n855_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(KEYINPUT57), .A3(new_n674_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n865_), .A2(new_n877_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n356_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n383_), .B2(new_n776_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n357_), .A2(new_n382_), .A3(new_n888_), .A4(new_n412_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n886_), .A2(new_n891_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n629_), .B(new_n652_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n836_), .B1(new_n894_), .B2(new_n412_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(KEYINPUT120), .B(new_n836_), .C1(new_n894_), .C2(new_n412_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n892_), .A2(new_n893_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n890_), .B1(new_n885_), .B2(new_n356_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n893_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT59), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n900_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n412_), .A2(new_n836_), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n897_), .A2(new_n898_), .B1(new_n904_), .B2(new_n905_), .ZN(G1340gat));
  NAND3_X1  g705(.A1(new_n900_), .A2(new_n679_), .A3(new_n903_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G120gat), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G120gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n382_), .A2(KEYINPUT60), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(G120gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n908_), .B1(new_n894_), .B2(new_n912_), .ZN(G1341gat));
  INV_X1    g712(.A(new_n894_), .ZN(new_n914_));
  AOI21_X1  g713(.A(G127gat), .B1(new_n914_), .B2(new_n355_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n356_), .A2(KEYINPUT122), .ZN(new_n916_));
  MUX2_X1   g715(.A(KEYINPUT122), .B(new_n916_), .S(G127gat), .Z(new_n917_));
  AOI21_X1  g716(.A(new_n915_), .B1(new_n904_), .B2(new_n917_), .ZN(G1342gat));
  NAND3_X1  g717(.A1(new_n900_), .A2(new_n306_), .A3(new_n903_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G134gat), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n674_), .A2(G134gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n894_), .B2(new_n921_), .ZN(G1343gat));
  NAND4_X1  g721(.A1(new_n628_), .A2(new_n652_), .A3(new_n663_), .A4(new_n637_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n901_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n776_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n679_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g727(.A1(new_n924_), .A2(new_n355_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT61), .B(G155gat), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1346gat));
  AOI21_X1  g730(.A(G162gat), .B1(new_n924_), .B2(new_n302_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n416_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT123), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n924_), .B2(new_n934_), .ZN(G1347gat));
  NOR3_X1   g734(.A1(new_n654_), .A2(new_n628_), .A3(new_n637_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n937_), .B1(new_n886_), .B2(new_n891_), .ZN(new_n938_));
  AOI211_X1 g737(.A(KEYINPUT62), .B(new_n510_), .C1(new_n938_), .C2(new_n776_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n776_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(G169gat), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n938_), .B(new_n776_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n939_), .B1(new_n942_), .B2(new_n943_), .ZN(G1348gat));
  NAND2_X1  g743(.A1(new_n938_), .A2(new_n679_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g745(.A1(new_n883_), .A2(new_n674_), .ZN(new_n947_));
  AOI22_X1  g746(.A1(new_n947_), .A2(new_n866_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n355_), .B1(new_n948_), .B2(new_n884_), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n355_), .B(new_n936_), .C1(new_n949_), .C2(new_n890_), .ZN(new_n950_));
  INV_X1    g749(.A(G183gat), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n953_));
  INV_X1    g752(.A(new_n526_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n938_), .A2(new_n954_), .A3(new_n355_), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n952_), .A2(new_n953_), .A3(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n953_), .B1(new_n952_), .B2(new_n955_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1350gat));
  INV_X1    g757(.A(new_n938_), .ZN(new_n959_));
  OAI21_X1  g758(.A(G190gat), .B1(new_n959_), .B2(new_n717_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n938_), .A2(new_n527_), .A3(new_n302_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1351gat));
  NOR4_X1   g761(.A1(new_n622_), .A2(new_n663_), .A3(new_n637_), .A4(new_n651_), .ZN(new_n963_));
  OAI211_X1 g762(.A(KEYINPUT125), .B(new_n963_), .C1(new_n949_), .C2(new_n890_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965_));
  INV_X1    g764(.A(new_n963_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n901_), .B2(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n964_), .A2(new_n967_), .ZN(new_n968_));
  AOI21_X1  g767(.A(G197gat), .B1(new_n968_), .B2(new_n776_), .ZN(new_n969_));
  AOI211_X1 g768(.A(new_n486_), .B(new_n412_), .C1(new_n964_), .C2(new_n967_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1352gat));
  NAND2_X1  g770(.A1(new_n968_), .A2(new_n679_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n972_), .A2(G204gat), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n968_), .A2(new_n487_), .A3(new_n679_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n973_), .A2(new_n974_), .ZN(G1353gat));
  AOI21_X1  g774(.A(new_n356_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n968_), .A2(new_n976_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(KEYINPUT126), .ZN(new_n979_));
  INV_X1    g778(.A(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n977_), .A2(new_n980_), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n968_), .A2(new_n979_), .A3(new_n976_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n981_), .A2(new_n982_), .ZN(G1354gat));
  NAND3_X1  g782(.A1(new_n968_), .A2(new_n493_), .A3(new_n302_), .ZN(new_n984_));
  AOI21_X1  g783(.A(new_n717_), .B1(new_n964_), .B2(new_n967_), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n984_), .B1(new_n493_), .B2(new_n985_), .ZN(G1355gat));
endmodule


