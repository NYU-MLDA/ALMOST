//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT18), .B(G64gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT19), .ZN(new_n207_));
  INV_X1    g006(.A(G204gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G197gat), .ZN(new_n209_));
  INV_X1    g008(.A(G197gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G204gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT21), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT21), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n209_), .A2(new_n211_), .A3(new_n215_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n213_), .A2(KEYINPUT87), .A3(new_n214_), .A4(new_n216_), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n213_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219_));
  INV_X1    g018(.A(new_n214_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n215_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n217_), .B1(new_n218_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT22), .B(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n229_), .B(new_n230_), .C1(G183gat), .C2(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n226_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT26), .B(G190gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT25), .B(G183gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT89), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT89), .ZN(new_n238_));
  INV_X1    g037(.A(G183gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(KEYINPUT25), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(G183gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n238_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n235_), .B1(new_n237_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G169gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n225_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT24), .A3(new_n232_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(new_n245_), .A3(new_n225_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n247_), .A2(new_n229_), .A3(new_n230_), .A4(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n233_), .B1(new_n244_), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n223_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n226_), .A2(KEYINPUT79), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT79), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n224_), .A2(new_n254_), .A3(new_n225_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n253_), .A2(new_n232_), .A3(new_n231_), .A4(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT76), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n239_), .B2(KEYINPUT25), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n234_), .B(new_n258_), .C1(new_n236_), .C2(new_n257_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n249_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT78), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n249_), .A2(new_n229_), .A3(KEYINPUT78), .A4(new_n230_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n247_), .B(KEYINPUT77), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n256_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n256_), .B(KEYINPUT80), .C1(new_n264_), .C2(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n252_), .B1(new_n270_), .B2(new_n223_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n207_), .B1(new_n271_), .B2(KEYINPUT20), .ZN(new_n272_));
  INV_X1    g071(.A(new_n223_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n268_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n223_), .A2(new_n251_), .ZN(new_n275_));
  AND4_X1   g074(.A1(KEYINPUT20), .A2(new_n274_), .A3(new_n207_), .A4(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n205_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n207_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n274_), .A2(KEYINPUT20), .A3(new_n278_), .A4(new_n275_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT93), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n251_), .A2(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n233_), .B(KEYINPUT93), .C1(new_n244_), .C2(new_n250_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n273_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT94), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n269_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT77), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n247_), .B(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n291_), .A2(new_n262_), .A3(new_n263_), .A4(new_n259_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT80), .B1(new_n292_), .B2(new_n256_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n223_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n284_), .A2(KEYINPUT94), .A3(new_n285_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n288_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n280_), .B1(new_n296_), .B2(new_n207_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n277_), .B(KEYINPUT27), .C1(new_n297_), .C2(new_n205_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT96), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n272_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n276_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n205_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n277_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n295_), .A2(new_n294_), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT94), .B1(new_n284_), .B2(new_n285_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n207_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n279_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n303_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n312_), .A2(KEYINPUT96), .A3(KEYINPUT27), .A4(new_n277_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n300_), .A2(new_n307_), .A3(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G141gat), .B(G148gat), .Z(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT1), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT82), .ZN(new_n320_));
  OR2_X1    g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n322_), .A3(KEYINPUT1), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n318_), .A2(KEYINPUT1), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n317_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n327_), .B1(new_n328_), .B2(KEYINPUT83), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT83), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n330_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(KEYINPUT83), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n321_), .B(new_n318_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n326_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT85), .B1(new_n337_), .B2(KEYINPUT29), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT85), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n326_), .A2(new_n336_), .A3(new_n339_), .A4(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n338_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n343_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n316_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n338_), .A2(new_n341_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n342_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n338_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n315_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT88), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT86), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n337_), .B2(KEYINPUT29), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n223_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(new_n356_), .A3(new_n223_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n351_), .A2(new_n352_), .A3(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n354_), .A2(new_n356_), .A3(new_n223_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n356_), .B1(new_n354_), .B2(new_n223_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT88), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n358_), .A2(new_n352_), .A3(new_n359_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n350_), .A2(new_n346_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n362_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n363_), .B1(new_n362_), .B2(new_n368_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G15gat), .B(G43gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT81), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT31), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT30), .B1(new_n289_), .B2(new_n293_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G127gat), .B(G134gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n268_), .A2(new_n378_), .A3(new_n269_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n374_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n377_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n373_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n377_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n379_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n378_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n374_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n373_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  AND3_X1   g191(.A1(new_n382_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n382_), .B2(new_n389_), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n369_), .A2(new_n370_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n363_), .ZN(new_n396_));
  AOI211_X1 g195(.A(KEYINPUT88), .B(new_n360_), .C1(new_n346_), .C2(new_n350_), .ZN(new_n397_));
  AND4_X1   g196(.A1(new_n367_), .A2(new_n346_), .A3(new_n366_), .A4(new_n350_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n392_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n389_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n388_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n400_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n382_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n362_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n399_), .A2(new_n403_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n395_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n337_), .A2(new_n383_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n326_), .A2(new_n336_), .A3(new_n377_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(KEYINPUT4), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n411_), .B(KEYINPUT90), .Z(new_n412_));
  OAI211_X1 g211(.A(new_n410_), .B(new_n412_), .C1(KEYINPUT4), .C2(new_n408_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n409_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n414_), .A2(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417_));
  INV_X1    g216(.A(G85gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT0), .B(G57gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n416_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT95), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n413_), .A2(new_n415_), .A3(new_n421_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT95), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n416_), .A2(new_n426_), .A3(new_n422_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n424_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n314_), .A2(new_n407_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n428_), .B(new_n432_), .C1(new_n297_), .C2(new_n431_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n425_), .B(KEYINPUT33), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n414_), .B(KEYINPUT91), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n412_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n410_), .B1(KEYINPUT4), .B2(new_n408_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n436_), .B(new_n422_), .C1(new_n412_), .C2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n434_), .A2(new_n304_), .A3(new_n277_), .A4(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n393_), .A2(new_n394_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n399_), .A2(new_n405_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n430_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT10), .B(G99gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT64), .B1(new_n445_), .B2(G106gat), .ZN(new_n446_));
  INV_X1    g245(.A(G99gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT10), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT10), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(G99gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT64), .ZN(new_n452_));
  INV_X1    g251(.A(G106gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n446_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n461_), .A2(KEYINPUT9), .ZN(new_n462_));
  OR2_X1    g261(.A1(G85gat), .A2(G92gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(KEYINPUT9), .A3(new_n461_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n460_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT66), .B1(new_n455_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT8), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT7), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n447_), .A3(new_n453_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n458_), .A3(new_n459_), .A4(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n463_), .A2(new_n461_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n467_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n465_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n446_), .A2(new_n454_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT66), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n466_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G57gat), .B(G64gat), .ZN(new_n483_));
  INV_X1    g282(.A(G71gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT65), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G71gat), .ZN(new_n487_));
  INV_X1    g286(.A(G78gat), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT11), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n486_), .A2(G71gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n484_), .A2(KEYINPUT65), .ZN(new_n494_));
  OAI21_X1  g293(.A(G78gat), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT11), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n483_), .B1(new_n492_), .B2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(KEYINPUT11), .A3(new_n496_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n483_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n482_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n481_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n491_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n500_), .B1(new_n504_), .B2(new_n499_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n499_), .A2(new_n500_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n474_), .A2(new_n475_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n482_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G230gat), .A2(G233gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n508_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n503_), .A2(new_n509_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n510_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n507_), .A2(new_n508_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n498_), .A2(new_n501_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n475_), .ZN(new_n516_));
  OAI22_X1  g315(.A1(new_n455_), .A2(new_n465_), .B1(new_n516_), .B2(new_n473_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n513_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n512_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT67), .B(G204gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT5), .B(G176gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G120gat), .B(G148gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n520_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n512_), .A2(new_n519_), .A3(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(KEYINPUT68), .B2(KEYINPUT13), .ZN(new_n530_));
  NOR2_X1   g329(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n531_));
  AND2_X1   g330(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n527_), .B(new_n528_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536_));
  INV_X1    g335(.A(G1gat), .ZN(new_n537_));
  INV_X1    g336(.A(G8gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT14), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G1gat), .B(G8gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G29gat), .B(G36gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G43gat), .B(G50gat), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n542_), .A2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT69), .B(KEYINPUT15), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n549_), .B(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n552_), .B2(new_n542_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n542_), .B(new_n549_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G169gat), .B(G197gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT75), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n559_), .B(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n535_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n444_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n542_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(new_n515_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT74), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT16), .B(G183gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT17), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(KEYINPUT17), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n570_), .A2(new_n571_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n572_), .A2(new_n578_), .A3(new_n579_), .A4(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n579_), .A2(KEYINPUT73), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(KEYINPUT73), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n570_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(KEYINPUT36), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n481_), .A2(new_n552_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT35), .Z(new_n595_));
  OAI211_X1 g394(.A(new_n592_), .B(new_n595_), .C1(new_n549_), .C2(new_n517_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n592_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT70), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n517_), .A2(new_n549_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT70), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n592_), .B2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n594_), .A2(KEYINPUT35), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n591_), .B(new_n596_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT71), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n603_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n596_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT71), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n591_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n589_), .B(KEYINPUT36), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n612_));
  AND4_X1   g411(.A1(KEYINPUT37), .A2(new_n605_), .A3(new_n610_), .A4(new_n612_), .ZN(new_n613_));
  OR3_X1    g412(.A1(new_n606_), .A2(KEYINPUT72), .A3(new_n607_), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT72), .B1(new_n606_), .B2(new_n607_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n611_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT37), .B1(new_n616_), .B2(new_n604_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n567_), .A2(new_n586_), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(new_n537_), .A3(new_n428_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT38), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n604_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI211_X1 g422(.A(new_n585_), .B(new_n623_), .C1(new_n430_), .C2(new_n443_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n566_), .B(KEYINPUT97), .Z(new_n625_));
  AND2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(new_n428_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n621_), .B1(new_n537_), .B2(new_n627_), .ZN(G1324gat));
  NAND3_X1  g427(.A1(new_n300_), .A2(new_n307_), .A3(new_n313_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n619_), .A2(new_n538_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n626_), .A2(new_n629_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(G8gat), .ZN(new_n633_));
  AOI211_X1 g432(.A(KEYINPUT39), .B(new_n538_), .C1(new_n626_), .C2(new_n629_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(G1325gat));
  INV_X1    g436(.A(G15gat), .ZN(new_n638_));
  INV_X1    g437(.A(new_n441_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n626_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT41), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n619_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  INV_X1    g443(.A(new_n442_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n626_), .B2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT42), .Z(new_n647_));
  NAND3_X1  g446(.A1(new_n619_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1327gat));
  NOR2_X1   g448(.A1(new_n622_), .A2(new_n586_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n567_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G29gat), .B1(new_n651_), .B2(new_n428_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n618_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT98), .B1(new_n613_), .B2(new_n617_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT43), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n444_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n444_), .B2(new_n653_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n625_), .B(new_n585_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n655_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n629_), .B1(new_n406_), .B2(new_n395_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(new_n429_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n664_), .B2(new_n618_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n444_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n659_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n667_), .A2(new_n625_), .A3(new_n585_), .A4(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n660_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n428_), .A2(G29gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n652_), .B1(new_n670_), .B2(new_n671_), .ZN(G1328gat));
  NAND3_X1  g471(.A1(new_n660_), .A2(new_n669_), .A3(new_n629_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G36gat), .ZN(new_n674_));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n629_), .A2(KEYINPUT100), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n629_), .A2(KEYINPUT100), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n567_), .A2(new_n675_), .A3(new_n650_), .A4(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n674_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n674_), .A2(KEYINPUT46), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1329gat));
  NAND2_X1  g486(.A1(new_n567_), .A2(new_n650_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n688_), .A2(G43gat), .A3(new_n441_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n660_), .A2(new_n669_), .A3(new_n639_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(G43gat), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT47), .B(new_n689_), .C1(new_n690_), .C2(G43gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1330gat));
  NAND3_X1  g494(.A1(new_n660_), .A2(new_n669_), .A3(new_n645_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G50gat), .ZN(new_n697_));
  OR3_X1    g496(.A1(new_n688_), .A2(G50gat), .A3(new_n442_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT102), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(new_n701_), .A3(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1331gat));
  INV_X1    g502(.A(new_n565_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n534_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n624_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(G57gat), .A3(new_n428_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT103), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n444_), .A2(new_n705_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n709_), .A2(new_n585_), .A3(new_n653_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n428_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n708_), .A2(new_n711_), .ZN(G1332gat));
  INV_X1    g511(.A(G64gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n706_), .B2(new_n679_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT48), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n710_), .A2(new_n713_), .A3(new_n679_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1333gat));
  NAND3_X1  g516(.A1(new_n710_), .A2(new_n484_), .A3(new_n639_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n484_), .B1(new_n706_), .B2(new_n639_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT49), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n719_), .A2(new_n720_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT104), .B(new_n718_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1334gat));
  AOI21_X1  g526(.A(new_n488_), .B1(new_n706_), .B2(new_n645_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n710_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n645_), .A2(new_n488_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT106), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n730_), .B1(new_n731_), .B2(new_n733_), .ZN(G1335gat));
  AND3_X1   g533(.A1(new_n444_), .A2(new_n650_), .A3(new_n705_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n428_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n705_), .A2(new_n585_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT107), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n667_), .A2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n429_), .A2(new_n418_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1336gat));
  AOI21_X1  g540(.A(G92gat), .B1(new_n735_), .B2(new_n629_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n679_), .A2(G92gat), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT108), .Z(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n744_), .B2(new_n739_), .ZN(G1337gat));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(KEYINPUT51), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n735_), .A2(new_n451_), .A3(new_n639_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT109), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n667_), .A2(new_n639_), .A3(new_n738_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G99gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n747_), .B1(new_n749_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n746_), .A2(KEYINPUT51), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT111), .Z(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n752_), .B(new_n755_), .ZN(G1338gat));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n667_), .A2(new_n645_), .A3(new_n738_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n757_), .B1(new_n759_), .B2(new_n453_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n735_), .A2(new_n453_), .A3(new_n645_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT112), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT53), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n760_), .A2(new_n762_), .A3(new_n766_), .A4(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1339gat));
  NOR3_X1   g567(.A1(new_n629_), .A2(new_n429_), .A3(new_n395_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT56), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT12), .B1(new_n515_), .B2(new_n517_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n518_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n510_), .B1(new_n773_), .B2(new_n503_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n512_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n503_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n777_), .A2(new_n775_), .A3(new_n513_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n771_), .B1(new_n780_), .B2(new_n526_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT56), .B(new_n525_), .C1(new_n776_), .C2(new_n779_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n783_), .A2(KEYINPUT114), .A3(new_n704_), .A4(new_n528_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n553_), .A2(new_n557_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n556_), .A2(new_n554_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n562_), .A3(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT115), .ZN(new_n788_));
  INV_X1    g587(.A(new_n559_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n563_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n529_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n775_), .B1(new_n777_), .B2(new_n513_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n512_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n526_), .B1(new_n794_), .B2(new_n778_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT56), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n771_), .B(new_n526_), .C1(new_n794_), .C2(new_n778_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n796_), .A2(new_n704_), .A3(new_n528_), .A4(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n784_), .A2(new_n791_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n622_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT116), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n801_), .A2(KEYINPUT57), .A3(new_n622_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n796_), .A2(new_n528_), .A3(new_n797_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n790_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(KEYINPUT58), .A3(new_n790_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n653_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n806_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT57), .B1(new_n801_), .B2(new_n622_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n805_), .A2(new_n813_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n585_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n586_), .A2(new_n534_), .A3(new_n565_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT113), .ZN(new_n820_));
  OR3_X1    g619(.A1(new_n820_), .A2(KEYINPUT54), .A3(new_n653_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT54), .B1(new_n820_), .B2(new_n653_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n770_), .B1(new_n818_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n704_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n818_), .A2(new_n823_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n769_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n806_), .A2(new_n812_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n585_), .B1(new_n828_), .B2(new_n814_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n823_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n770_), .A2(KEYINPUT59), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n827_), .A2(KEYINPUT59), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n704_), .A2(G113gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n825_), .B1(new_n832_), .B2(new_n833_), .ZN(G1340gat));
  NAND2_X1  g633(.A1(new_n830_), .A2(new_n831_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n535_), .B(new_n835_), .C1(new_n824_), .C2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G120gat), .ZN(new_n838_));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n534_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n824_), .B(new_n840_), .C1(KEYINPUT60), .C2(new_n839_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(G1341gat));
  AOI21_X1  g641(.A(G127gat), .B1(new_n824_), .B2(new_n586_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n586_), .A2(G127gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n832_), .B2(new_n844_), .ZN(G1342gat));
  AOI21_X1  g644(.A(G134gat), .B1(new_n824_), .B2(new_n623_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n653_), .A2(G134gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n832_), .B2(new_n847_), .ZN(G1343gat));
  NOR2_X1   g647(.A1(new_n406_), .A2(new_n429_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n826_), .A2(new_n704_), .A3(new_n678_), .A4(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g650(.A1(new_n826_), .A2(new_n535_), .A3(new_n678_), .A4(new_n849_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT117), .B(G148gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1345gat));
  NAND4_X1  g653(.A1(new_n826_), .A2(new_n586_), .A3(new_n678_), .A4(new_n849_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  AND3_X1   g656(.A1(new_n826_), .A2(new_n678_), .A3(new_n849_), .ZN(new_n858_));
  INV_X1    g657(.A(G162gat), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n618_), .A2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT118), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n826_), .A2(new_n623_), .A3(new_n678_), .A4(new_n849_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n858_), .A2(new_n861_), .B1(new_n862_), .B2(new_n859_), .ZN(G1347gat));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n676_), .A2(new_n429_), .A3(new_n704_), .A4(new_n677_), .ZN(new_n865_));
  OR3_X1    g664(.A1(new_n865_), .A2(KEYINPUT119), .A3(new_n441_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT119), .B1(new_n865_), .B2(new_n441_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n866_), .A2(new_n442_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n245_), .B1(new_n868_), .B2(new_n830_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n864_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n866_), .A2(new_n442_), .A3(new_n867_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n823_), .B2(new_n829_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT120), .B(KEYINPUT62), .C1(new_n873_), .C2(new_n245_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n869_), .A2(new_n870_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n871_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n678_), .A2(new_n428_), .A3(new_n395_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n830_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n704_), .A2(new_n224_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT121), .Z(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n881_), .ZN(G1348gat));
  NAND3_X1  g681(.A1(new_n878_), .A2(new_n225_), .A3(new_n535_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n826_), .A2(new_n535_), .A3(new_n877_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n225_), .ZN(G1349gat));
  NAND3_X1  g684(.A1(new_n826_), .A2(new_n586_), .A3(new_n877_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n586_), .A2(new_n243_), .A3(new_n237_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n886_), .A2(new_n239_), .B1(new_n878_), .B2(new_n887_), .ZN(G1350gat));
  NOR2_X1   g687(.A1(new_n622_), .A2(new_n235_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT122), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n878_), .A2(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n878_), .A2(new_n653_), .ZN(new_n892_));
  INV_X1    g691(.A(G190gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(G1351gat));
  INV_X1    g693(.A(new_n406_), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT123), .B1(new_n895_), .B2(new_n429_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n678_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n895_), .A2(KEYINPUT123), .A3(new_n429_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n815_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n901_));
  AOI211_X1 g700(.A(KEYINPUT116), .B(KEYINPUT57), .C1(new_n801_), .C2(new_n622_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n586_), .B1(new_n903_), .B2(new_n813_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n823_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n704_), .B(new_n900_), .C1(new_n904_), .C2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n210_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n906_), .B2(new_n210_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n906_), .A2(new_n210_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n908_), .A2(new_n909_), .A3(new_n910_), .ZN(G1352gat));
  AOI21_X1  g710(.A(new_n905_), .B1(new_n817_), .B2(new_n585_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n912_), .A2(new_n534_), .A3(new_n899_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n208_), .A2(KEYINPUT125), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n208_), .A2(KEYINPUT125), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n913_), .B2(new_n914_), .ZN(G1353gat));
  AOI21_X1  g716(.A(new_n585_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n900_), .B(new_n918_), .C1(new_n904_), .C2(new_n905_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT126), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n919_), .A2(new_n920_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n920_), .B1(new_n919_), .B2(new_n922_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n919_), .A2(new_n922_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(G1354gat));
  NOR2_X1   g725(.A1(new_n912_), .A2(new_n899_), .ZN(new_n927_));
  AOI21_X1  g726(.A(G218gat), .B1(new_n927_), .B2(new_n623_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n653_), .A2(G218gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(G1355gat));
endmodule


