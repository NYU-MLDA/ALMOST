//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  XNOR2_X1  g000(.A(KEYINPUT75), .B(G15gat), .ZN(new_n202_));
  INV_X1    g001(.A(G22gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT76), .B(G8gat), .Z(new_n205_));
  INV_X1    g004(.A(G1gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n204_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G29gat), .B(G36gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT78), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n219_), .A3(new_n216_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n213_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n216_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n221_), .A2(new_n222_), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n216_), .B(KEYINPUT15), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n218_), .A2(new_n220_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n228_), .B2(new_n222_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G113gat), .B(G141gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G169gat), .B(G197gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n230_), .B(new_n231_), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n232_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n226_), .B(new_n234_), .C1(new_n228_), .C2(new_n222_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT23), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT79), .B(G183gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n239_), .B1(G190gat), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT82), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n239_), .B(KEYINPUT82), .C1(G190gat), .C2(new_n240_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT81), .ZN(new_n245_));
  AOI21_X1  g044(.A(G176gat), .B1(new_n245_), .B2(KEYINPUT22), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G169gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G169gat), .ZN(new_n249_));
  INV_X1    g048(.A(G176gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT24), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(KEYINPUT24), .A3(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n239_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n240_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(G183gat), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n259_), .A2(KEYINPUT80), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(KEYINPUT80), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n256_), .B1(new_n258_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n248_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G71gat), .B(G99gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(G43gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n265_), .B(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G127gat), .B(G134gat), .Z(new_n269_));
  XOR2_X1   g068(.A(G113gat), .B(G120gat), .Z(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n268_), .B(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G227gat), .A2(G233gat), .ZN(new_n273_));
  INV_X1    g072(.A(G15gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT30), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT31), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n272_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT91), .ZN(new_n279_));
  XOR2_X1   g078(.A(G211gat), .B(G218gat), .Z(new_n280_));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n281_));
  INV_X1    g080(.A(G204gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(G197gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(G197gat), .ZN(new_n284_));
  INV_X1    g083(.A(G197gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n280_), .B1(new_n287_), .B2(KEYINPUT21), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(G204gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT21), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n284_), .A3(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n291_), .A2(KEYINPUT86), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(KEYINPUT86), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n288_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n280_), .A2(KEYINPUT87), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n290_), .B1(new_n289_), .B2(new_n284_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n294_), .A2(KEYINPUT88), .A3(new_n300_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n265_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT20), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n279_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n294_), .A2(KEYINPUT88), .A3(new_n300_), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT88), .B1(new_n294_), .B2(new_n300_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(KEYINPUT91), .B(KEYINPUT20), .C1(new_n313_), .C2(new_n265_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n239_), .B1(G183gat), .B2(G190gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT22), .B(G169gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n250_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n253_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n261_), .ZN(new_n319_));
  INV_X1    g118(.A(G183gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT25), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n259_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT92), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n259_), .A2(new_n321_), .A3(KEYINPUT92), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n319_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n318_), .B1(new_n255_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n301_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n307_), .A2(new_n310_), .A3(new_n314_), .A4(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT95), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n303_), .A2(new_n304_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n265_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n306_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n334_), .A2(KEYINPUT91), .B1(new_n301_), .B2(new_n327_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n335_), .A2(KEYINPUT95), .A3(new_n310_), .A4(new_n307_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT20), .B1(new_n327_), .B2(new_n301_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n313_), .B2(new_n265_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT94), .B1(new_n338_), .B2(new_n310_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT94), .ZN(new_n340_));
  INV_X1    g139(.A(new_n310_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n332_), .A2(new_n333_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n340_), .B(new_n341_), .C1(new_n342_), .C2(new_n337_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n331_), .A2(new_n336_), .A3(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT18), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n345_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT27), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n342_), .A2(new_n341_), .A3(new_n337_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n307_), .A2(new_n328_), .A3(new_n314_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(new_n341_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n352_), .B1(new_n355_), .B2(new_n349_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G155gat), .B(G162gat), .Z(new_n358_));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n361_), .A2(KEYINPUT83), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(KEYINPUT83), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n360_), .A2(new_n364_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n361_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT2), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n358_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n367_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT29), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n301_), .ZN(new_n378_));
  AND2_X1   g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n376_), .B2(KEYINPUT29), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n303_), .A2(new_n381_), .A3(new_n304_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n383_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT89), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n389_), .A2(new_n385_), .A3(new_n390_), .A4(new_n384_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n376_), .A2(KEYINPUT29), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n392_), .A2(KEYINPUT28), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(KEYINPUT28), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G22gat), .B(G50gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n393_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n396_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n388_), .A2(new_n391_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n376_), .A2(new_n271_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n269_), .B(new_n270_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(new_n367_), .A3(new_n375_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n402_), .A2(KEYINPUT4), .A3(new_n404_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n376_), .A2(new_n271_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n406_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G85gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT0), .B(G57gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  OR3_X1    g216(.A1(new_n408_), .A2(new_n412_), .A3(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n400_), .A2(new_n401_), .A3(new_n420_), .ZN(new_n421_));
  AOI211_X1 g220(.A(new_n350_), .B(new_n353_), .C1(new_n354_), .C2(new_n341_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n314_), .A2(new_n328_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n332_), .A2(new_n333_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT91), .B1(new_n424_), .B2(KEYINPUT20), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n341_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n353_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n349_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n352_), .B1(new_n422_), .B2(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n357_), .A2(new_n421_), .A3(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n400_), .A2(new_n401_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n418_), .A2(new_n419_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n433_), .B2(new_n355_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n345_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n422_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n428_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n419_), .A2(KEYINPUT93), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT93), .ZN(new_n442_));
  OAI221_X1 g241(.A(new_n417_), .B1(new_n442_), .B2(KEYINPUT33), .C1(new_n408_), .C2(new_n412_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n405_), .A2(new_n407_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n409_), .A2(new_n406_), .A3(new_n411_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n416_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n441_), .A2(new_n443_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n438_), .A2(new_n439_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n431_), .B1(new_n437_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n278_), .B1(new_n430_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n431_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n278_), .A2(new_n420_), .ZN(new_n453_));
  AND4_X1   g252(.A1(new_n452_), .A2(new_n357_), .A3(new_n453_), .A4(new_n429_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n237_), .B1(new_n451_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G230gat), .A2(G233gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G85gat), .ZN(new_n459_));
  INV_X1    g258(.A(G92gat), .ZN(new_n460_));
  OR3_X1    g259(.A1(new_n459_), .A2(new_n460_), .A3(KEYINPUT9), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n460_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G85gat), .A2(G92gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(KEYINPUT9), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT65), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT65), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT6), .ZN(new_n468_));
  AND2_X1   g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n466_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n469_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n461_), .B(new_n464_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n473_));
  NAND2_X1  g272(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n473_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT10), .ZN(new_n478_));
  INV_X1    g277(.A(G99gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(KEYINPUT64), .A3(new_n474_), .ZN(new_n481_));
  AOI21_X1  g280(.A(G106gat), .B1(new_n477_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT66), .B1(new_n472_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(G106gat), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n475_), .A2(new_n476_), .A3(new_n473_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT64), .B1(new_n480_), .B2(new_n474_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n484_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n461_), .A2(new_n464_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT66), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n467_), .A2(KEYINPUT6), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n465_), .A2(KEYINPUT65), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n466_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .A4(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n483_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n479_), .A2(new_n484_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT7), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n479_), .A2(new_n484_), .A3(KEYINPUT67), .A4(KEYINPUT7), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n493_), .A2(new_n494_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n462_), .A2(new_n463_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(KEYINPUT68), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT8), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n502_), .B1(G99gat), .B2(G106gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n504_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n507_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n497_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G57gat), .B(G64gat), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(KEYINPUT11), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(KEYINPUT11), .ZN(new_n520_));
  XOR2_X1   g319(.A(G71gat), .B(G78gat), .Z(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n520_), .A2(new_n521_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n517_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n497_), .A2(new_n516_), .A3(new_n524_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(KEYINPUT12), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n517_), .A2(new_n529_), .A3(new_n525_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n458_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n524_), .B1(new_n497_), .B2(new_n516_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT69), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n457_), .B1(new_n533_), .B2(new_n527_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n533_), .A2(new_n527_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n531_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G120gat), .B(G148gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT5), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G176gat), .B(G204gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT70), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n536_), .A2(new_n541_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT13), .ZN(new_n544_));
  OR4_X1    g343(.A1(KEYINPUT71), .A2(new_n542_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n544_), .A2(KEYINPUT71), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(KEYINPUT71), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n546_), .B(new_n547_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n550_));
  NAND2_X1  g349(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n517_), .A2(new_n227_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT73), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  OAI221_X1 g355(.A(new_n552_), .B1(KEYINPUT35), .B2(new_n556_), .C1(new_n224_), .C2(new_n517_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(KEYINPUT35), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n559_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n560_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n563_), .B(KEYINPUT36), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n560_), .B2(new_n565_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n550_), .B(new_n551_), .C1(new_n567_), .C2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n572_), .A2(KEYINPUT74), .A3(KEYINPUT37), .A4(new_n566_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n213_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n524_), .B(KEYINPUT77), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT16), .ZN(new_n580_));
  XOR2_X1   g379(.A(G183gat), .B(G211gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT17), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n578_), .B1(new_n585_), .B2(new_n582_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n549_), .A2(new_n574_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n456_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n420_), .A2(new_n206_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT97), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n590_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT98), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n567_), .A2(new_n570_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n451_), .B2(new_n455_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n587_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n549_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n597_), .A2(new_n236_), .A3(new_n598_), .A4(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G1gat), .B1(new_n600_), .B2(new_n432_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n593_), .A2(new_n595_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT99), .ZN(G1324gat));
  AND2_X1   g402(.A1(new_n357_), .A2(new_n429_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G8gat), .B1(new_n600_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT39), .ZN(new_n606_));
  INV_X1    g405(.A(new_n589_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n604_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n205_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g410(.A(G15gat), .B1(new_n600_), .B2(new_n278_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT100), .Z(new_n613_));
  OR2_X1    g412(.A1(new_n613_), .A2(KEYINPUT41), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(KEYINPUT41), .ZN(new_n615_));
  INV_X1    g414(.A(new_n278_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n607_), .A2(new_n274_), .A3(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n615_), .A3(new_n617_), .ZN(G1326gat));
  OAI21_X1  g417(.A(G22gat), .B1(new_n600_), .B2(new_n452_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT42), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n607_), .A2(new_n203_), .A3(new_n431_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1327gat));
  NAND2_X1  g421(.A1(new_n596_), .A2(new_n587_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n549_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n456_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(G29gat), .B1(new_n626_), .B2(new_n420_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n329_), .A2(new_n330_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n433_), .B1(new_n628_), .B2(new_n336_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n426_), .A2(new_n433_), .A3(new_n427_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n420_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n422_), .A2(new_n428_), .A3(new_n447_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n452_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n357_), .A2(new_n421_), .A3(new_n429_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n616_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n574_), .B1(new_n636_), .B2(new_n454_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT43), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n639_), .B(new_n574_), .C1(new_n636_), .C2(new_n454_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n599_), .A2(new_n236_), .A3(new_n587_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT44), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  AOI211_X1 g444(.A(new_n645_), .B(new_n642_), .C1(new_n638_), .C2(new_n640_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n420_), .A2(G29gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n627_), .B1(new_n647_), .B2(new_n648_), .ZN(G1328gat));
  INV_X1    g448(.A(new_n647_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G36gat), .B1(new_n650_), .B2(new_n604_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n625_), .A2(G36gat), .A3(new_n604_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT46), .ZN(G1329gat));
  NAND3_X1  g455(.A1(new_n647_), .A2(G43gat), .A3(new_n616_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n625_), .A2(new_n278_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(G43gat), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1330gat));
  OAI21_X1  g460(.A(G50gat), .B1(new_n650_), .B2(new_n452_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n452_), .A2(G50gat), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT103), .Z(new_n664_));
  OAI21_X1  g463(.A(new_n662_), .B1(new_n625_), .B2(new_n664_), .ZN(G1331gat));
  NAND2_X1  g464(.A1(new_n451_), .A2(new_n455_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n574_), .A2(new_n587_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n666_), .A2(new_n237_), .A3(new_n667_), .A4(new_n549_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G57gat), .B1(new_n669_), .B2(new_n420_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n549_), .A2(new_n237_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n587_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n597_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n432_), .A2(KEYINPUT104), .ZN(new_n675_));
  MUX2_X1   g474(.A(KEYINPUT104), .B(new_n675_), .S(G57gat), .Z(new_n676_));
  AOI21_X1  g475(.A(new_n670_), .B1(new_n674_), .B2(new_n676_), .ZN(G1332gat));
  OAI21_X1  g476(.A(G64gat), .B1(new_n673_), .B2(new_n604_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT48), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n604_), .A2(G64gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n668_), .B2(new_n680_), .ZN(G1333gat));
  OAI21_X1  g480(.A(G71gat), .B1(new_n673_), .B2(new_n278_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT49), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n278_), .A2(G71gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n668_), .B2(new_n684_), .ZN(G1334gat));
  OAI21_X1  g484(.A(G78gat), .B1(new_n673_), .B2(new_n452_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT50), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n452_), .A2(G78gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n668_), .B2(new_n688_), .ZN(G1335gat));
  AOI21_X1  g488(.A(new_n623_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n690_), .B(new_n237_), .C1(new_n636_), .C2(new_n454_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n459_), .A3(new_n420_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n549_), .A2(new_n237_), .A3(new_n587_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n639_), .B1(new_n666_), .B2(new_n574_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n640_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n695_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT105), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n641_), .A2(new_n700_), .A3(new_n695_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n432_), .B1(new_n699_), .B2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n693_), .B1(new_n702_), .B2(new_n459_), .ZN(G1336gat));
  NOR3_X1   g502(.A1(new_n691_), .A2(G92gat), .A3(new_n604_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n699_), .A2(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n608_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n706_), .B2(G92gat), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT106), .Z(G1337gat));
  AOI21_X1  g507(.A(new_n479_), .B1(new_n705_), .B2(new_n616_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n485_), .A2(new_n486_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n278_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n692_), .A2(KEYINPUT107), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713_));
  INV_X1    g512(.A(new_n711_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n691_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT51), .B1(new_n709_), .B2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n700_), .B1(new_n641_), .B2(new_n695_), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT105), .B(new_n694_), .C1(new_n638_), .C2(new_n640_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n616_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G99gat), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n716_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT109), .B1(new_n722_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727_));
  AOI211_X1 g526(.A(new_n727_), .B(new_n724_), .C1(new_n721_), .C2(G99gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n718_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT110), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n718_), .B(new_n731_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1338gat));
  NAND3_X1  g532(.A1(new_n692_), .A2(new_n484_), .A3(new_n431_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n641_), .A2(new_n431_), .A3(new_n695_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G106gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G106gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XOR2_X1   g538(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(G1339gat));
  NAND2_X1  g540(.A1(new_n527_), .A2(KEYINPUT12), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(new_n532_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n530_), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT55), .B(new_n457_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n528_), .A2(new_n458_), .A3(new_n530_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n531_), .A2(KEYINPUT55), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n540_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n457_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n540_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(new_n750_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n749_), .A2(new_n750_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n536_), .A2(new_n755_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n236_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT113), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n233_), .A2(new_n235_), .B1(new_n536_), .B2(new_n755_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n540_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n756_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n761_), .B(new_n762_), .C1(new_n763_), .C2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n228_), .A2(new_n222_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n221_), .A2(new_n225_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n767_), .B(new_n234_), .C1(new_n768_), .C2(new_n222_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n233_), .B(new_n769_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n760_), .A2(new_n766_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n596_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n771_), .A2(KEYINPUT57), .A3(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n749_), .A2(new_n750_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n764_), .A2(KEYINPUT114), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n754_), .A2(new_n779_), .A3(new_n756_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n778_), .A3(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n758_), .A2(new_n233_), .A3(new_n769_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(KEYINPUT58), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n781_), .A2(new_n782_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n781_), .A2(KEYINPUT115), .A3(KEYINPUT58), .A4(new_n782_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n785_), .A2(new_n788_), .A3(new_n574_), .A4(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n775_), .A2(new_n776_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT116), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n775_), .A2(new_n790_), .A3(new_n793_), .A4(new_n776_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n587_), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n599_), .A2(new_n237_), .A3(new_n667_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n588_), .A2(new_n237_), .A3(new_n797_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n795_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT117), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n795_), .A2(new_n805_), .A3(new_n802_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n608_), .A2(new_n431_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(new_n420_), .A3(new_n616_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n804_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(G113gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n236_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n808_), .A2(KEYINPUT59), .ZN(new_n814_));
  INV_X1    g613(.A(new_n776_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n775_), .A2(new_n790_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n775_), .A2(KEYINPUT118), .A3(new_n790_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n587_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n814_), .B1(new_n821_), .B2(new_n802_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n237_), .B(new_n822_), .C1(new_n810_), .C2(KEYINPUT59), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n813_), .B1(new_n823_), .B2(new_n812_), .ZN(G1340gat));
  AOI211_X1 g623(.A(new_n599_), .B(new_n822_), .C1(new_n810_), .C2(KEYINPUT59), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT119), .B(G120gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n599_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(KEYINPUT60), .B2(new_n826_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n825_), .A2(new_n826_), .B1(new_n810_), .B2(new_n828_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n811_), .A2(new_n830_), .A3(new_n598_), .ZN(new_n831_));
  AOI211_X1 g630(.A(new_n587_), .B(new_n822_), .C1(new_n810_), .C2(KEYINPUT59), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n830_), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n811_), .A2(new_n834_), .A3(new_n596_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n574_), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n836_), .B(new_n822_), .C1(new_n810_), .C2(KEYINPUT59), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n837_), .B2(new_n834_), .ZN(G1343gat));
  NAND2_X1  g637(.A1(new_n804_), .A2(new_n806_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n452_), .A2(new_n616_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n608_), .A2(new_n841_), .A3(new_n432_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n839_), .A2(new_n237_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(G141gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1344gat));
  NOR3_X1   g645(.A1(new_n839_), .A2(new_n599_), .A3(new_n843_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT120), .B(G148gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1345gat));
  NAND4_X1  g648(.A1(new_n804_), .A2(new_n598_), .A3(new_n806_), .A4(new_n842_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT121), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n598_), .B1(new_n791_), .B2(KEYINPUT116), .ZN(new_n852_));
  AOI211_X1 g651(.A(KEYINPUT117), .B(new_n801_), .C1(new_n852_), .C2(new_n794_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n805_), .B1(new_n795_), .B2(new_n802_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n598_), .A4(new_n842_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT61), .B(G155gat), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n851_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n851_), .B2(new_n857_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1346gat));
  NOR2_X1   g660(.A1(new_n839_), .A2(new_n843_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G162gat), .B1(new_n862_), .B2(new_n596_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n574_), .A2(G162gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT122), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n862_), .B2(new_n865_), .ZN(G1347gat));
  NAND2_X1  g665(.A1(new_n821_), .A2(new_n802_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n604_), .A2(new_n420_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n278_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n867_), .A2(new_n236_), .A3(new_n452_), .A4(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT123), .B1(new_n871_), .B2(G169gat), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n598_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n452_), .B(new_n870_), .C1(new_n874_), .C2(new_n801_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n237_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n872_), .A2(new_n873_), .B1(new_n316_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n876_), .B2(new_n249_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n871_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(KEYINPUT62), .A3(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n881_), .ZN(G1348gat));
  NOR2_X1   g681(.A1(new_n839_), .A2(new_n431_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n870_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n884_), .A2(new_n599_), .A3(new_n250_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n431_), .B1(new_n821_), .B2(new_n802_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n549_), .A3(new_n870_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n883_), .A2(new_n885_), .B1(new_n887_), .B2(new_n250_), .ZN(G1349gat));
  NOR2_X1   g687(.A1(new_n884_), .A2(new_n587_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n240_), .B1(new_n883_), .B2(new_n889_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n889_), .A2(new_n325_), .A3(new_n324_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n886_), .B2(new_n891_), .ZN(G1350gat));
  NAND4_X1  g691(.A1(new_n886_), .A2(new_n261_), .A3(new_n596_), .A4(new_n870_), .ZN(new_n893_));
  INV_X1    g692(.A(G190gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n875_), .A2(new_n836_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT124), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n893_), .B(new_n898_), .C1(new_n894_), .C2(new_n895_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1351gat));
  NOR2_X1   g699(.A1(new_n869_), .A2(new_n841_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n855_), .A2(new_n236_), .A3(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g702(.A(new_n599_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n855_), .A2(new_n901_), .A3(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n905_), .B(new_n906_), .Z(G1353gat));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n908_));
  INV_X1    g707(.A(G211gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(new_n909_), .A3(KEYINPUT126), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n598_), .B(new_n910_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n855_), .A2(new_n901_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(KEYINPUT126), .B1(new_n908_), .B2(new_n909_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1354gat));
  NAND4_X1  g714(.A1(new_n804_), .A2(new_n574_), .A3(new_n806_), .A4(new_n901_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G218gat), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n772_), .A2(G218gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n855_), .A2(new_n901_), .A3(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT127), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n917_), .A2(new_n922_), .A3(new_n919_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1355gat));
endmodule


