//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n865_, new_n866_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n208_));
  OR2_X1    g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n208_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT22), .B(G169gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(new_n214_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT75), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT76), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n207_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT24), .B1(new_n220_), .B2(new_n221_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n205_), .A2(new_n206_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT76), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n215_), .A2(new_n223_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT25), .B(G183gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT26), .B(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n230_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n218_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n240_), .B(KEYINPUT79), .Z(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT78), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n218_), .A2(new_n238_), .A3(new_n242_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G15gat), .B(G43gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT30), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G71gat), .B(G99gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(new_n248_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n251_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n202_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n255_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(KEYINPUT80), .A3(new_n253_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G127gat), .B(G134gat), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n259_), .A2(G113gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(G113gat), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n260_), .A2(G120gat), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(G120gat), .B1(new_n260_), .B2(new_n261_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT31), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n256_), .A2(new_n258_), .A3(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n267_), .B1(new_n258_), .B2(new_n266_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G1gat), .B(G29gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G57gat), .B(G85gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  INV_X1    g073(.A(KEYINPUT96), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT83), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n276_), .A2(KEYINPUT82), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(KEYINPUT82), .ZN(new_n278_));
  OAI22_X1  g077(.A1(new_n277_), .A2(new_n278_), .B1(G155gat), .B2(G162gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT2), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT81), .B1(G141gat), .B2(G148gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n285_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(KEYINPUT2), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT3), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT86), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT86), .ZN(new_n296_));
  OAI22_X1  g095(.A1(new_n296_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n283_), .B(new_n284_), .C1(new_n292_), .C2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT84), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT1), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT84), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n303_), .A3(new_n284_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n300_), .A2(KEYINPUT1), .A3(G155gat), .A4(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(new_n282_), .A3(new_n279_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT85), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n288_), .A2(new_n293_), .A3(new_n289_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n299_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n264_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n264_), .B(new_n299_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT94), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT94), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n317_), .A3(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G225gat), .A2(G233gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n275_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n320_), .ZN(new_n322_));
  AOI211_X1 g121(.A(KEYINPUT96), .B(new_n322_), .C1(new_n316_), .C2(new_n318_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n314_), .A2(KEYINPUT4), .ZN(new_n325_));
  AOI211_X1 g124(.A(new_n320_), .B(new_n325_), .C1(new_n319_), .C2(KEYINPUT4), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n274_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT99), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n319_), .A2(KEYINPUT4), .ZN(new_n329_));
  INV_X1    g128(.A(new_n325_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n322_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n274_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n331_), .B(new_n332_), .C1(new_n321_), .C2(new_n323_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n327_), .A2(new_n328_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n324_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n335_), .A2(KEYINPUT99), .A3(new_n331_), .A4(new_n332_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n269_), .A2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n339_));
  INV_X1    g138(.A(G197gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT87), .B1(new_n340_), .B2(G204gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT87), .ZN(new_n342_));
  INV_X1    g141(.A(G204gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(G197gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(G204gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT21), .ZN(new_n347_));
  XOR2_X1   g146(.A(G211gat), .B(G218gat), .Z(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT88), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(new_n340_), .B2(G204gat), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n343_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n352_));
  OAI22_X1  g151(.A1(new_n351_), .A2(new_n352_), .B1(new_n340_), .B2(G204gat), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n347_), .B(new_n349_), .C1(new_n353_), .C2(KEYINPUT21), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT21), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n348_), .B2(KEYINPUT89), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n356_), .B(new_n353_), .C1(KEYINPUT89), .C2(new_n348_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n312_), .A2(new_n339_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n354_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n311_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n298_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(G155gat), .B2(G162gat), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n362_), .A2(new_n363_), .B1(new_n365_), .B2(new_n283_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n361_), .B(new_n359_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n360_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G78gat), .ZN(new_n370_));
  INV_X1    g169(.A(G78gat), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n368_), .B(new_n371_), .C1(new_n359_), .C2(new_n358_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(G106gat), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G106gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n360_), .B2(new_n368_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n372_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n374_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n366_), .A2(new_n367_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G22gat), .B(G50gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT28), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n380_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(KEYINPUT91), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n373_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT91), .B1(new_n381_), .B2(new_n382_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  AOI211_X1 g186(.A(KEYINPUT91), .B(KEYINPUT92), .C1(new_n381_), .C2(new_n382_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n387_), .A2(new_n388_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n391_), .A2(new_n373_), .A3(new_n383_), .A4(new_n377_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n232_), .A2(new_n224_), .A3(new_n207_), .A4(new_n235_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n207_), .A2(new_n209_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n217_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n361_), .A2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT20), .B(new_n398_), .C1(new_n239_), .C2(new_n361_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT19), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n216_), .A2(new_n214_), .ZN(new_n403_));
  NOR4_X1   g202(.A1(new_n210_), .A2(new_n211_), .A3(new_n215_), .A4(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n236_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n361_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n401_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n357_), .A2(new_n354_), .A3(new_n394_), .A4(new_n396_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n406_), .A2(KEYINPUT20), .A3(new_n407_), .A4(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n402_), .A2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT18), .B(G64gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G92gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G8gat), .B(G36gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n414_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n410_), .A2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n402_), .A2(new_n415_), .A3(new_n416_), .A4(new_n409_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(KEYINPUT93), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT27), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT93), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n410_), .A2(new_n422_), .A3(new_n417_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  OR2_X1    g223(.A1(KEYINPUT97), .A2(KEYINPUT20), .ZN(new_n425_));
  NAND2_X1  g224(.A1(KEYINPUT97), .A2(KEYINPUT20), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n408_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n427_), .A2(KEYINPUT98), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT98), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n408_), .A2(new_n429_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n406_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n401_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n399_), .A2(new_n401_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n417_), .B(KEYINPUT100), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(KEYINPUT101), .A3(KEYINPUT27), .A4(new_n419_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT101), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n419_), .A2(KEYINPUT27), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n435_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n424_), .A2(new_n438_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n393_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n338_), .A2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n415_), .A2(KEYINPUT32), .A3(new_n416_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n410_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n434_), .A2(new_n447_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n334_), .A2(new_n336_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n335_), .A2(KEYINPUT33), .A3(new_n331_), .A4(new_n332_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n333_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n420_), .A2(new_n423_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n329_), .A2(new_n320_), .A3(new_n330_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n319_), .A2(new_n322_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n274_), .A3(new_n456_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n451_), .A2(new_n453_), .A3(new_n454_), .A4(new_n457_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n450_), .A2(new_n393_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n443_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n268_), .B1(new_n460_), .B2(new_n393_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT102), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n337_), .A2(new_n444_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n393_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n450_), .A2(new_n393_), .A3(new_n458_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT102), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .A4(new_n268_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n446_), .B1(new_n462_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT12), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT10), .B(G99gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT64), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n374_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n473_), .A2(KEYINPUT65), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n475_), .B(KEYINPUT6), .Z(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT66), .B(G92gat), .ZN(new_n478_));
  INV_X1    g277(.A(G85gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT67), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n476_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n473_), .A2(KEYINPUT65), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n474_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G85gat), .B(G92gat), .Z(new_n486_));
  NOR2_X1   g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT7), .Z(new_n488_));
  OAI21_X1  g287(.A(new_n486_), .B1(new_n488_), .B2(new_n476_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT8), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G57gat), .B(G64gat), .Z(new_n492_));
  INV_X1    g291(.A(KEYINPUT11), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G71gat), .A2(G78gat), .ZN(new_n495_));
  INV_X1    g294(.A(G71gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n371_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n492_), .A2(new_n493_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n470_), .B1(new_n491_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G230gat), .A2(G233gat), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n498_), .A2(KEYINPUT68), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(KEYINPUT68), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n505_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n501_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n485_), .B(new_n490_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n485_), .A2(new_n490_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n507_), .A2(new_n508_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT12), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n503_), .A2(new_n504_), .A3(new_n509_), .A4(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n509_), .B(KEYINPUT69), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n491_), .A2(new_n502_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n513_), .B1(new_n516_), .B2(new_n504_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G120gat), .B(G148gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(new_n343_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT5), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(new_n214_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n513_), .B(new_n521_), .C1(new_n516_), .C2(new_n504_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT13), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n523_), .B(new_n524_), .C1(KEYINPUT70), .C2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G29gat), .B(G36gat), .ZN(new_n531_));
  INV_X1    g330(.A(G43gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n533_), .A2(G50gat), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(G50gat), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537_));
  INV_X1    g336(.A(G1gat), .ZN(new_n538_));
  INV_X1    g337(.A(G8gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT14), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G1gat), .B(G8gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  OR2_X1    g342(.A1(new_n536_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n536_), .A2(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(KEYINPUT73), .A3(new_n545_), .ZN(new_n546_));
  OR3_X1    g345(.A1(new_n536_), .A2(KEYINPUT73), .A3(new_n543_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n546_), .A2(G229gat), .A3(G233gat), .A4(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n536_), .B(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n549_), .B(new_n545_), .C1(new_n551_), .C2(new_n543_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n548_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G169gat), .B(G197gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT74), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(G113gat), .ZN(new_n556_));
  INV_X1    g355(.A(G141gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n553_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n548_), .A2(new_n552_), .A3(new_n558_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n530_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n491_), .A2(new_n536_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT34), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n565_), .B(new_n568_), .C1(new_n551_), .C2(new_n491_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(G134gat), .ZN(new_n573_));
  INV_X1    g372(.A(G162gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT36), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n575_), .B(KEYINPUT36), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n578_), .B1(new_n579_), .B2(new_n571_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT37), .Z(new_n581_));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT71), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n543_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n511_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT16), .B(G183gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G211gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n589_), .A2(new_n590_), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n585_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n585_), .A2(new_n591_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  MUX2_X1   g394(.A(new_n593_), .B(new_n595_), .S(KEYINPUT72), .Z(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n581_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n469_), .A2(new_n564_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n337_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n538_), .A3(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT38), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n469_), .A2(new_n564_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n580_), .B(KEYINPUT103), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(new_n596_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n337_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n602_), .A2(new_n608_), .ZN(G1324gat));
  NAND3_X1  g408(.A1(new_n599_), .A2(new_n539_), .A3(new_n443_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611_));
  INV_X1    g410(.A(new_n607_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n443_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n613_), .B2(G8gat), .ZN(new_n614_));
  AOI211_X1 g413(.A(KEYINPUT39), .B(new_n539_), .C1(new_n612_), .C2(new_n443_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n610_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g416(.A(G15gat), .B1(new_n607_), .B2(new_n268_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT41), .Z(new_n619_));
  INV_X1    g418(.A(G15gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n599_), .A2(new_n620_), .A3(new_n269_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(G1326gat));
  OAI21_X1  g421(.A(G22gat), .B1(new_n607_), .B2(new_n393_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT42), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n623_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(G22gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n599_), .A2(new_n627_), .A3(new_n464_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1327gat));
  NOR2_X1   g428(.A1(new_n469_), .A2(new_n604_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n564_), .A2(new_n597_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(G29gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n600_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT106), .B1(new_n469_), .B2(new_n581_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT43), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT106), .B(new_n637_), .C1(new_n469_), .C2(new_n581_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT107), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n641_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n639_), .A2(new_n643_), .A3(new_n644_), .A4(new_n631_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n636_), .A2(new_n644_), .A3(new_n631_), .A4(new_n638_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n642_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n337_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n634_), .B1(new_n648_), .B2(new_n633_), .ZN(G1328gat));
  INV_X1    g448(.A(G36gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n632_), .A2(new_n650_), .A3(new_n443_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT45), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n444_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(new_n650_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT108), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(KEYINPUT46), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  OAI221_X1 g456(.A(new_n652_), .B1(new_n655_), .B2(KEYINPUT46), .C1(new_n653_), .C2(new_n650_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1329gat));
  AND2_X1   g458(.A1(new_n646_), .A2(new_n642_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n646_), .A2(new_n642_), .ZN(new_n661_));
  OAI211_X1 g460(.A(G43gat), .B(new_n269_), .C1(new_n660_), .C2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n632_), .A2(new_n269_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n532_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n662_), .A2(KEYINPUT47), .A3(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT47), .B1(new_n662_), .B2(new_n664_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1330gat));
  INV_X1    g466(.A(G50gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n632_), .A2(new_n668_), .A3(new_n464_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n464_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(G50gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n670_), .B2(G50gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(G1331gat));
  NOR2_X1   g473(.A1(new_n469_), .A2(new_n563_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n530_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n606_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n678_), .A2(G57gat), .A3(new_n600_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n598_), .A2(new_n530_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n675_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G57gat), .B1(new_n682_), .B2(new_n600_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n679_), .A2(new_n683_), .ZN(G1332gat));
  OR3_X1    g483(.A1(new_n681_), .A2(G64gat), .A3(new_n444_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G64gat), .B1(new_n677_), .B2(new_n444_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT110), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT110), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n687_), .A2(KEYINPUT48), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT48), .B1(new_n687_), .B2(new_n688_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n689_), .B2(new_n690_), .ZN(G1333gat));
  OAI21_X1  g490(.A(G71gat), .B1(new_n677_), .B2(new_n268_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT49), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n682_), .A2(new_n496_), .A3(new_n269_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1334gat));
  OAI21_X1  g494(.A(G78gat), .B1(new_n677_), .B2(new_n393_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT50), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n682_), .A2(new_n371_), .A3(new_n464_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1335gat));
  NAND3_X1  g498(.A1(new_n676_), .A2(new_n596_), .A3(new_n562_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n469_), .A2(new_n604_), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G85gat), .B1(new_n701_), .B2(new_n600_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n530_), .A2(new_n597_), .A3(new_n563_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT111), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n639_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(G85gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n702_), .B1(new_n706_), .B2(new_n600_), .ZN(G1336gat));
  AOI21_X1  g506(.A(G92gat), .B1(new_n701_), .B2(new_n443_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n444_), .A2(new_n478_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n705_), .B2(new_n709_), .ZN(G1337gat));
  NAND3_X1  g509(.A1(new_n701_), .A2(new_n472_), .A3(new_n269_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT112), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT113), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n636_), .A2(new_n704_), .A3(new_n269_), .A4(new_n638_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G99gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n712_), .A2(new_n713_), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n713_), .B1(new_n712_), .B2(new_n715_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n717_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n712_), .A2(new_n715_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT113), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT51), .B1(new_n722_), .B2(new_n716_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n720_), .A2(new_n723_), .ZN(G1338gat));
  NAND3_X1  g523(.A1(new_n701_), .A2(new_n374_), .A3(new_n464_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n636_), .A2(new_n704_), .A3(new_n464_), .A4(new_n638_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(G106gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n726_), .B2(G106gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g530(.A1(new_n581_), .A2(new_n597_), .A3(new_n562_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT54), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n733_), .A2(new_n530_), .A3(new_n736_), .A4(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n734_), .B(new_n735_), .C1(new_n732_), .C2(new_n676_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n546_), .A2(new_n549_), .A3(new_n547_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n545_), .B1(new_n551_), .B2(new_n543_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n741_), .B(new_n559_), .C1(new_n742_), .C2(new_n549_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT119), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n561_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(new_n561_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n525_), .A2(new_n747_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n503_), .A2(new_n504_), .A3(new_n512_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT117), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(KEYINPUT55), .A4(new_n509_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT117), .B1(new_n513_), .B2(new_n752_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n513_), .A2(new_n752_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n513_), .A2(KEYINPUT115), .A3(new_n752_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n504_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n503_), .A2(new_n512_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n514_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT116), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n760_), .C1(new_n514_), .C2(new_n761_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n754_), .A2(new_n759_), .A3(new_n763_), .A4(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n766_), .A2(KEYINPUT118), .A3(new_n767_), .A4(new_n522_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n513_), .A2(KEYINPUT115), .A3(new_n752_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT115), .B1(new_n513_), .B2(new_n752_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n753_), .B(new_n751_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n763_), .A2(new_n765_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n522_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n768_), .A2(new_n563_), .A3(new_n775_), .A4(new_n524_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(KEYINPUT56), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n748_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT120), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n779_), .A2(new_n604_), .A3(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n779_), .B2(new_n604_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n747_), .A2(new_n785_), .A3(new_n524_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n524_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n745_), .A2(new_n746_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT121), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT122), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n767_), .B(new_n522_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n790_), .A2(new_n777_), .A3(new_n792_), .A4(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n791_), .A2(KEYINPUT122), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n581_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n793_), .A2(new_n792_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n799_), .A2(new_n795_), .A3(new_n777_), .A4(new_n790_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n797_), .A2(new_n798_), .A3(new_n800_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n783_), .A2(new_n784_), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n740_), .B1(new_n802_), .B2(new_n597_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n445_), .A2(new_n337_), .A3(new_n268_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT123), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G113gat), .B1(new_n807_), .B2(new_n563_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(KEYINPUT59), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n562_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n808_), .B1(new_n812_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g612(.A(G120gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n530_), .B2(KEYINPUT60), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n807_), .B(new_n815_), .C1(KEYINPUT60), .C2(new_n814_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n530_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n814_), .ZN(G1341gat));
  AOI21_X1  g617(.A(G127gat), .B1(new_n807_), .B2(new_n597_), .ZN(new_n819_));
  INV_X1    g618(.A(G127gat), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n597_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n820_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n819_), .B1(new_n823_), .B2(new_n824_), .ZN(G1342gat));
  AOI21_X1  g624(.A(G134gat), .B1(new_n807_), .B2(new_n605_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n581_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g627(.A1(new_n269_), .A2(new_n393_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n784_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n801_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n779_), .A2(new_n604_), .A3(new_n782_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n596_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n830_), .B1(new_n835_), .B2(new_n740_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(new_n600_), .A3(new_n444_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n562_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(new_n557_), .ZN(G1344gat));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n530_), .ZN(new_n840_));
  INV_X1    g639(.A(G148gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1345gat));
  NOR2_X1   g641(.A1(new_n837_), .A2(new_n596_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT61), .B(G155gat), .Z(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1346gat));
  NOR3_X1   g644(.A1(new_n837_), .A2(new_n574_), .A3(new_n581_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n837_), .A2(new_n604_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n574_), .B2(new_n847_), .ZN(G1347gat));
  XNOR2_X1  g647(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n338_), .B1(new_n835_), .B2(new_n740_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n464_), .A2(new_n444_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n850_), .A2(new_n563_), .A3(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n849_), .B1(new_n852_), .B2(new_n213_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n851_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n563_), .A2(new_n216_), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT126), .Z(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G169gat), .B1(new_n854_), .B2(new_n562_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT62), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n853_), .B(new_n858_), .C1(new_n859_), .C2(new_n861_), .ZN(G1348gat));
  NOR2_X1   g661(.A1(new_n854_), .A2(new_n530_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(new_n214_), .ZN(G1349gat));
  NAND3_X1  g663(.A1(new_n855_), .A2(new_n597_), .A3(new_n233_), .ZN(new_n865_));
  OAI21_X1  g664(.A(G183gat), .B1(new_n854_), .B2(new_n596_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1350gat));
  NAND3_X1  g666(.A1(new_n855_), .A2(new_n605_), .A3(new_n234_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G190gat), .B1(new_n854_), .B2(new_n581_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1351gat));
  NOR2_X1   g669(.A1(new_n600_), .A2(new_n444_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT127), .B1(new_n836_), .B2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n803_), .A2(KEYINPUT127), .A3(new_n829_), .A4(new_n871_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n563_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G197gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n803_), .A2(new_n829_), .A3(new_n871_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT127), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n873_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(new_n340_), .A3(new_n563_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n881_), .ZN(G1352gat));
  AOI21_X1  g681(.A(G204gat), .B1(new_n880_), .B2(new_n676_), .ZN(new_n883_));
  AOI211_X1 g682(.A(new_n343_), .B(new_n530_), .C1(new_n879_), .C2(new_n873_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1353gat));
  XNOR2_X1  g684(.A(KEYINPUT63), .B(G211gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n880_), .A2(new_n597_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n596_), .B1(new_n879_), .B2(new_n873_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(G1354gat));
  AOI21_X1  g689(.A(G218gat), .B1(new_n880_), .B2(new_n605_), .ZN(new_n891_));
  INV_X1    g690(.A(G218gat), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n892_), .B(new_n581_), .C1(new_n879_), .C2(new_n873_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1355gat));
endmodule


