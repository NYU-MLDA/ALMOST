//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_;
  OR2_X1    g000(.A1(KEYINPUT70), .A2(G22gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(KEYINPUT70), .A2(G22gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G15gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n202_), .A2(G15gat), .A3(new_n203_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G1gat), .B(G8gat), .Z(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n206_), .A2(new_n212_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G50gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218_));
  INV_X1    g017(.A(G43gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G29gat), .A2(G36gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n219_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n217_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n223_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G50gat), .A3(new_n221_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n216_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT73), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n214_), .A2(new_n215_), .A3(new_n226_), .A4(new_n224_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n216_), .A2(KEYINPUT73), .A3(new_n227_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT15), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT15), .B1(new_n224_), .B2(new_n226_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n216_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n232_), .B(new_n230_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G113gat), .B(G141gat), .ZN(new_n243_));
  INV_X1    g042(.A(G169gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n242_), .A2(new_n247_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G99gat), .A2(G106gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT6), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT6), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(G99gat), .A3(G106gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NOR3_X1   g060(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n259_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n253_), .A2(new_n255_), .A3(KEYINPUT65), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT7), .ZN(new_n265_));
  INV_X1    g064(.A(G99gat), .ZN(new_n266_));
  INV_X1    g065(.A(G106gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT66), .A3(new_n260_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n258_), .A2(new_n263_), .A3(new_n264_), .A4(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT8), .ZN(new_n271_));
  INV_X1    g070(.A(G85gat), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n272_), .A2(G92gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(G92gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n271_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G57gat), .ZN(new_n277_));
  INV_X1    g076(.A(G64gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G57gat), .A2(G64gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT11), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G71gat), .B(G78gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT11), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n279_), .A2(new_n285_), .A3(new_n280_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n281_), .A2(new_n283_), .A3(KEYINPUT11), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n273_), .A2(new_n274_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n253_), .A2(new_n255_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n268_), .A2(new_n260_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n271_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(KEYINPUT9), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT10), .B(G99gat), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n267_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n272_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(G85gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(G92gat), .B1(new_n298_), .B2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n295_), .A2(new_n297_), .A3(new_n256_), .A4(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n276_), .A2(new_n289_), .A3(new_n294_), .A4(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G230gat), .A2(G233gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT67), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n276_), .A2(new_n294_), .A3(new_n302_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n289_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT12), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n307_), .A2(KEYINPUT12), .A3(new_n308_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n303_), .A2(new_n313_), .A3(new_n304_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n306_), .A2(new_n311_), .A3(new_n312_), .A4(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n303_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G230gat), .A3(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318_));
  INV_X1    g117(.A(G204gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT5), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n315_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n315_), .A2(new_n317_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n323_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n315_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT68), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT13), .B1(new_n327_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n307_), .A2(new_n227_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G232gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT34), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT35), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n307_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n337_), .A2(KEYINPUT35), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n335_), .A2(new_n338_), .A3(new_n339_), .A4(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n294_), .A2(new_n302_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT15), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n227_), .A2(new_n343_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n342_), .A2(new_n276_), .B1(new_n344_), .B2(new_n236_), .ZN(new_n345_));
  OAI211_X1 g144(.A(KEYINPUT35), .B(new_n337_), .C1(new_n345_), .C2(new_n334_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G190gat), .B(G218gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(G134gat), .ZN(new_n349_));
  INV_X1    g148(.A(G162gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT36), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT37), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n349_), .B(G162gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT36), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n347_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(new_n355_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT69), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n353_), .A2(new_n357_), .A3(new_n360_), .ZN(new_n362_));
  AOI211_X1 g161(.A(new_n361_), .B(new_n362_), .C1(new_n341_), .C2(new_n346_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n347_), .A2(new_n353_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT37), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n359_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n216_), .B(new_n308_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G231gat), .A2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G127gat), .B(G155gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G183gat), .B(G211gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT17), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n374_), .A2(KEYINPUT17), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n369_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n376_), .B2(new_n369_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n326_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n330_), .A2(KEYINPUT68), .A3(new_n331_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT13), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n333_), .A2(new_n366_), .A3(new_n379_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT72), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n251_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G1gat), .B(G29gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G57gat), .B(G85gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n389_), .B(new_n390_), .Z(new_n391_));
  NOR2_X1   g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G155gat), .A2(G162gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(KEYINPUT81), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(KEYINPUT3), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n398_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT2), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n397_), .B1(KEYINPUT81), .B2(new_n399_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n403_), .A2(new_n405_), .A3(KEYINPUT82), .A4(new_n406_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n396_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n404_), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n395_), .B(KEYINPUT1), .Z(new_n413_));
  AOI211_X1 g212(.A(new_n397_), .B(new_n412_), .C1(new_n413_), .C2(new_n394_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G127gat), .B(G134gat), .ZN(new_n416_));
  INV_X1    g215(.A(G113gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G120gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n421_), .A2(KEYINPUT4), .A3(new_n422_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n422_), .A2(KEYINPUT4), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n391_), .B(new_n425_), .C1(new_n428_), .C2(new_n424_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT96), .ZN(new_n430_));
  INV_X1    g229(.A(new_n391_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n423_), .A2(new_n424_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n429_), .A2(new_n430_), .A3(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n432_), .A2(new_n433_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT96), .A3(new_n391_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT98), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(KEYINPUT98), .A3(new_n437_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT21), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n246_), .A2(G204gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT84), .B(G197gat), .Z(new_n446_));
  OAI211_X1 g245(.A(new_n443_), .B(new_n445_), .C1(new_n446_), .C2(new_n319_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G211gat), .B(G218gat), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(KEYINPUT85), .A3(new_n319_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n246_), .A2(G204gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT85), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT84), .B(G197gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(G204gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n450_), .B1(KEYINPUT21), .B2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n444_), .B1(new_n454_), .B2(G204gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n448_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT21), .B1(new_n458_), .B2(new_n459_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT87), .B1(new_n457_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT29), .B1(new_n411_), .B2(new_n414_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n456_), .A2(KEYINPUT21), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n448_), .B1(new_n458_), .B2(new_n443_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n449_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n470_), .B(KEYINPUT21), .C1(new_n459_), .C2(new_n458_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n464_), .A2(new_n465_), .A3(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(G228gat), .A3(G233gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n457_), .A2(new_n463_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G228gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT83), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n465_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G78gat), .B(G106gat), .Z(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n411_), .A2(new_n414_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n484_), .A2(KEYINPUT29), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G22gat), .B(G50gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT28), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n485_), .B(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n481_), .B(KEYINPUT88), .Z(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n474_), .A2(new_n490_), .A3(new_n479_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n483_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n480_), .A2(new_n489_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n491_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n487_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n485_), .B(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT89), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n474_), .A2(new_n490_), .A3(new_n479_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n490_), .B1(new_n474_), .B2(new_n479_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT89), .B(new_n497_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n493_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G15gat), .B(G43gat), .Z(new_n504_));
  XOR2_X1   g303(.A(new_n419_), .B(new_n504_), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G183gat), .ZN(new_n507_));
  INV_X1    g306(.A(G190gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT23), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT78), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT23), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(G183gat), .A3(G190gat), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n509_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n508_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G169gat), .A2(G176gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT22), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT77), .B1(new_n519_), .B2(G169gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT22), .B(G169gat), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n322_), .B(new_n520_), .C1(new_n521_), .C2(KEYINPUT77), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(new_n518_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n244_), .A2(new_n322_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT24), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT25), .B(G183gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G190gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT74), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n525_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(KEYINPUT24), .A3(new_n518_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT75), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT76), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n512_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(new_n509_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n528_), .A2(KEYINPUT74), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n531_), .A2(new_n534_), .A3(new_n537_), .A4(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n523_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n540_), .B1(new_n523_), .B2(new_n539_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT31), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n523_), .A2(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT30), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT31), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n523_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G227gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT79), .ZN(new_n550_));
  XOR2_X1   g349(.A(G71gat), .B(G99gat), .Z(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n543_), .A2(new_n548_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n553_), .B1(new_n543_), .B2(new_n548_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n506_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n543_), .A2(new_n548_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n552_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n543_), .A2(new_n548_), .A3(new_n553_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n505_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n503_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n497_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n501_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n561_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n493_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n442_), .B1(new_n562_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT20), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n476_), .B2(new_n544_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n525_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n515_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n537_), .A2(new_n516_), .B1(G169gat), .B2(G176gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n521_), .B(KEYINPUT90), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n322_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n572_), .A2(new_n573_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n475_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G226gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT19), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n577_), .A2(new_n475_), .A3(KEYINPUT92), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n571_), .A2(new_n580_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n468_), .A2(new_n523_), .A3(new_n539_), .A4(new_n471_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n586_), .B(KEYINPUT20), .C1(new_n577_), .C2(new_n475_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n587_), .A2(KEYINPUT91), .A3(new_n582_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT91), .B1(new_n587_), .B2(new_n582_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n585_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT18), .B(G64gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(G92gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G8gat), .B(G36gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n594_), .B(new_n585_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT27), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n464_), .A2(new_n472_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n577_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n583_), .B1(new_n600_), .B2(new_n571_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n587_), .A2(new_n582_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n595_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n597_), .A2(KEYINPUT27), .A3(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n598_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n594_), .A2(KEYINPUT32), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n606_), .B(new_n585_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n607_));
  OAI211_X1 g406(.A(KEYINPUT32), .B(new_n594_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT97), .B1(new_n438_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n437_), .A4(new_n435_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n587_), .A2(new_n582_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n587_), .A2(KEYINPUT91), .A3(new_n582_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n594_), .B1(new_n618_), .B2(new_n585_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n597_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT93), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT93), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n596_), .A2(new_n622_), .A3(new_n597_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n434_), .A2(KEYINPUT95), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT33), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n431_), .B1(new_n428_), .B2(new_n424_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n424_), .B2(new_n423_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n434_), .A2(KEYINPUT95), .A3(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n610_), .B(new_n613_), .C1(new_n624_), .C2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n503_), .A2(new_n567_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n569_), .A2(new_n605_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n386_), .B(new_n634_), .C1(new_n385_), .C2(new_n384_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n207_), .A3(new_n442_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT100), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n354_), .A2(new_n358_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n382_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n251_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n379_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n634_), .A2(new_n641_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n207_), .B1(new_n649_), .B2(new_n442_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n639_), .A2(new_n651_), .ZN(G1324gat));
  INV_X1    g451(.A(new_n605_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n635_), .A2(new_n208_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n649_), .A2(new_n653_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(G8gat), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT39), .B(new_n208_), .C1(new_n649_), .C2(new_n653_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT101), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n661_), .B(new_n654_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(KEYINPUT40), .A3(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1325gat));
  AOI21_X1  g466(.A(new_n205_), .B1(new_n649_), .B2(new_n567_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT41), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n635_), .A2(new_n205_), .A3(new_n567_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT102), .Z(G1326gat));
  NAND2_X1  g471(.A1(new_n649_), .A2(new_n503_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G22gat), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT103), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n676_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n635_), .A2(new_n503_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n677_), .B(new_n678_), .C1(G22gat), .C2(new_n679_), .ZN(G1327gat));
  INV_X1    g479(.A(new_n379_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n647_), .A2(new_n681_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n634_), .A2(new_n640_), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G29gat), .B1(new_n683_), .B2(new_n442_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n682_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n632_), .A2(new_n633_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n441_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT98), .B1(new_n435_), .B2(new_n437_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n567_), .B1(new_n566_), .B2(new_n493_), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n561_), .B(new_n492_), .C1(new_n565_), .C2(new_n501_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n690_), .B(new_n605_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n687_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n366_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n686_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT43), .B(new_n366_), .C1(new_n687_), .C2(new_n693_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT44), .B(new_n685_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n634_), .B2(new_n366_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n694_), .A2(new_n686_), .A3(new_n695_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n682_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT104), .B1(new_n702_), .B2(KEYINPUT44), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n685_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n704_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n699_), .B1(new_n703_), .B2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n442_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n684_), .B1(new_n709_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n708_), .B2(new_n653_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n683_), .A2(new_n712_), .A3(new_n653_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n714_), .B(new_n715_), .Z(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n711_), .B1(new_n713_), .B2(new_n717_), .ZN(new_n718_));
  AOI211_X1 g517(.A(new_n605_), .B(new_n699_), .C1(new_n703_), .C2(new_n707_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT46), .B(new_n716_), .C1(new_n719_), .C2(new_n712_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1329gat));
  XNOR2_X1  g520(.A(KEYINPUT106), .B(G43gat), .ZN(new_n722_));
  INV_X1    g521(.A(new_n683_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n561_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n702_), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n705_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n726_));
  OAI211_X1 g525(.A(G43gat), .B(new_n698_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n727_), .B2(new_n561_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT47), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n730_), .B(new_n724_), .C1(new_n727_), .C2(new_n561_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1330gat));
  AOI21_X1  g531(.A(G50gat), .B1(new_n683_), .B2(new_n503_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n503_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n734_), .A2(new_n217_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n708_), .B2(new_n735_), .ZN(G1331gat));
  NOR2_X1   g535(.A1(new_n634_), .A2(new_n251_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n644_), .A2(new_n681_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n640_), .A3(new_n738_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n739_), .A2(new_n277_), .A3(new_n690_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(new_n366_), .A3(new_n738_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n442_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n740_), .B1(new_n277_), .B2(new_n743_), .ZN(G1332gat));
  OAI21_X1  g543(.A(G64gat), .B1(new_n739_), .B2(new_n605_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT48), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(new_n278_), .A3(new_n653_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1333gat));
  OR3_X1    g547(.A1(new_n741_), .A2(G71gat), .A3(new_n561_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n739_), .A2(new_n561_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G71gat), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT107), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n753_), .A3(G71gat), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n752_), .A2(KEYINPUT49), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT49), .B1(new_n752_), .B2(new_n754_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n749_), .B1(new_n755_), .B2(new_n756_), .ZN(G1334gat));
  OAI21_X1  g556(.A(G78gat), .B1(new_n739_), .B2(new_n734_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT50), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n734_), .A2(G78gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n741_), .B2(new_n760_), .ZN(G1335gat));
  NAND3_X1  g560(.A1(new_n645_), .A2(new_n681_), .A3(new_n646_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n634_), .A2(new_n640_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G85gat), .B1(new_n763_), .B2(new_n442_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n762_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n700_), .A2(KEYINPUT108), .A3(new_n701_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n300_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n299_), .A2(G85gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n690_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n764_), .B1(new_n769_), .B2(new_n772_), .ZN(G1336gat));
  AOI21_X1  g572(.A(G92gat), .B1(new_n763_), .B2(new_n653_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n769_), .A2(new_n653_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(G92gat), .ZN(G1337gat));
  NAND4_X1  g575(.A1(new_n766_), .A2(new_n768_), .A3(new_n567_), .A4(new_n767_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(G99gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n763_), .A2(new_n296_), .A3(new_n567_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g580(.A1(new_n762_), .A2(new_n734_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n784_), .B2(new_n267_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n782_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(G106gat), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n763_), .A2(new_n267_), .A3(new_n503_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT109), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(KEYINPUT53), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n793_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n790_), .ZN(new_n798_));
  AOI211_X1 g597(.A(KEYINPUT109), .B(new_n798_), .C1(new_n785_), .C2(new_n788_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n796_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n795_), .A2(new_n800_), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n690_), .A2(new_n653_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n324_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n315_), .A2(new_n804_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n307_), .A2(KEYINPUT12), .A3(new_n308_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT12), .B1(new_n307_), .B2(new_n308_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n808_), .A2(KEYINPUT55), .A3(new_n306_), .A4(new_n314_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n311_), .A2(new_n303_), .A3(new_n312_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(G230gat), .A3(G233gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n805_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n329_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n329_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n803_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n231_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n247_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n816_), .B2(new_n247_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n233_), .B(new_n230_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n248_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n641_), .B1(new_n815_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT57), .B1(new_n824_), .B2(KEYINPUT113), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n251_), .A2(new_n331_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n812_), .A2(new_n329_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n329_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n826_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n822_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n640_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n825_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n829_), .A2(KEYINPUT116), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n830_), .A2(KEYINPUT115), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n812_), .A2(new_n840_), .A3(KEYINPUT56), .A4(new_n329_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n814_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n838_), .A2(new_n839_), .A3(new_n841_), .A4(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n822_), .A2(new_n331_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n822_), .A2(KEYINPUT114), .A3(new_n331_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n844_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n844_), .A2(new_n849_), .A3(KEYINPUT58), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n695_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n379_), .B1(new_n837_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n644_), .A2(new_n379_), .A3(new_n366_), .A4(new_n646_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(KEYINPUT54), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT54), .B1(new_n384_), .B2(new_n251_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT111), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n384_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n862_), .A2(KEYINPUT110), .A3(new_n863_), .A4(new_n646_), .ZN(new_n864_));
  OAI211_X1 g663(.A(KEYINPUT111), .B(KEYINPUT54), .C1(new_n384_), .C2(new_n251_), .ZN(new_n865_));
  AND4_X1   g664(.A1(new_n858_), .A2(new_n861_), .A3(new_n864_), .A4(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n692_), .B(new_n802_), .C1(new_n855_), .C2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G113gat), .B1(new_n868_), .B2(new_n251_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n844_), .A2(KEYINPUT58), .A3(new_n849_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT58), .B1(new_n844_), .B2(new_n849_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n366_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n825_), .A2(new_n836_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n681_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n858_), .A2(new_n861_), .A3(new_n864_), .A4(new_n865_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n568_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(KEYINPUT59), .B1(new_n877_), .B2(new_n802_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n867_), .A2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n870_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n877_), .A2(KEYINPUT59), .A3(new_n802_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n867_), .A2(new_n879_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(new_n883_), .A3(KEYINPUT117), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n646_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n869_), .B1(new_n885_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g685(.A(G120gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n644_), .B2(KEYINPUT60), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n868_), .B(new_n888_), .C1(KEYINPUT60), .C2(new_n887_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n644_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n887_), .ZN(G1341gat));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT119), .B(G127gat), .Z(new_n893_));
  NOR2_X1   g692(.A1(new_n681_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n896_));
  INV_X1    g695(.A(G127gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n867_), .B2(new_n681_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT118), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n892_), .B1(new_n896_), .B2(new_n899_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n882_), .A2(new_n883_), .A3(KEYINPUT117), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT117), .B1(new_n882_), .B2(new_n883_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n894_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n898_), .B(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(KEYINPUT120), .A3(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n900_), .A2(new_n906_), .ZN(G1342gat));
  AOI21_X1  g706(.A(G134gat), .B1(new_n868_), .B2(new_n641_), .ZN(new_n908_));
  INV_X1    g707(.A(G134gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n910_), .B2(new_n695_), .ZN(G1343gat));
  AOI21_X1  g710(.A(new_n562_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n802_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n646_), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n644_), .ZN(new_n916_));
  XOR2_X1   g715(.A(new_n916_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g716(.A1(new_n913_), .A2(new_n681_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT61), .B(G155gat), .Z(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1346gat));
  NOR3_X1   g719(.A1(new_n913_), .A2(new_n350_), .A3(new_n366_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n913_), .A2(new_n640_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(G162gat), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n923_), .A2(KEYINPUT121), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(KEYINPUT121), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n921_), .B1(new_n924_), .B2(new_n925_), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n442_), .A2(new_n605_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n877_), .A2(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928_), .B2(new_n646_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n929_), .A2(KEYINPUT122), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(KEYINPUT122), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n930_), .A2(KEYINPUT62), .A3(new_n931_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n877_), .A2(new_n251_), .A3(new_n575_), .A4(new_n927_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT62), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n929_), .A2(KEYINPUT122), .A3(new_n934_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n932_), .A2(new_n933_), .A3(new_n935_), .ZN(G1348gat));
  AOI211_X1 g735(.A(new_n644_), .B(new_n928_), .C1(KEYINPUT123), .C2(new_n322_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n322_), .A2(KEYINPUT123), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(KEYINPUT124), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n937_), .B(new_n939_), .ZN(G1349gat));
  NOR2_X1   g739(.A1(new_n928_), .A2(new_n681_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n526_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n942_), .B1(new_n507_), .B2(new_n941_), .ZN(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n928_), .B2(new_n366_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n641_), .A2(new_n527_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n928_), .B2(new_n945_), .ZN(G1351gat));
  OAI211_X1 g745(.A(new_n691_), .B(new_n927_), .C1(new_n855_), .C2(new_n866_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n646_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n246_), .ZN(G1352gat));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n950_), .B1(new_n947_), .B2(new_n644_), .ZN(new_n951_));
  NAND4_X1  g750(.A1(new_n912_), .A2(KEYINPUT125), .A3(new_n645_), .A4(new_n927_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n951_), .A2(new_n952_), .A3(G204gat), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n947_), .A2(new_n644_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n954_), .B1(new_n955_), .B2(new_n319_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n953_), .A2(new_n956_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n951_), .A2(new_n952_), .A3(new_n954_), .A4(G204gat), .ZN(new_n959_));
  AND3_X1   g758(.A1(new_n957_), .A2(new_n958_), .A3(new_n959_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n958_), .B1(new_n957_), .B2(new_n959_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1353gat));
  INV_X1    g761(.A(new_n947_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n963_), .A2(new_n379_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  AND2_X1   g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n964_), .A2(new_n965_), .A3(new_n966_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n967_), .B1(new_n964_), .B2(new_n965_), .ZN(G1354gat));
  INV_X1    g767(.A(G218gat), .ZN(new_n969_));
  NOR3_X1   g768(.A1(new_n947_), .A2(new_n969_), .A3(new_n366_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n963_), .A2(new_n641_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n970_), .B1(new_n971_), .B2(new_n969_), .ZN(G1355gat));
endmodule


