//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G127gat), .A2(G134gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G127gat), .A2(G134gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(G113gat), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G127gat), .ZN(new_n207_));
  INV_X1    g006(.A(G134gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G113gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(new_n203_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(G120gat), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(G120gat), .B1(new_n206_), .B2(new_n211_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n202_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n214_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(KEYINPUT87), .A3(new_n212_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT31), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT78), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n225_), .A2(KEYINPUT79), .A3(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT79), .B1(new_n225_), .B2(new_n226_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n221_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT77), .B1(new_n232_), .B2(G183gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT26), .B(G190gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT25), .B(G183gat), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n233_), .B(new_n234_), .C1(new_n235_), .C2(KEYINPUT77), .ZN(new_n236_));
  OAI211_X1 g035(.A(KEYINPUT80), .B(new_n221_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n231_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT81), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT81), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n231_), .A2(new_n240_), .A3(new_n236_), .A4(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n225_), .A2(new_n226_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT79), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n225_), .A2(KEYINPUT79), .A3(new_n226_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n220_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT82), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G183gat), .A2(G190gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT23), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n246_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n247_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n239_), .A2(new_n241_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT30), .ZN(new_n254_));
  OR2_X1    g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n249_), .A2(new_n255_), .B1(G169gat), .B2(G176gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n223_), .A2(KEYINPUT22), .ZN(new_n257_));
  AOI21_X1  g056(.A(G176gat), .B1(new_n257_), .B2(KEYINPUT83), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT83), .B1(KEYINPUT84), .B2(G169gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT22), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT84), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n223_), .A2(KEYINPUT22), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n258_), .B(new_n260_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n256_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n253_), .A2(new_n254_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n254_), .B1(new_n253_), .B2(new_n264_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT86), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT86), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n265_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G71gat), .B(G99gat), .Z(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT85), .B(G15gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G43gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n274_), .B(new_n276_), .Z(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n268_), .A2(new_n271_), .A3(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(KEYINPUT86), .B(new_n277_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n219_), .B1(new_n281_), .B2(KEYINPUT88), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(KEYINPUT88), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT88), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(new_n280_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n282_), .B1(new_n286_), .B2(new_n219_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G78gat), .B(G106gat), .Z(new_n288_));
  XNOR2_X1  g087(.A(G197gat), .B(G204gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT21), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT91), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G197gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(G204gat), .ZN(new_n297_));
  INV_X1    g096(.A(G204gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(G197gat), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n292_), .B(KEYINPUT21), .C1(new_n297_), .C2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n289_), .A2(new_n290_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(new_n293_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT92), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G228gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT29), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT3), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT89), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n309_), .B(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n308_), .B(new_n312_), .C1(new_n314_), .C2(KEYINPUT2), .ZN(new_n315_));
  INV_X1    g114(.A(G155gat), .ZN(new_n316_));
  INV_X1    g115(.A(G162gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n316_), .A2(new_n317_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n315_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT1), .B1(new_n316_), .B2(new_n317_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n309_), .B(KEYINPUT89), .ZN(new_n326_));
  INV_X1    g125(.A(new_n307_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n321_), .A2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n304_), .B(new_n305_), .C1(new_n306_), .C2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n306_), .B1(new_n321_), .B2(new_n328_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n295_), .A2(new_n302_), .ZN(new_n332_));
  OAI211_X1 g131(.A(G228gat), .B(G233gat), .C1(new_n331_), .C2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n288_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n321_), .A2(new_n328_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G22gat), .B(G50gat), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n335_), .A2(KEYINPUT29), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n335_), .B2(KEYINPUT29), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n340_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n336_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n343_), .B1(new_n329_), .B2(new_n306_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n342_), .B1(new_n344_), .B2(new_n337_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT93), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n330_), .A2(new_n333_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n288_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n330_), .A2(KEYINPUT93), .A3(new_n288_), .A4(new_n333_), .ZN(new_n351_));
  AOI211_X1 g150(.A(new_n334_), .B(new_n346_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n348_), .B1(new_n353_), .B2(new_n288_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n330_), .A2(KEYINPUT94), .A3(new_n349_), .A4(new_n333_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n346_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n253_), .A2(new_n264_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n304_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n235_), .A2(new_n234_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n242_), .A2(new_n220_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n229_), .A2(new_n249_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n262_), .A2(new_n257_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n256_), .B1(G176gat), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n332_), .A3(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n366_), .A2(KEYINPUT20), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT19), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n304_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n253_), .A2(new_n264_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n375_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n369_), .A2(new_n371_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(new_n303_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(new_n379_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n364_), .B1(new_n376_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n378_), .A2(new_n382_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n375_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n372_), .A2(KEYINPUT95), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT95), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n369_), .A2(new_n332_), .A3(new_n371_), .A4(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n387_), .A2(KEYINPUT20), .A3(new_n379_), .A4(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n366_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n386_), .A2(new_n364_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT27), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT99), .B1(new_n384_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT27), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n379_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n390_), .B1(new_n365_), .B2(new_n304_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(new_n364_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n397_), .A2(new_n398_), .A3(new_n363_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n396_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n372_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n365_), .B2(new_n304_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n379_), .B1(new_n404_), .B2(KEYINPUT20), .ZN(new_n405_));
  INV_X1    g204(.A(new_n383_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n363_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n396_), .B1(new_n399_), .B2(new_n364_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT99), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n358_), .A2(new_n395_), .A3(new_n402_), .A4(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G85gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT0), .ZN(new_n414_));
  INV_X1    g213(.A(G57gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G225gat), .A2(G233gat), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n217_), .A2(new_n215_), .B1(new_n321_), .B2(new_n328_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n213_), .A2(new_n214_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n321_), .A2(new_n420_), .A3(new_n328_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT4), .B1(new_n419_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT4), .B1(new_n218_), .B2(new_n335_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n418_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n218_), .A2(new_n335_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n418_), .A3(new_n421_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n417_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n421_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n424_), .B1(new_n431_), .B2(KEYINPUT4), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n428_), .B(new_n416_), .C1(new_n432_), .C2(new_n418_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n287_), .A2(new_n411_), .A3(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n409_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n352_), .A2(new_n434_), .A3(new_n357_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n438_), .A2(KEYINPUT100), .A3(new_n439_), .A4(new_n402_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n400_), .A2(new_n401_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n418_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n427_), .A2(new_n442_), .A3(new_n421_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n417_), .B(new_n443_), .C1(new_n432_), .C2(new_n442_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT97), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n433_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n445_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n423_), .A2(new_n425_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n442_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n451_), .A2(KEYINPUT33), .A3(new_n428_), .A4(new_n416_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n448_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n441_), .A2(new_n446_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n399_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n434_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n455_), .B1(new_n376_), .B2(new_n383_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT98), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(KEYINPUT32), .B(new_n364_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT98), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n434_), .A4(new_n456_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n454_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n358_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n395_), .A2(new_n439_), .A3(new_n402_), .A4(new_n410_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT100), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n440_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n435_), .B1(new_n468_), .B2(new_n287_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT73), .ZN(new_n471_));
  INV_X1    g270(.A(G15gat), .ZN(new_n472_));
  INV_X1    g271(.A(G22gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G15gat), .A2(G22gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G1gat), .A2(G8gat), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n474_), .A2(new_n475_), .B1(KEYINPUT14), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n471_), .B(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G231gat), .A2(G233gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G57gat), .B(G64gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G71gat), .B(G78gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n481_), .A2(KEYINPUT11), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n480_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT74), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G127gat), .B(G155gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT16), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G183gat), .ZN(new_n492_));
  INV_X1    g291(.A(G211gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n489_), .B(new_n496_), .Z(new_n497_));
  INV_X1    g296(.A(new_n488_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(new_n495_), .A3(new_n494_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT65), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT6), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n502_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(G99gat), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n510_), .A2(KEYINPUT10), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(KEYINPUT10), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(KEYINPUT9), .A3(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT66), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n515_), .A2(KEYINPUT9), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n508_), .A2(new_n517_), .A3(new_n518_), .A4(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n513_), .B(new_n516_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT66), .B1(new_n522_), .B2(new_n519_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n524_));
  OR3_X1    g323(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n524_), .B(new_n525_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n514_), .A2(new_n515_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n521_), .B(new_n523_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G29gat), .B(G36gat), .ZN(new_n532_));
  INV_X1    g331(.A(G43gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G50gat), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G232gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT34), .ZN(new_n538_));
  INV_X1    g337(.A(G50gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n534_), .B(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT15), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT15), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n535_), .A2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n521_), .A2(new_n523_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n530_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT68), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT68), .B1(new_n529_), .B2(new_n530_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n545_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  OAI221_X1 g350(.A(new_n536_), .B1(KEYINPUT35), .B2(new_n538_), .C1(new_n544_), .C2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n538_), .A2(KEYINPUT35), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n544_), .A2(new_n551_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n555_), .A2(KEYINPUT35), .A3(new_n538_), .A4(new_n536_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G134gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n317_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT36), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n560_), .A2(new_n561_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n554_), .B(new_n556_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT37), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n563_), .A2(new_n569_), .A3(new_n566_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n469_), .A2(new_n500_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n478_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT75), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n478_), .A2(new_n535_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT75), .B1(new_n574_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n478_), .B(new_n535_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(G229gat), .A3(G233gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT76), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(G169gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(new_n296_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n586_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n579_), .A2(new_n581_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n545_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n547_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n529_), .A2(new_n530_), .A3(KEYINPUT68), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(KEYINPUT12), .A3(new_n487_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT64), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT12), .B1(new_n531_), .B2(new_n487_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n531_), .A2(new_n487_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n595_), .A2(new_n597_), .A3(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n531_), .B(new_n487_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n597_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(KEYINPUT69), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT71), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n605_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT13), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT72), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n572_), .A2(new_n590_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(G1gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n434_), .B(KEYINPUT101), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n615_), .A2(new_n590_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n469_), .A2(new_n625_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n567_), .A2(KEYINPUT103), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n567_), .A2(KEYINPUT103), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(new_n500_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n626_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(new_n434_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n623_), .B1(new_n619_), .B2(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(G8gat), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n438_), .A2(new_n402_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n618_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n636_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G8gat), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(KEYINPUT39), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(KEYINPUT39), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(new_n287_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n472_), .B1(new_n632_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT41), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n618_), .A2(new_n472_), .A3(new_n645_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1326gat));
  INV_X1    g448(.A(new_n358_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n473_), .B1(new_n632_), .B2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT42), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n618_), .A2(new_n473_), .A3(new_n650_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1327gat));
  INV_X1    g453(.A(new_n500_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n629_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n626_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G29gat), .B1(new_n658_), .B2(new_n434_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n468_), .A2(new_n287_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n435_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n663_), .A3(new_n571_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n571_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n469_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n624_), .A3(new_n500_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n667_), .A2(KEYINPUT44), .A3(new_n624_), .A4(new_n500_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(G29gat), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n659_), .B1(new_n672_), .B2(new_n620_), .ZN(G1328gat));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n626_), .A2(new_n674_), .A3(new_n636_), .A4(new_n656_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT45), .Z(new_n676_));
  NAND3_X1  g475(.A1(new_n670_), .A2(new_n636_), .A3(new_n671_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(G36gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT104), .B(KEYINPUT46), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n678_), .B(new_n679_), .Z(G1329gat));
  NAND2_X1  g479(.A1(KEYINPUT105), .A2(G43gat), .ZN(new_n681_));
  OR2_X1    g480(.A1(KEYINPUT105), .A2(G43gat), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n681_), .B(new_n682_), .C1(new_n657_), .C2(new_n287_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT106), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n670_), .A2(G43gat), .A3(new_n645_), .A4(new_n671_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT47), .ZN(G1330gat));
  AND3_X1   g486(.A1(new_n670_), .A2(new_n650_), .A3(new_n671_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n358_), .A2(G50gat), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT107), .ZN(new_n690_));
  OAI22_X1  g489(.A1(new_n688_), .A2(new_n539_), .B1(new_n657_), .B2(new_n690_), .ZN(G1331gat));
  NOR2_X1   g490(.A1(new_n615_), .A2(new_n590_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n572_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT108), .ZN(new_n694_));
  AOI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n620_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n617_), .A2(new_n590_), .A3(new_n469_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n631_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n415_), .B(new_n697_), .C1(new_n430_), .C2(new_n433_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n695_), .A2(new_n698_), .ZN(G1332gat));
  NAND3_X1  g498(.A1(new_n696_), .A2(new_n636_), .A3(new_n631_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G64gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT48), .ZN(new_n702_));
  INV_X1    g501(.A(G64gat), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n636_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n693_), .B2(new_n704_), .ZN(G1333gat));
  OR3_X1    g504(.A1(new_n693_), .A2(G71gat), .A3(new_n287_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n696_), .A2(new_n645_), .A3(new_n631_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G71gat), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n708_), .A2(KEYINPUT109), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(KEYINPUT109), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(KEYINPUT49), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT49), .B1(new_n709_), .B2(new_n710_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n706_), .B1(new_n711_), .B2(new_n712_), .ZN(G1334gat));
  OR3_X1    g512(.A1(new_n693_), .A2(G78gat), .A3(new_n358_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G78gat), .B1(new_n697_), .B2(new_n358_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n715_), .A2(KEYINPUT110), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(KEYINPUT110), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(KEYINPUT50), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT50), .B1(new_n716_), .B2(new_n717_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n718_), .B2(new_n719_), .ZN(G1335gat));
  NOR3_X1   g519(.A1(new_n615_), .A2(new_n655_), .A3(new_n590_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n667_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n434_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n696_), .A2(new_n656_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n620_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(G85gat), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n723_), .A2(G85gat), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT111), .ZN(G1336gat));
  AOI21_X1  g527(.A(G92gat), .B1(new_n724_), .B2(new_n636_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n636_), .A2(G92gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n722_), .B2(new_n730_), .ZN(G1337gat));
  OAI211_X1 g530(.A(new_n724_), .B(new_n645_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(KEYINPUT112), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n722_), .A2(new_n645_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n510_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT51), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n733_), .B(new_n737_), .C1(new_n510_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1338gat));
  AOI21_X1  g538(.A(new_n663_), .B1(new_n662_), .B2(new_n571_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n469_), .A2(KEYINPUT43), .A3(new_n665_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n650_), .B(new_n721_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n667_), .A2(KEYINPUT113), .A3(new_n650_), .A4(new_n721_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(G106gat), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT52), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n744_), .A2(new_n748_), .A3(G106gat), .A4(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n724_), .A2(new_n509_), .A3(new_n650_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n750_), .A2(new_n754_), .A3(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  NAND2_X1  g555(.A1(new_n580_), .A2(new_n576_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n575_), .A2(new_n578_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n586_), .B(new_n757_), .C1(new_n758_), .C2(new_n576_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(new_n589_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n605_), .A2(new_n611_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n601_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n595_), .A2(new_n600_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n603_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n595_), .A2(KEYINPUT55), .A3(new_n600_), .A4(new_n597_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n601_), .A2(KEYINPUT114), .A3(new_n762_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n765_), .A2(new_n767_), .A3(new_n768_), .A4(new_n769_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n770_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT56), .B1(new_n770_), .B2(new_n610_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n760_), .B(new_n761_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  INV_X1    g575(.A(new_n769_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n767_), .A2(new_n768_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT114), .B1(new_n601_), .B2(new_n762_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n780_), .B2(new_n611_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n770_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n783_), .A2(KEYINPUT58), .A3(new_n760_), .A4(new_n761_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n775_), .A2(new_n571_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n590_), .A2(new_n761_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n614_), .A2(new_n760_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n629_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT57), .B(new_n629_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n785_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n571_), .A2(new_n500_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n590_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n615_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n796_), .A2(KEYINPUT54), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(KEYINPUT54), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n793_), .A2(new_n500_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(new_n287_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n411_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n620_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT115), .ZN(new_n803_));
  NOR4_X1   g602(.A1(new_n799_), .A2(new_n287_), .A3(new_n411_), .A4(new_n725_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G113gat), .B1(new_n807_), .B2(new_n590_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n802_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n812_));
  NAND4_X1  g611(.A1(new_n800_), .A2(new_n801_), .A3(new_n620_), .A4(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n795_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n808_), .B1(G113gat), .B2(new_n814_), .ZN(G1340gat));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  INV_X1    g615(.A(G120gat), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(KEYINPUT60), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n615_), .A2(KEYINPUT60), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n817_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n818_), .B(new_n821_), .C1(new_n803_), .C2(new_n806_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n809_), .A2(new_n810_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n813_), .B1(new_n804_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n817_), .B1(new_n824_), .B2(new_n616_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n816_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n818_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n802_), .A2(KEYINPUT115), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n804_), .A2(new_n805_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n827_), .B(new_n820_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n617_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n830_), .B(KEYINPUT117), .C1(new_n831_), .C2(new_n817_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n826_), .A2(new_n832_), .ZN(G1341gat));
  AND3_X1   g632(.A1(new_n824_), .A2(G127gat), .A3(new_n655_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n807_), .A2(new_n655_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(KEYINPUT118), .A3(new_n207_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n500_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(G127gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n834_), .B1(new_n836_), .B2(new_n839_), .ZN(G1342gat));
  AOI21_X1  g639(.A(G134gat), .B1(new_n807_), .B2(new_n630_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT119), .B(G134gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n665_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(G1343gat));
  NOR2_X1   g643(.A1(new_n636_), .A2(new_n358_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NOR4_X1   g645(.A1(new_n799_), .A2(new_n645_), .A3(new_n725_), .A4(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n590_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n616_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g650(.A1(new_n793_), .A2(new_n500_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n797_), .A2(new_n798_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n645_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n620_), .A3(new_n845_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n500_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT120), .B1(new_n847_), .B2(new_n655_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT61), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n855_), .B2(new_n500_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n847_), .A2(KEYINPUT120), .A3(new_n655_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT61), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n859_), .A2(G155gat), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G155gat), .B1(new_n859_), .B2(new_n863_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1346gat));
  AOI21_X1  g665(.A(G162gat), .B1(new_n847_), .B2(new_n630_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n665_), .A2(new_n317_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n847_), .B2(new_n868_), .ZN(G1347gat));
  NAND2_X1  g668(.A1(new_n852_), .A2(new_n853_), .ZN(new_n870_));
  AOI211_X1 g669(.A(new_n620_), .B(new_n650_), .C1(new_n438_), .C2(new_n402_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n870_), .A2(new_n590_), .A3(new_n645_), .A4(new_n871_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(G169gat), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT122), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n872_), .A2(G169gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n873_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n872_), .A2(new_n879_), .A3(G169gat), .A4(new_n874_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n876_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n800_), .A2(new_n871_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n800_), .A2(new_n871_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT123), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n795_), .A2(new_n370_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n884_), .A2(new_n886_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n881_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT124), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n881_), .A2(new_n888_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1348gat));
  NOR3_X1   g692(.A1(new_n885_), .A2(new_n224_), .A3(new_n617_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n884_), .A2(new_n886_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n895_), .A2(new_n615_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n896_), .B2(new_n224_), .ZN(G1349gat));
  AOI21_X1  g696(.A(G183gat), .B1(new_n882_), .B2(new_n655_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n500_), .A2(new_n235_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(G1350gat));
  OAI21_X1  g700(.A(G190gat), .B1(new_n895_), .B2(new_n665_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n630_), .A2(new_n234_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n895_), .B2(new_n903_), .ZN(G1351gat));
  NAND3_X1  g703(.A1(new_n854_), .A2(new_n439_), .A3(new_n636_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n590_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n616_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n655_), .B1(new_n912_), .B2(new_n493_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT126), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n905_), .A2(new_n906_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n439_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n799_), .A2(new_n645_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(KEYINPUT125), .B1(new_n917_), .B2(new_n636_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n914_), .B1(new_n915_), .B2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT127), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n920_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923_));
  INV_X1    g722(.A(new_n920_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n907_), .A2(new_n923_), .A3(new_n924_), .A4(new_n914_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n921_), .A2(new_n922_), .A3(new_n925_), .ZN(G1354gat));
  AOI21_X1  g725(.A(G218gat), .B1(new_n907_), .B2(new_n630_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n907_), .A2(new_n571_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(G218gat), .B2(new_n928_), .ZN(G1355gat));
endmodule


