//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT78), .B(G176gat), .Z(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT22), .B1(new_n206_), .B2(KEYINPUT77), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n206_), .A2(KEYINPUT22), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n205_), .B(new_n207_), .C1(KEYINPUT77), .C2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT25), .B(G183gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n206_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n214_), .A2(new_n203_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n211_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G71gat), .B(G99gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(G43gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n220_), .B(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G127gat), .B(G134gat), .Z(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n223_), .B(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G227gat), .A2(G233gat), .ZN(new_n228_));
  INV_X1    g027(.A(G15gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT31), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n227_), .B(new_n232_), .Z(new_n233_));
  NAND2_X1  g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n234_), .B1(new_n235_), .B2(KEYINPUT1), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT80), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n238_), .B(new_n234_), .C1(new_n235_), .C2(KEYINPUT1), .ZN(new_n239_));
  AND2_X1   g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(KEYINPUT79), .A2(G141gat), .A3(G148gat), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n246_), .B(new_n247_), .C1(G141gat), .C2(G148gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT2), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT82), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT2), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n246_), .A2(new_n247_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(KEYINPUT81), .A3(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G141gat), .ZN(new_n262_));
  INV_X1    g061(.A(G148gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT81), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n255_), .A2(new_n258_), .A3(new_n261_), .A4(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT83), .A3(new_n234_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT83), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n240_), .B2(new_n235_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n250_), .A2(new_n273_), .A3(KEYINPUT84), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT84), .B1(new_n250_), .B2(new_n273_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT91), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT90), .B(KEYINPUT4), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n226_), .A4(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n269_), .A2(new_n271_), .ZN(new_n281_));
  NOR4_X1   g080(.A1(new_n265_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT81), .B1(new_n256_), .B2(new_n257_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n259_), .A2(new_n260_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n281_), .B1(new_n285_), .B2(new_n255_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n236_), .A2(KEYINPUT80), .B1(new_n241_), .B2(new_n240_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n248_), .B1(new_n287_), .B2(new_n239_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n280_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n250_), .A2(new_n273_), .A3(KEYINPUT84), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(new_n226_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n250_), .A2(new_n273_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(new_n226_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(KEYINPUT4), .A3(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n289_), .A2(new_n290_), .A3(new_n226_), .A4(new_n278_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT91), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n279_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT92), .B(KEYINPUT0), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT93), .ZN(new_n305_));
  XOR2_X1   g104(.A(G1gat), .B(G29gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G57gat), .B(G85gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n303_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT94), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n301_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(new_n309_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n303_), .A2(new_n312_), .A3(new_n310_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n205_), .ZN(new_n317_));
  XOR2_X1   g116(.A(KEYINPUT22), .B(G169gat), .Z(new_n318_));
  OAI211_X1 g117(.A(new_n204_), .B(new_n210_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n219_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G211gat), .B(G218gat), .Z(new_n321_));
  INV_X1    g120(.A(KEYINPUT21), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G197gat), .B(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n323_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(new_n321_), .A3(KEYINPUT21), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT20), .B1(new_n320_), .B2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n328_), .A2(new_n220_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G226gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT19), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n320_), .A2(new_n328_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n336_), .B(KEYINPUT20), .C1(new_n220_), .C2(new_n328_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G8gat), .B(G36gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT32), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n333_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n337_), .B2(new_n333_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n348_), .B2(new_n345_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n315_), .A2(new_n316_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n303_), .A2(KEYINPUT33), .A3(new_n310_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n313_), .B2(new_n309_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n335_), .A2(new_n338_), .A3(new_n344_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n344_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n291_), .A2(new_n299_), .A3(new_n293_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n309_), .B(new_n358_), .C1(new_n297_), .C2(new_n299_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n351_), .A2(new_n353_), .A3(new_n357_), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n350_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G228gat), .A2(G233gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n289_), .A2(new_n290_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n362_), .B(new_n328_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT86), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n243_), .A2(new_n249_), .B1(new_n267_), .B2(new_n272_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(new_n364_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n292_), .A2(KEYINPUT86), .A3(KEYINPUT29), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n328_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT87), .ZN(new_n371_));
  INV_X1    g170(.A(new_n362_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n371_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n365_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G78gat), .B(G106gat), .Z(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n378_), .B(new_n365_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT28), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n383_));
  AOI211_X1 g182(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n289_), .C2(new_n290_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT85), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT28), .B1(new_n276_), .B2(KEYINPUT29), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n363_), .A2(new_n382_), .A3(new_n364_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G22gat), .B(G50gat), .Z(new_n390_));
  AND3_X1   g189(.A1(new_n385_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n385_), .B2(new_n389_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n381_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n390_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n383_), .A2(new_n384_), .A3(KEYINPUT85), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n387_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n385_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(KEYINPUT88), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n380_), .B1(new_n393_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n398_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n401_), .A2(new_n381_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n361_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT27), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT96), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n354_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n344_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n348_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT95), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n348_), .A2(KEYINPUT95), .A3(new_n408_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n335_), .A2(new_n338_), .A3(KEYINPUT96), .A4(new_n344_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n407_), .A2(new_n411_), .A3(new_n412_), .A4(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n405_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n315_), .A2(new_n316_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n417_), .B(new_n418_), .C1(new_n400_), .C2(new_n402_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n233_), .B1(new_n404_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n403_), .A2(new_n417_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n233_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G29gat), .B(G36gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G43gat), .B(G50gat), .Z(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G43gat), .B(G50gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT15), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G15gat), .B(G22gat), .ZN(new_n434_));
  INV_X1    g233(.A(G1gat), .ZN(new_n435_));
  INV_X1    g234(.A(G8gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT14), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G1gat), .B(G8gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n428_), .A2(KEYINPUT15), .A3(new_n430_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n433_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n438_), .A2(new_n439_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n439_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n431_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G229gat), .A2(G233gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n446_), .B(KEYINPUT74), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n431_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n440_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n445_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n446_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n442_), .A2(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G113gat), .B(G141gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G169gat), .B(G197gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n455_), .B(new_n456_), .Z(new_n457_));
  NOR2_X1   g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n449_), .A2(new_n442_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n452_), .A2(new_n453_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n457_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT75), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT75), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n454_), .A2(new_n463_), .A3(new_n457_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n458_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT76), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n424_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468_));
  XOR2_X1   g267(.A(G85gat), .B(G92gat), .Z(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT6), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n472_));
  INV_X1    g271(.A(G99gat), .ZN(new_n473_));
  INV_X1    g272(.A(G106gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n471_), .B1(new_n478_), .B2(KEYINPUT64), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT64), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT8), .B(new_n469_), .C1(new_n479_), .C2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n470_), .B(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n469_), .B1(new_n484_), .B2(new_n477_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT8), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT10), .B(G99gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n474_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n469_), .A2(KEYINPUT9), .ZN(new_n490_));
  INV_X1    g289(.A(G85gat), .ZN(new_n491_));
  INV_X1    g290(.A(G92gat), .ZN(new_n492_));
  OR3_X1    g291(.A1(new_n491_), .A2(new_n492_), .A3(KEYINPUT9), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n489_), .A2(new_n490_), .A3(new_n471_), .A4(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n482_), .A2(new_n487_), .A3(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n433_), .A2(new_n441_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT35), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT34), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n495_), .A2(new_n496_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n482_), .A2(KEYINPUT65), .A3(new_n487_), .A4(new_n494_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n487_), .A2(new_n494_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n469_), .A2(KEYINPUT8), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n484_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n481_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n503_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n502_), .A2(new_n509_), .A3(new_n431_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n501_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n500_), .A2(new_n497_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n501_), .B(new_n510_), .C1(new_n497_), .C2(new_n500_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G190gat), .B(G218gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G134gat), .B(G162gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT69), .Z(new_n520_));
  NAND3_X1  g319(.A1(new_n513_), .A2(new_n514_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT70), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT70), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n513_), .A2(new_n523_), .A3(new_n514_), .A4(new_n520_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n513_), .A2(new_n514_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n517_), .B(KEYINPUT36), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT71), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n468_), .B1(new_n525_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n527_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n533_));
  AOI211_X1 g332(.A(KEYINPUT37), .B(new_n533_), .C1(new_n522_), .C2(new_n524_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G127gat), .B(G155gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT16), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G183gat), .B(G211gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n544_));
  XOR2_X1   g343(.A(G71gat), .B(G78gat), .Z(new_n545_));
  OR2_X1    g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n545_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT72), .ZN(new_n552_));
  INV_X1    g351(.A(new_n550_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n546_), .B(new_n553_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n551_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n552_), .B1(new_n551_), .B2(new_n554_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n440_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n548_), .A2(new_n547_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n553_), .B1(new_n558_), .B2(new_n546_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n554_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT72), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n440_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n551_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n542_), .B1(new_n557_), .B2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n540_), .A2(new_n541_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n557_), .A2(new_n566_), .A3(new_n564_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT73), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n557_), .A2(new_n564_), .A3(KEYINPUT73), .A4(new_n566_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n565_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n536_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n502_), .A2(new_n509_), .A3(new_n549_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n549_), .B1(new_n502_), .B2(new_n509_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G120gat), .B(G148gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT5), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n502_), .A2(new_n509_), .A3(new_n549_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n549_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n495_), .A2(KEYINPUT12), .A3(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT66), .B(KEYINPUT12), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n583_), .B(new_n585_), .C1(new_n576_), .C2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n577_), .B(new_n582_), .C1(new_n588_), .C2(new_n574_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT67), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n502_), .A2(new_n509_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n587_), .B1(new_n592_), .B2(new_n584_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n583_), .A2(new_n585_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n596_), .A3(new_n573_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n597_), .A2(KEYINPUT67), .A3(new_n577_), .A4(new_n582_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n591_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n577_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n581_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT68), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT13), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n599_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n572_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n467_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n418_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n435_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n380_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n391_), .A2(new_n392_), .A3(new_n381_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT88), .B1(new_n397_), .B2(new_n398_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n393_), .A2(new_n380_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n416_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n620_), .A2(new_n418_), .B1(new_n361_), .B2(new_n403_), .ZN(new_n621_));
  OAI22_X1  g420(.A1(new_n621_), .A2(new_n233_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n533_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n607_), .A2(new_n465_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n622_), .A2(new_n571_), .A3(new_n624_), .A4(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n418_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n612_), .A2(new_n613_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n614_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT97), .ZN(G1324gat));
  OAI21_X1  g429(.A(G8gat), .B1(new_n626_), .B2(new_n417_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT98), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(KEYINPUT98), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(KEYINPUT39), .A3(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n610_), .A2(new_n436_), .A3(new_n416_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n634_), .B(new_n635_), .C1(KEYINPUT39), .C2(new_n633_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1325gat));
  INV_X1    g437(.A(new_n233_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G15gat), .B1(new_n626_), .B2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT41), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n610_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1326gat));
  OAI21_X1  g442(.A(G22gat), .B1(new_n626_), .B2(new_n403_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT42), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n403_), .A2(G22gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n645_), .B1(new_n609_), .B2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(new_n571_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n625_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n530_), .A2(new_n534_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n622_), .B2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n651_), .B(new_n652_), .C1(new_n420_), .C2(new_n423_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n650_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(KEYINPUT44), .B(new_n650_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n418_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT100), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G29gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n661_), .A2(KEYINPUT100), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n607_), .A2(new_n571_), .A3(new_n624_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n467_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n418_), .A2(G29gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT101), .ZN(new_n668_));
  OAI22_X1  g467(.A1(new_n663_), .A2(new_n664_), .B1(new_n666_), .B2(new_n668_), .ZN(G1328gat));
  NOR3_X1   g468(.A1(new_n666_), .A2(G36gat), .A3(new_n417_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT45), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n658_), .A2(new_n416_), .A3(new_n659_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n672_), .A2(new_n673_), .A3(G36gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n672_), .B2(G36gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI211_X1 g477(.A(KEYINPUT46), .B(new_n671_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1329gat));
  AND2_X1   g479(.A1(new_n233_), .A2(G43gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n658_), .A2(new_n659_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n658_), .A2(KEYINPUT103), .A3(new_n659_), .A4(new_n681_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT104), .B(G43gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n666_), .B2(new_n639_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n685_), .A3(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g488(.A(new_n403_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G50gat), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n666_), .A2(new_n403_), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n660_), .A2(new_n691_), .B1(G50gat), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT105), .Z(G1331gat));
  INV_X1    g493(.A(G57gat), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n462_), .A2(new_n464_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n458_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n424_), .A2(new_n698_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n699_), .A2(new_n607_), .A3(new_n571_), .A4(new_n536_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n695_), .B1(new_n700_), .B2(new_n418_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT106), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n599_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n599_), .A2(new_n601_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n605_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n698_), .A2(KEYINPUT76), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT76), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n465_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n571_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n705_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n622_), .A2(new_n624_), .A3(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n711_), .A2(new_n695_), .A3(new_n418_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n702_), .A2(new_n712_), .ZN(G1332gat));
  OAI21_X1  g512(.A(G64gat), .B1(new_n711_), .B2(new_n417_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT48), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n417_), .A2(G64gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n700_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT107), .ZN(G1333gat));
  OAI21_X1  g517(.A(G71gat), .B1(new_n711_), .B2(new_n639_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT49), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n639_), .A2(G71gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n700_), .B2(new_n721_), .ZN(G1334gat));
  OAI21_X1  g521(.A(G78gat), .B1(new_n711_), .B2(new_n403_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT50), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n403_), .A2(G78gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n700_), .B2(new_n725_), .ZN(G1335gat));
  OR2_X1    g525(.A1(new_n653_), .A2(new_n655_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n705_), .A2(new_n698_), .A3(new_n571_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n418_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n699_), .A2(new_n607_), .A3(new_n648_), .A4(new_n623_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n491_), .A3(new_n611_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1336gat));
  OAI21_X1  g533(.A(G92gat), .B1(new_n729_), .B2(new_n417_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n492_), .A3(new_n416_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1337gat));
  NAND3_X1  g536(.A1(new_n732_), .A2(new_n233_), .A3(new_n488_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n727_), .A2(new_n233_), .A3(new_n728_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(new_n740_), .A3(G99gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n739_), .B2(G99gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g543(.A1(new_n732_), .A2(new_n474_), .A3(new_n690_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n727_), .A2(new_n690_), .A3(new_n728_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n747_), .A3(G106gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(G106gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n709_), .A2(new_n752_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n571_), .A2(new_n706_), .A3(KEYINPUT109), .A4(new_n708_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n753_), .B(new_n754_), .C1(new_n530_), .C2(new_n534_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT54), .B1(new_n607_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT109), .B1(new_n466_), .B2(new_n571_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n754_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n705_), .A2(new_n759_), .A3(new_n536_), .A4(new_n760_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n756_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n599_), .A2(new_n601_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n457_), .B1(new_n452_), .B2(new_n448_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n442_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n696_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT111), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n696_), .A2(new_n770_), .A3(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n764_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT55), .B1(new_n573_), .B2(KEYINPUT110), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n581_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(KEYINPUT55), .B2(new_n573_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n588_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n774_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n582_), .B1(new_n588_), .B2(new_n776_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n782_), .B(KEYINPUT56), .C1(new_n588_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(new_n698_), .A3(new_n599_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n623_), .B1(new_n773_), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n763_), .B1(new_n786_), .B2(KEYINPUT57), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n781_), .A2(new_n783_), .B1(new_n591_), .B2(new_n598_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n698_), .A2(new_n789_), .B1(new_n764_), .B2(new_n772_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT112), .B(new_n788_), .C1(new_n790_), .C2(new_n623_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n784_), .A2(KEYINPUT58), .A3(new_n599_), .A4(new_n772_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n789_), .A2(new_n772_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n652_), .B(new_n792_), .C1(new_n793_), .C2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n786_), .A2(KEYINPUT57), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n787_), .A2(new_n791_), .A3(new_n796_), .A4(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n762_), .B1(new_n798_), .B2(new_n648_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n403_), .A2(new_n611_), .A3(new_n417_), .A4(new_n233_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(G113gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n698_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n800_), .A2(KEYINPUT59), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n790_), .A2(new_n788_), .A3(new_n623_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n792_), .A2(new_n531_), .A3(new_n535_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n795_), .B1(new_n789_), .B2(new_n772_), .ZN(new_n807_));
  OAI22_X1  g606(.A1(new_n786_), .A2(KEYINPUT57), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n805_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n796_), .B(KEYINPUT114), .C1(KEYINPUT57), .C2(new_n786_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n571_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n804_), .B1(new_n812_), .B2(new_n762_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT59), .B1(new_n799_), .B2(new_n800_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n466_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n803_), .B1(new_n818_), .B2(new_n802_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT116), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n803_), .C1(new_n818_), .C2(new_n802_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1340gat));
  NOR2_X1   g622(.A1(new_n705_), .A2(KEYINPUT60), .ZN(new_n824_));
  MUX2_X1   g623(.A(new_n824_), .B(KEYINPUT60), .S(G120gat), .Z(new_n825_));
  NAND2_X1  g624(.A1(new_n801_), .A2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT117), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n813_), .A2(new_n814_), .A3(new_n607_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(G120gat), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1341gat));
  INV_X1    g629(.A(G127gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n801_), .A2(new_n831_), .A3(new_n571_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n816_), .A2(new_n817_), .A3(new_n648_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n831_), .ZN(G1342gat));
  INV_X1    g633(.A(G134gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n801_), .A2(new_n835_), .A3(new_n623_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n816_), .A2(new_n817_), .A3(new_n536_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n835_), .ZN(G1343gat));
  NOR2_X1   g637(.A1(new_n799_), .A2(new_n233_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n403_), .A2(new_n418_), .A3(new_n416_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n465_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT118), .B(G141gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1344gat));
  NOR2_X1   g643(.A1(new_n841_), .A2(new_n705_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT119), .B(G148gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1345gat));
  OR3_X1    g646(.A1(new_n841_), .A2(KEYINPUT120), .A3(new_n648_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT120), .B1(new_n841_), .B2(new_n648_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT61), .B(G155gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1346gat));
  INV_X1    g651(.A(new_n841_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n853_), .A2(G162gat), .A3(new_n652_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G162gat), .B1(new_n853_), .B2(new_n623_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n855_), .A2(KEYINPUT121), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(KEYINPUT121), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n854_), .B1(new_n856_), .B2(new_n857_), .ZN(G1347gat));
  NAND2_X1  g657(.A1(new_n810_), .A2(new_n811_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n762_), .B1(new_n859_), .B2(new_n648_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n611_), .A2(new_n417_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n403_), .A3(new_n233_), .ZN(new_n862_));
  OR3_X1    g661(.A1(new_n860_), .A2(KEYINPUT123), .A3(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT123), .B1(new_n860_), .B2(new_n862_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n465_), .A2(new_n318_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n862_), .A2(new_n465_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n868_), .B(new_n869_), .C1(new_n812_), .C2(new_n762_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n870_), .A2(G169gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n869_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT122), .B1(new_n860_), .B2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n867_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  AND4_X1   g673(.A1(new_n867_), .A2(new_n873_), .A3(G169gat), .A4(new_n870_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n866_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT124), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n878_), .B(new_n866_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1348gat));
  NAND2_X1  g679(.A1(new_n863_), .A2(new_n864_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n317_), .B1(new_n882_), .B2(new_n607_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n799_), .A2(new_n690_), .ZN(new_n884_));
  AND4_X1   g683(.A1(G176gat), .A2(new_n607_), .A3(new_n861_), .A4(new_n233_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1349gat));
  NOR2_X1   g685(.A1(new_n648_), .A2(new_n212_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  AND4_X1   g687(.A1(new_n233_), .A2(new_n884_), .A3(new_n571_), .A4(new_n861_), .ZN(new_n889_));
  OAI22_X1  g688(.A1(new_n881_), .A2(new_n888_), .B1(G183gat), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n881_), .B2(new_n536_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n623_), .A2(new_n213_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n881_), .B2(new_n894_), .ZN(G1351gat));
  AND3_X1   g694(.A1(new_n839_), .A2(new_n690_), .A3(new_n861_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n698_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT126), .B(G197gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n897_), .B2(new_n900_), .ZN(G1352gat));
  NAND2_X1  g700(.A1(new_n896_), .A2(new_n607_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g702(.A(new_n648_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT127), .Z(new_n905_));
  NAND2_X1  g704(.A1(new_n896_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  XOR2_X1   g706(.A(new_n906_), .B(new_n907_), .Z(G1354gat));
  INV_X1    g707(.A(G218gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n896_), .A2(new_n909_), .A3(new_n623_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n896_), .A2(new_n652_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n909_), .ZN(G1355gat));
endmodule


