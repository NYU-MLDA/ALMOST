//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT34), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n208_));
  OAI22_X1  g007(.A1(new_n208_), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT64), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT65), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G85gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n213_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n207_), .B1(new_n212_), .B2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT6), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT6), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n222_), .A2(new_n223_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n219_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n214_), .A2(new_n213_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n225_), .A2(new_n227_), .ZN(new_n240_));
  AOI211_X1 g039(.A(new_n231_), .B(new_n235_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT7), .ZN(new_n242_));
  INV_X1    g041(.A(G99gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n223_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n226_), .B1(G99gat), .B2(G106gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n224_), .A2(KEYINPUT6), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n236_), .B(new_n244_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n235_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n230_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n229_), .B1(new_n241_), .B2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G29gat), .B(G36gat), .Z(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT70), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G29gat), .B(G36gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G43gat), .B(G50gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n252_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n206_), .B1(new_n250_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT15), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n252_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n257_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n259_), .A2(KEYINPUT15), .A3(new_n260_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n250_), .A2(KEYINPUT68), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n229_), .B(new_n272_), .C1(new_n241_), .C2(new_n249_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(KEYINPUT71), .B(new_n206_), .C1(new_n250_), .C2(new_n261_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n264_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n205_), .B(new_n206_), .C1(new_n250_), .C2(new_n261_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n278_), .A2(new_n274_), .A3(KEYINPUT74), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT74), .B1(new_n278_), .B2(new_n274_), .ZN(new_n280_));
  OAI22_X1  g079(.A1(new_n205_), .A2(new_n276_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G190gat), .B(G218gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT72), .ZN(new_n283_));
  XOR2_X1   g082(.A(G134gat), .B(G162gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n281_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n285_), .B(KEYINPUT36), .Z(new_n289_));
  NAND2_X1  g088(.A1(new_n281_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n202_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n281_), .A2(new_n292_), .A3(new_n289_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(new_n281_), .B2(new_n289_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n202_), .B(new_n288_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n290_), .A2(KEYINPUT75), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n281_), .A2(new_n292_), .A3(new_n289_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n300_), .A2(KEYINPUT76), .A3(new_n202_), .A4(new_n288_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n291_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G155gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G183gat), .B(G211gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n307_), .A2(KEYINPUT17), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(KEYINPUT17), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G1gat), .B(G8gat), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G15gat), .B(G22gat), .Z(new_n313_));
  INV_X1    g112(.A(KEYINPUT14), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n314_), .B1(G1gat), .B2(G8gat), .ZN(new_n315_));
  OR3_X1    g114(.A1(new_n313_), .A2(KEYINPUT77), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT77), .B1(new_n313_), .B2(new_n315_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n317_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n312_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(new_n311_), .A3(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G231gat), .A2(G233gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(KEYINPUT67), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G57gat), .B(G64gat), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n328_), .B1(new_n329_), .B2(KEYINPUT11), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n329_), .A2(KEYINPUT11), .ZN(new_n332_));
  XOR2_X1   g131(.A(G71gat), .B(G78gat), .Z(new_n333_));
  NAND3_X1  g132(.A1(new_n329_), .A2(new_n328_), .A3(KEYINPUT11), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .A4(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(KEYINPUT11), .B2(new_n329_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n334_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n330_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n327_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n327_), .A2(new_n339_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n310_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n342_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(new_n340_), .A3(new_n308_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n302_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT80), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n335_), .A2(new_n338_), .A3(KEYINPUT12), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n271_), .A2(new_n273_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT12), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n247_), .A2(new_n248_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n231_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n247_), .A2(new_n230_), .A3(new_n248_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n353_), .A2(new_n354_), .B1(new_n219_), .B2(new_n228_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n351_), .B1(new_n355_), .B2(new_n339_), .ZN(new_n356_));
  AND2_X1   g155(.A1(G230gat), .A2(G233gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(new_n355_), .B2(new_n339_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n350_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n250_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n355_), .A2(new_n339_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n357_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G120gat), .B(G148gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT5), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G176gat), .B(G204gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n368_), .A2(KEYINPUT69), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n363_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT13), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n371_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n261_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G229gat), .A2(G233gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n322_), .A2(new_n324_), .A3(new_n270_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n378_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n322_), .A2(new_n324_), .A3(new_n261_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n376_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G113gat), .B(G141gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G169gat), .B(G197gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n384_), .B1(KEYINPUT81), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(KEYINPUT81), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n375_), .A2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT22), .B(G169gat), .ZN(new_n396_));
  INV_X1    g195(.A(G176gat), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT23), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(G183gat), .A3(G190gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT82), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G183gat), .A2(G190gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT23), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G183gat), .A2(G190gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n398_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G197gat), .B(G204gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT21), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n408_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G211gat), .B(G218gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  OR3_X1    g211(.A1(new_n407_), .A2(new_n411_), .A3(new_n408_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT24), .ZN(new_n417_));
  OR3_X1    g216(.A1(new_n395_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT25), .B(G183gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT26), .B(G190gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n416_), .A2(new_n417_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n418_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n403_), .A2(new_n400_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n406_), .A2(new_n415_), .A3(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT92), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G226gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT19), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT20), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(new_n427_), .B2(KEYINPUT92), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n398_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n425_), .B1(G183gat), .B2(G190gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n398_), .A2(new_n434_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n437_), .A2(new_n438_), .B1(new_n404_), .B2(new_n423_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(KEYINPUT91), .A3(new_n414_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT91), .B1(new_n439_), .B2(new_n414_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n428_), .B(new_n433_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n406_), .A2(new_n426_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n414_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n445_), .B(KEYINPUT20), .C1(new_n439_), .C2(new_n414_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n430_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G8gat), .B(G36gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT18), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G64gat), .B(G92gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(new_n447_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT27), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n427_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n442_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(new_n440_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT94), .B1(new_n457_), .B2(new_n431_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT94), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n441_), .A2(new_n442_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n459_), .B(new_n430_), .C1(new_n460_), .C2(new_n455_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n446_), .A2(new_n430_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n451_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n453_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G29gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(G85gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT0), .B(G57gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G127gat), .B(G134gat), .Z(new_n471_));
  XOR2_X1   g270(.A(G113gat), .B(G120gat), .Z(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G155gat), .B(G162gat), .Z(new_n475_));
  INV_X1    g274(.A(KEYINPUT1), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n478_));
  INV_X1    g277(.A(G141gat), .ZN(new_n479_));
  INV_X1    g278(.A(G148gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n479_), .A2(new_n480_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n477_), .A2(new_n478_), .A3(new_n481_), .A4(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT3), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n489_), .B(new_n490_), .C1(new_n482_), .C2(KEYINPUT2), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n475_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n484_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n474_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n484_), .A2(new_n492_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n473_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G225gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n494_), .A2(KEYINPUT4), .A3(new_n496_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n496_), .A2(KEYINPUT4), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n470_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n500_), .A2(new_n503_), .A3(new_n470_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n443_), .A2(new_n447_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n464_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT27), .B1(new_n509_), .B2(new_n452_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n465_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G22gat), .B(G50gat), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT28), .B1(new_n495_), .B2(KEYINPUT29), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT87), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT29), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n484_), .A2(new_n492_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n514_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n515_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n513_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n518_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT87), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n514_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n512_), .A3(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(new_n525_), .A3(KEYINPUT90), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G78gat), .B(G106gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT89), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n521_), .A2(new_n525_), .A3(KEYINPUT90), .A4(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n521_), .A2(new_n525_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT90), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n414_), .B1(new_n493_), .B2(new_n517_), .ZN(new_n536_));
  AND2_X1   g335(.A1(G228gat), .A2(G233gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT88), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n536_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(KEYINPUT88), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n532_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G71gat), .B(G99gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n544_), .B(G43gat), .Z(new_n545_));
  NAND2_X1  g344(.A1(new_n439_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G227gat), .A2(G233gat), .ZN(new_n547_));
  INV_X1    g346(.A(G15gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n550_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n552_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n398_), .A2(new_n434_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n557_), .A2(new_n436_), .A3(new_n435_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n401_), .A2(new_n403_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n424_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n545_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n546_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n556_), .B1(new_n546_), .B2(new_n562_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT84), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n562_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n561_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n567_));
  OAI22_X1  g366(.A1(new_n566_), .A2(new_n567_), .B1(new_n555_), .B2(new_n554_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT84), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n546_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n565_), .A2(new_n473_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n473_), .B1(new_n565_), .B2(new_n571_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n529_), .A2(new_n535_), .A3(new_n541_), .A4(new_n531_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n543_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT85), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n563_), .A2(new_n564_), .A3(KEYINPUT84), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n569_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n474_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n565_), .A2(new_n571_), .A3(new_n473_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT85), .A3(new_n582_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n543_), .A2(new_n575_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n511_), .B1(new_n576_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n543_), .A2(new_n575_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n505_), .A2(KEYINPUT33), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n497_), .A2(new_n499_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n469_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n501_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT33), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n504_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n588_), .A2(new_n593_), .A3(new_n509_), .A4(new_n452_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n451_), .A2(KEYINPUT32), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n463_), .A2(new_n596_), .ZN(new_n597_));
  OAI22_X1  g396(.A1(new_n505_), .A2(new_n506_), .B1(new_n508_), .B2(new_n596_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n578_), .A2(new_n583_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n587_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n394_), .B1(new_n585_), .B2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n348_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(G1gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n507_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n606_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n300_), .A2(new_n288_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n585_), .B2(new_n601_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n346_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n393_), .A4(new_n375_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT96), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n614_), .A2(new_n507_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n607_), .B(new_n608_), .C1(new_n604_), .C2(new_n615_), .ZN(G1324gat));
  NOR2_X1   g415(.A1(new_n465_), .A2(new_n510_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G8gat), .B1(new_n613_), .B2(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n618_), .A2(KEYINPUT97), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(KEYINPUT97), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(KEYINPUT39), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(G8gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n617_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n603_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n621_), .B(new_n624_), .C1(KEYINPUT39), .C2(new_n620_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g425(.A(new_n600_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n548_), .B1(new_n614_), .B2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT41), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n603_), .A2(new_n548_), .A3(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1326gat));
  INV_X1    g430(.A(G22gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n614_), .B2(new_n586_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT42), .Z(new_n634_));
  NAND2_X1  g433(.A1(new_n586_), .A2(new_n632_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT98), .Z(new_n636_));
  NAND2_X1  g435(.A1(new_n603_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(G1327gat));
  NOR2_X1   g437(.A1(new_n612_), .A2(new_n609_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n602_), .A2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT101), .Z(new_n641_));
  INV_X1    g440(.A(G29gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n507_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n585_), .A2(new_n601_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT43), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(new_n302_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT99), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n644_), .A2(new_n648_), .A3(new_n645_), .A4(new_n302_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n644_), .A2(new_n302_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT43), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n647_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n394_), .A2(new_n612_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n652_), .A2(KEYINPUT44), .A3(new_n653_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(KEYINPUT100), .A3(new_n507_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G29gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT100), .B1(new_n658_), .B2(new_n507_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n643_), .B1(new_n660_), .B2(new_n661_), .ZN(G1328gat));
  INV_X1    g461(.A(G36gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n641_), .A2(new_n663_), .A3(new_n623_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT45), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n656_), .A2(new_n623_), .A3(new_n657_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n663_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n665_), .B(KEYINPUT46), .C1(new_n666_), .C2(new_n663_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1329gat));
  AND2_X1   g470(.A1(new_n574_), .A2(G43gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n641_), .A2(new_n627_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT102), .B(G43gat), .ZN(new_n674_));
  AOI22_X1  g473(.A1(new_n658_), .A2(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g475(.A(G50gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n641_), .A2(new_n677_), .A3(new_n586_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n656_), .A2(new_n586_), .A3(new_n657_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n679_), .A2(KEYINPUT103), .A3(G50gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT103), .B1(new_n679_), .B2(G50gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT104), .B(new_n678_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1331gat));
  NAND4_X1  g485(.A1(new_n611_), .A2(new_n612_), .A3(new_n392_), .A4(new_n374_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n507_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G57gat), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n393_), .B1(new_n585_), .B2(new_n601_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n375_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n348_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n688_), .A2(G57gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n689_), .B1(new_n695_), .B2(new_n696_), .ZN(G1332gat));
  OAI21_X1  g496(.A(G64gat), .B1(new_n687_), .B2(new_n617_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT48), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n617_), .A2(G64gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n695_), .B2(new_n700_), .ZN(G1333gat));
  OAI21_X1  g500(.A(G71gat), .B1(new_n687_), .B2(new_n600_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n600_), .A2(G71gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n695_), .B2(new_n705_), .ZN(G1334gat));
  OAI21_X1  g505(.A(G78gat), .B1(new_n687_), .B2(new_n587_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT50), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n587_), .A2(G78gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n695_), .B2(new_n709_), .ZN(G1335gat));
  NAND2_X1  g509(.A1(new_n694_), .A2(new_n639_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G85gat), .B1(new_n712_), .B2(new_n507_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n346_), .A2(new_n392_), .A3(new_n374_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n652_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n652_), .A2(new_n715_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n714_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n688_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT108), .Z(new_n720_));
  AOI21_X1  g519(.A(new_n713_), .B1(new_n718_), .B2(new_n720_), .ZN(G1336gat));
  NAND3_X1  g520(.A1(new_n712_), .A2(new_n213_), .A3(new_n623_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n718_), .A2(new_n623_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n213_), .ZN(G1337gat));
  NAND2_X1  g523(.A1(new_n718_), .A2(new_n627_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n574_), .A2(new_n222_), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n725_), .A2(G99gat), .B1(new_n712_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(G1338gat));
  AND4_X1   g528(.A1(new_n223_), .A2(new_n694_), .A3(new_n586_), .A4(new_n639_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n714_), .A2(new_n587_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n223_), .B1(new_n652_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT52), .Z(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n732_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n732_), .B2(new_n735_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1339gat));
  INV_X1    g538(.A(new_n302_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT54), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n346_), .A2(new_n374_), .A3(new_n393_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n740_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n740_), .B2(new_n742_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n377_), .A2(new_n381_), .A3(new_n379_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n378_), .B1(new_n382_), .B2(new_n376_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n387_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n388_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n749_));
  OR3_X1    g548(.A1(new_n748_), .A2(new_n749_), .A3(KEYINPUT113), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT113), .B1(new_n748_), .B2(new_n749_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n363_), .A2(new_n367_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n751_), .A3(new_n753_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n350_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n355_), .A2(new_n339_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n350_), .A2(new_n756_), .A3(new_n356_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n755_), .A2(KEYINPUT55), .B1(new_n757_), .B2(new_n357_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT111), .B1(new_n359_), .B2(new_n760_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n359_), .A2(KEYINPUT111), .A3(new_n760_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n758_), .B(new_n759_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n359_), .A2(new_n760_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n359_), .A2(KEYINPUT111), .A3(new_n760_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n759_), .B1(new_n769_), .B2(new_n758_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n367_), .B1(new_n764_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n758_), .B1(new_n762_), .B2(new_n761_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT112), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n763_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n367_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n754_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n302_), .B1(new_n778_), .B2(KEYINPUT58), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n750_), .A2(new_n751_), .A3(new_n753_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT56), .B1(new_n776_), .B2(new_n367_), .ZN(new_n781_));
  AOI211_X1 g580(.A(new_n772_), .B(new_n368_), .C1(new_n775_), .C2(new_n763_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n780_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT114), .B1(new_n779_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n784_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n778_), .A2(KEYINPUT58), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .A4(new_n302_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n753_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n750_), .A2(new_n751_), .A3(new_n370_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n609_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n791_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n610_), .B1(new_n799_), .B2(new_n793_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT57), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n786_), .A2(new_n790_), .A3(new_n797_), .A4(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n612_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n800_), .A2(KEYINPUT57), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n796_), .B(new_n610_), .C1(new_n799_), .C2(new_n793_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(KEYINPUT115), .A3(new_n790_), .A4(new_n786_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n745_), .B1(new_n804_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n617_), .A2(new_n507_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n576_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n809_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OR3_X1    g613(.A1(new_n814_), .A2(G113gat), .A3(new_n392_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n812_), .A2(KEYINPUT59), .ZN(new_n816_));
  INV_X1    g615(.A(new_n745_), .ZN(new_n817_));
  OAI22_X1  g616(.A1(new_n779_), .A2(new_n785_), .B1(new_n800_), .B2(KEYINPUT57), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n806_), .B1(new_n818_), .B2(KEYINPUT116), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n797_), .B(new_n820_), .C1(new_n785_), .C2(new_n779_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n612_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n817_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  AOI211_X1 g623(.A(KEYINPUT117), .B(new_n612_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n816_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT59), .B1(new_n809_), .B2(new_n812_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n393_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(G113gat), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n815_), .A2(new_n829_), .ZN(G1340gat));
  NAND2_X1  g629(.A1(new_n802_), .A2(new_n803_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n808_), .A3(new_n346_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n817_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n812_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT118), .B(G120gat), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n375_), .B2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n833_), .A2(new_n834_), .A3(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n826_), .A2(new_n839_), .A3(new_n827_), .A4(new_n374_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n837_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n813_), .A2(new_n835_), .A3(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1341gat));
  AOI21_X1  g642(.A(G127gat), .B1(new_n813_), .B2(new_n612_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n826_), .A2(new_n827_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n612_), .A2(G127gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT119), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n844_), .B1(new_n845_), .B2(new_n847_), .ZN(G1342gat));
  OR3_X1    g647(.A1(new_n814_), .A2(G134gat), .A3(new_n609_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n826_), .A2(new_n302_), .A3(new_n827_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(G134gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1343gat));
  XNOR2_X1  g651(.A(KEYINPUT121), .B(G141gat), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n810_), .A2(new_n627_), .A3(new_n587_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT120), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n809_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n855_), .B1(new_n859_), .B2(new_n393_), .ZN(new_n860_));
  NOR4_X1   g659(.A1(new_n809_), .A2(KEYINPUT122), .A3(new_n392_), .A4(new_n858_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n854_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n833_), .A2(new_n857_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT122), .B1(new_n863_), .B2(new_n392_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n855_), .A3(new_n393_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n853_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n866_), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n859_), .A2(new_n374_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT123), .B(G148gat), .Z(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1345gat));
  NAND2_X1  g669(.A1(new_n859_), .A2(new_n612_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  OR3_X1    g672(.A1(new_n863_), .A2(G162gat), .A3(new_n609_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G162gat), .B1(new_n863_), .B2(new_n740_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1347gat));
  NOR3_X1   g675(.A1(new_n617_), .A2(new_n600_), .A3(new_n507_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n586_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n393_), .B(new_n879_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(G169gat), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n824_), .A2(new_n825_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n884_), .A2(new_n396_), .A3(new_n393_), .A4(new_n879_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n880_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n885_), .A3(new_n886_), .ZN(G1348gat));
  NAND3_X1  g686(.A1(new_n877_), .A2(G176gat), .A3(new_n374_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n809_), .A2(new_n586_), .A3(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n884_), .A2(new_n374_), .A3(new_n879_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n397_), .ZN(G1349gat));
  NOR2_X1   g690(.A1(new_n346_), .A2(new_n419_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n879_), .B(new_n892_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n878_), .A2(new_n346_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n833_), .A2(new_n587_), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G183gat), .B1(new_n897_), .B2(KEYINPUT124), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n894_), .B1(new_n898_), .B2(new_n900_), .ZN(G1350gat));
  NAND3_X1  g700(.A1(new_n884_), .A2(new_n302_), .A3(new_n879_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G190gat), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n884_), .A2(new_n610_), .A3(new_n420_), .A4(new_n879_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1351gat));
  NAND2_X1  g704(.A1(new_n584_), .A2(new_n688_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n623_), .B1(new_n906_), .B2(KEYINPUT125), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n809_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n393_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n833_), .A2(new_n911_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n375_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1353gat));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  NOR4_X1   g720(.A1(new_n916_), .A2(new_n346_), .A3(new_n920_), .A4(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n913_), .A2(new_n612_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n920_), .ZN(G1354gat));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n913_), .B2(new_n302_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n609_), .A2(G218gat), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n833_), .A2(new_n911_), .A3(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT127), .B1(new_n926_), .B2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G218gat), .B1(new_n916_), .B2(new_n740_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n913_), .A2(new_n927_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n929_), .A2(new_n933_), .ZN(G1355gat));
endmodule


