//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G183gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT80), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G190gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT79), .B(G183gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT25), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n206_), .A3(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT81), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(KEYINPUT81), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT24), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT23), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT82), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n216_), .B(new_n218_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n212_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n207_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n218_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n220_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n229_), .B(KEYINPUT22), .C1(new_n230_), .C2(new_n214_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232_));
  OAI211_X1 g031(.A(KEYINPUT84), .B(G169gat), .C1(new_n232_), .C2(KEYINPUT83), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n230_), .B1(new_n214_), .B2(KEYINPUT22), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n231_), .A2(new_n233_), .A3(new_n215_), .A4(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n227_), .A2(new_n228_), .A3(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G15gat), .B(G43gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT86), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n224_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n222_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n236_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n238_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(G71gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G99gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n240_), .A2(new_n243_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n252_));
  OR3_X1    g051(.A1(new_n251_), .A2(new_n252_), .A3(KEYINPUT87), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT87), .B1(new_n251_), .B2(new_n252_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G127gat), .B(G134gat), .Z(new_n255_));
  XOR2_X1   g054(.A(G113gat), .B(G120gat), .Z(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT31), .Z(new_n258_));
  NAND3_X1  g057(.A1(new_n253_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  OAI211_X1 g059(.A(KEYINPUT87), .B(new_n260_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT28), .B(G22gat), .ZN(new_n263_));
  INV_X1    g062(.A(G50gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT90), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT88), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n268_), .A2(new_n269_), .A3(KEYINPUT1), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(new_n268_), .B2(KEYINPUT1), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n272_));
  OR2_X1    g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .A4(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G141gat), .B(G148gat), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT2), .ZN(new_n277_));
  INV_X1    g076(.A(G141gat), .ZN(new_n278_));
  INV_X1    g077(.A(G148gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(KEYINPUT89), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(KEYINPUT89), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n283_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n273_), .A2(new_n268_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n276_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n267_), .B1(new_n289_), .B2(KEYINPUT29), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT92), .ZN(new_n291_));
  INV_X1    g090(.A(new_n289_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n266_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n290_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G204gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(G197gat), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT91), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(KEYINPUT91), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n296_), .A2(G197gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(KEYINPUT21), .ZN(new_n302_));
  XOR2_X1   g101(.A(G211gat), .B(G218gat), .Z(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n297_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n304_), .B2(KEYINPUT21), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n303_), .A2(KEYINPUT21), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n301_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(G228gat), .A3(G233gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G228gat), .A2(G233gat), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n309_), .B(new_n312_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n295_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT93), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT93), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n295_), .A2(new_n311_), .A3(new_n316_), .A4(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n290_), .A2(new_n294_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(new_n291_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G78gat), .B(G106gat), .Z(new_n322_));
  INV_X1    g121(.A(new_n320_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n321_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n322_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n262_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n262_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n321_), .A2(new_n324_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n322_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n332_), .A3(new_n325_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G8gat), .B(G36gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT18), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G64gat), .B(G92gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n335_), .B(new_n336_), .Z(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT19), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n309_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n224_), .B2(new_n236_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n218_), .A2(new_n216_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT95), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n213_), .B1(G169gat), .B2(G176gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT94), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n346_), .A2(new_n347_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT25), .B(G183gat), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n348_), .A2(new_n349_), .B1(new_n206_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n345_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n218_), .B1(G183gat), .B2(G190gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(KEYINPUT22), .B(G169gat), .Z(new_n354_));
  OAI211_X1 g153(.A(new_n353_), .B(new_n228_), .C1(G176gat), .C2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT20), .B1(new_n356_), .B2(new_n309_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n341_), .B1(new_n343_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n359_), .B1(new_n356_), .B2(new_n309_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n224_), .A2(new_n342_), .A3(new_n236_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n340_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n338_), .B1(new_n358_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT98), .B(KEYINPUT20), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n343_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT99), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n309_), .B1(new_n356_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(new_n369_), .B2(new_n356_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n341_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n360_), .A2(new_n361_), .A3(new_n341_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n365_), .B1(new_n374_), .B2(new_n337_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n358_), .A2(new_n362_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(new_n337_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n364_), .B1(new_n377_), .B2(new_n363_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n257_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n292_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n289_), .A2(new_n257_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n382_), .B(KEYINPUT4), .C1(KEYINPUT96), .C2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT96), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n289_), .A2(new_n385_), .A3(new_n386_), .A4(new_n257_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n380_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n380_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G1gat), .B(G29gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G85gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT0), .B(G57gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT100), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n395_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n391_), .A2(KEYINPUT100), .A3(new_n396_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n379_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n328_), .A2(new_n333_), .A3(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n384_), .A2(new_n380_), .A3(new_n387_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n382_), .A2(new_n389_), .A3(new_n383_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n406_), .A2(new_n396_), .A3(new_n407_), .ZN(new_n408_));
  OR3_X1    g207(.A1(new_n377_), .A2(new_n363_), .A3(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n399_), .B(KEYINPUT33), .Z(new_n410_));
  NAND2_X1  g209(.A1(new_n337_), .A2(KEYINPUT32), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT97), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n376_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n376_), .A2(KEYINPUT97), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n413_), .A2(new_n374_), .B1(new_n414_), .B2(new_n411_), .ZN(new_n415_));
  OAI22_X1  g214(.A1(new_n409_), .A2(new_n410_), .B1(new_n415_), .B2(new_n402_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n332_), .A2(new_n325_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n262_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n405_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G230gat), .A2(G233gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n420_), .B(KEYINPUT64), .Z(new_n421_));
  XOR2_X1   g220(.A(KEYINPUT10), .B(G99gat), .Z(new_n422_));
  INV_X1    g221(.A(G106gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G99gat), .A2(G106gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT6), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(G99gat), .A3(G106gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G85gat), .A2(G92gat), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n430_), .A2(KEYINPUT9), .ZN(new_n431_));
  OR2_X1    g230(.A1(G85gat), .A2(G92gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(KEYINPUT9), .A3(new_n430_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n424_), .A2(new_n429_), .A3(new_n431_), .A4(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT7), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(new_n247_), .A3(new_n423_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT65), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT65), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n440_), .A2(new_n436_), .A3(new_n247_), .A4(new_n423_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n438_), .A2(new_n429_), .A3(new_n439_), .A4(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n432_), .A2(new_n430_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(KEYINPUT66), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT8), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT8), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(new_n447_), .A3(new_n444_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n435_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G57gat), .B(G64gat), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n452_));
  XOR2_X1   g251(.A(G71gat), .B(G78gat), .Z(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n452_), .A2(new_n453_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n449_), .A2(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n442_), .A2(new_n447_), .A3(new_n444_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n447_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n434_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n456_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n421_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n462_), .A3(KEYINPUT12), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT12), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n460_), .A2(new_n465_), .A3(new_n461_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n463_), .B1(new_n467_), .B2(new_n421_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G120gat), .B(G148gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT5), .ZN(new_n470_));
  XOR2_X1   g269(.A(G176gat), .B(G204gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n468_), .A2(new_n473_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(KEYINPUT13), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT13), .B1(new_n474_), .B2(new_n475_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480_));
  INV_X1    g279(.A(G1gat), .ZN(new_n481_));
  INV_X1    g280(.A(G8gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G1gat), .B(G8gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G29gat), .B(G36gat), .Z(new_n487_));
  XOR2_X1   g286(.A(G43gat), .B(G50gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n486_), .B(new_n493_), .Z(new_n494_));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT15), .B1(new_n489_), .B2(new_n492_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n486_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n486_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n493_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n504_), .A3(new_n495_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n497_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G113gat), .B(G141gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT78), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G169gat), .B(G197gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(new_n510_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n479_), .A2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n419_), .A2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n434_), .B(new_n493_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT34), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(KEYINPUT35), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n493_), .B(new_n498_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n521_), .B1(new_n449_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n460_), .A2(KEYINPUT67), .A3(new_n501_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n520_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n518_), .A2(KEYINPUT35), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT68), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n516_), .A2(new_n519_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n460_), .A2(KEYINPUT67), .A3(new_n501_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT67), .B1(new_n460_), .B2(new_n501_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT68), .ZN(new_n532_));
  INV_X1    g331(.A(new_n526_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n526_), .B(KEYINPUT70), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n528_), .B(new_n535_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n523_), .A2(new_n524_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n539_), .A2(KEYINPUT71), .A3(new_n528_), .A4(new_n535_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n527_), .A2(new_n534_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G190gat), .B(G218gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT69), .ZN(new_n543_));
  XOR2_X1   g342(.A(G134gat), .B(G162gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT36), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT72), .B1(new_n541_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n527_), .A2(new_n534_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n538_), .A2(new_n540_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT72), .ZN(new_n551_));
  INV_X1    g350(.A(new_n546_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n545_), .A2(KEYINPUT36), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n541_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n547_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(KEYINPUT37), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n550_), .A2(new_n552_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n559_), .A2(new_n555_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n557_), .B1(new_n556_), .B2(KEYINPUT37), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G127gat), .B(G155gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT76), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT17), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n486_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(new_n456_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n575_), .A2(new_n570_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT77), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n565_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n515_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT101), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n481_), .A3(new_n403_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT38), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n584_), .A2(KEYINPUT38), .A3(new_n481_), .A4(new_n403_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n560_), .B1(new_n405_), .B2(new_n418_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n579_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n514_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n481_), .B1(new_n591_), .B2(new_n403_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT102), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(new_n588_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT103), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(G1324gat));
  NAND3_X1  g395(.A1(new_n584_), .A2(new_n482_), .A3(new_n379_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n482_), .B1(new_n591_), .B2(new_n379_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g402(.A(G15gat), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n591_), .B2(new_n329_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT41), .ZN(new_n606_));
  INV_X1    g405(.A(new_n583_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n604_), .A3(new_n329_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(G1326gat));
  INV_X1    g408(.A(G22gat), .ZN(new_n610_));
  INV_X1    g409(.A(new_n417_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n591_), .B2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT42), .Z(new_n613_));
  NAND3_X1  g412(.A1(new_n607_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1327gat));
  INV_X1    g414(.A(new_n560_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n580_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n515_), .A2(new_n617_), .ZN(new_n618_));
  OR3_X1    g417(.A1(new_n618_), .A2(G29gat), .A3(new_n402_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n419_), .A2(new_n565_), .A3(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(new_n581_), .ZN(new_n623_));
  OR2_X1    g422(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n405_), .A2(new_n418_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n556_), .A2(KEYINPUT37), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT73), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n562_), .A3(new_n558_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n620_), .B(new_n624_), .C1(new_n625_), .C2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n623_), .A2(new_n514_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT106), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n623_), .A2(new_n629_), .A3(KEYINPUT44), .A4(new_n514_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n403_), .A4(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(G29gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n632_), .A2(new_n403_), .A3(new_n634_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT106), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT107), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  AND4_X1   g438(.A1(KEYINPUT107), .A2(new_n638_), .A3(G29gat), .A4(new_n635_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n619_), .B1(new_n639_), .B2(new_n640_), .ZN(G1328gat));
  INV_X1    g440(.A(new_n379_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n618_), .A2(G36gat), .A3(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT45), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n632_), .A2(new_n379_), .A3(new_n634_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G36gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1329gat));
  NAND4_X1  g448(.A1(new_n632_), .A2(G43gat), .A3(new_n329_), .A4(new_n634_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT108), .ZN(new_n651_));
  INV_X1    g450(.A(new_n618_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G43gat), .B1(new_n652_), .B2(new_n329_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(KEYINPUT108), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT47), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT47), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n651_), .A2(new_n657_), .A3(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1330gat));
  AND3_X1   g458(.A1(new_n632_), .A2(new_n611_), .A3(new_n634_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n611_), .A2(new_n264_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT109), .ZN(new_n662_));
  OAI22_X1  g461(.A1(new_n660_), .A2(new_n264_), .B1(new_n618_), .B2(new_n662_), .ZN(G1331gat));
  INV_X1    g462(.A(new_n479_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n513_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n589_), .A2(new_n580_), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G57gat), .B1(new_n667_), .B2(new_n402_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT110), .B1(new_n625_), .B2(new_n665_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n665_), .B1(new_n405_), .B2(new_n418_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n664_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n672_), .A3(new_n582_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n402_), .A2(G57gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n668_), .B1(new_n673_), .B2(new_n674_), .ZN(G1332gat));
  OAI21_X1  g474(.A(G64gat), .B1(new_n667_), .B2(new_n642_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT48), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n642_), .A2(G64gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n673_), .B2(new_n678_), .ZN(G1333gat));
  OAI21_X1  g478(.A(G71gat), .B1(new_n667_), .B2(new_n262_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT49), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n329_), .A2(new_n245_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n673_), .B2(new_n682_), .ZN(G1334gat));
  OAI21_X1  g482(.A(G78gat), .B1(new_n667_), .B2(new_n417_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT50), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n417_), .A2(G78gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n673_), .B2(new_n686_), .ZN(G1335gat));
  NAND3_X1  g486(.A1(new_n669_), .A2(new_n672_), .A3(new_n617_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT111), .Z(new_n689_));
  INV_X1    g488(.A(G85gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n403_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n623_), .A2(new_n629_), .A3(new_n666_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G85gat), .B1(new_n692_), .B2(new_n402_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1336gat));
  AOI21_X1  g493(.A(G92gat), .B1(new_n689_), .B2(new_n379_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n379_), .A2(G92gat), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT112), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n695_), .B1(new_n696_), .B2(new_n698_), .ZN(G1337gat));
  NAND3_X1  g498(.A1(new_n689_), .A2(new_n422_), .A3(new_n329_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G99gat), .B1(new_n692_), .B2(new_n262_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT51), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT51), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n700_), .A2(new_n704_), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1338gat));
  OAI21_X1  g505(.A(G106gat), .B1(new_n692_), .B2(new_n417_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT52), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n689_), .A2(new_n423_), .A3(new_n611_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n708_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1339gat));
  NOR2_X1   g512(.A1(new_n479_), .A2(new_n665_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n580_), .B(new_n714_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT54), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT54), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n628_), .A2(new_n717_), .A3(new_n580_), .A4(new_n714_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n563_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n494_), .A2(new_n495_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n502_), .A2(new_n504_), .A3(new_n496_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n510_), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT114), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n511_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n724_), .B2(new_n723_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(new_n475_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n729_));
  INV_X1    g528(.A(new_n421_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n464_), .A2(new_n730_), .A3(new_n466_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT55), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n467_), .A2(new_n421_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n467_), .A2(KEYINPUT55), .A3(new_n421_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n473_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n729_), .B1(new_n736_), .B2(KEYINPUT56), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(KEYINPUT56), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n736_), .A2(new_n729_), .A3(KEYINPUT56), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n728_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT58), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n728_), .B(KEYINPUT58), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n720_), .A2(new_n743_), .A3(new_n744_), .A4(new_n627_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n513_), .B1(new_n468_), .B2(new_n473_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n736_), .A2(KEYINPUT56), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n748_), .B(new_n473_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n474_), .A2(new_n475_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n727_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT57), .B1(new_n753_), .B2(new_n616_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT57), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n755_), .B(new_n560_), .C1(new_n750_), .C2(new_n752_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n590_), .B1(new_n745_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT116), .B1(new_n719_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n745_), .A2(new_n757_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n579_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n716_), .A2(new_n718_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n761_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n611_), .A2(new_n262_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n379_), .A2(new_n402_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n759_), .A2(new_n764_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT117), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n759_), .A2(new_n764_), .A3(new_n770_), .A4(new_n767_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n769_), .A2(new_n665_), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(G113gat), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n772_), .A2(KEYINPUT118), .A3(new_n773_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT119), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n768_), .A2(KEYINPUT59), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n767_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n760_), .A2(new_n581_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(new_n763_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n778_), .B1(new_n779_), .B2(new_n784_), .ZN(new_n785_));
  AOI211_X1 g584(.A(KEYINPUT119), .B(new_n783_), .C1(new_n768_), .C2(KEYINPUT59), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n665_), .A2(G113gat), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT120), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n776_), .A2(new_n777_), .B1(new_n787_), .B2(new_n789_), .ZN(G1340gat));
  INV_X1    g589(.A(KEYINPUT60), .ZN(new_n791_));
  AOI21_X1  g590(.A(G120gat), .B1(new_n479_), .B2(new_n791_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT121), .Z(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n791_), .B2(G120gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n769_), .A2(new_n771_), .A3(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT122), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n779_), .A2(new_n479_), .A3(new_n784_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(G120gat), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1341gat));
  INV_X1    g598(.A(G127gat), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n769_), .A2(new_n800_), .A3(new_n580_), .A4(new_n771_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n785_), .A2(new_n786_), .A3(new_n579_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n800_), .ZN(G1342gat));
  INV_X1    g602(.A(G134gat), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n769_), .A2(new_n804_), .A3(new_n560_), .A4(new_n771_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n785_), .A2(new_n786_), .A3(new_n628_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n804_), .ZN(G1343gat));
  AND2_X1   g606(.A1(new_n759_), .A2(new_n764_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n808_), .A2(new_n611_), .A3(new_n262_), .A4(new_n766_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n513_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT123), .B(G141gat), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(G1344gat));
  NOR2_X1   g611(.A1(new_n809_), .A2(new_n664_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(new_n279_), .ZN(G1345gat));
  NOR2_X1   g613(.A1(new_n809_), .A2(new_n581_), .ZN(new_n815_));
  XOR2_X1   g614(.A(KEYINPUT61), .B(G155gat), .Z(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(G1346gat));
  OAI21_X1  g616(.A(G162gat), .B1(new_n809_), .B2(new_n628_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n616_), .A2(G162gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n809_), .B2(new_n819_), .ZN(G1347gat));
  NAND2_X1  g619(.A1(new_n782_), .A2(new_n763_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n642_), .A2(new_n403_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n765_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n824_), .A2(new_n513_), .A3(new_n354_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n824_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n214_), .B1(new_n826_), .B2(new_n665_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n827_), .B2(KEYINPUT62), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(KEYINPUT62), .B2(new_n827_), .ZN(G1348gat));
  NAND2_X1  g628(.A1(new_n822_), .A2(new_n329_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n830_), .A2(new_n215_), .A3(new_n664_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n808_), .A2(new_n417_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n215_), .B1(new_n824_), .B2(new_n664_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n833_), .A2(KEYINPUT124), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(KEYINPUT124), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n832_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT125), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT125), .B(new_n832_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1349gat));
  NOR3_X1   g639(.A1(new_n824_), .A2(new_n579_), .A3(new_n350_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n830_), .A2(new_n581_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n808_), .A2(new_n417_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n843_), .B2(new_n207_), .ZN(G1350gat));
  OAI21_X1  g643(.A(G190gat), .B1(new_n824_), .B2(new_n628_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n560_), .A2(new_n206_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n824_), .B2(new_n846_), .ZN(G1351gat));
  NAND4_X1  g646(.A1(new_n808_), .A2(new_n611_), .A3(new_n262_), .A4(new_n822_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n513_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT126), .B(G197gat), .Z(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1352gat));
  INV_X1    g650(.A(KEYINPUT127), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n479_), .B1(new_n852_), .B2(new_n296_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n848_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1353gat));
  NOR2_X1   g655(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n857_));
  AND2_X1   g656(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n858_));
  NOR4_X1   g657(.A1(new_n848_), .A2(new_n579_), .A3(new_n857_), .A4(new_n858_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n848_), .A2(new_n579_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n857_), .ZN(G1354gat));
  OAI21_X1  g660(.A(G218gat), .B1(new_n848_), .B2(new_n628_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n616_), .A2(G218gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n848_), .B2(new_n863_), .ZN(G1355gat));
endmodule


