//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(KEYINPUT92), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT92), .ZN(new_n211_));
  OAI22_X1  g010(.A1(new_n211_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n203_), .B(new_n204_), .C1(new_n207_), .C2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n203_), .A2(KEYINPUT1), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G155gat), .A3(G162gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n217_), .A3(new_n204_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G141gat), .B(G148gat), .Z(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT91), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT91), .B1(new_n218_), .B2(new_n219_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n214_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G127gat), .B(G134gat), .Z(new_n224_));
  XOR2_X1   g023(.A(G113gat), .B(G120gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n218_), .A2(new_n219_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT91), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n220_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(new_n226_), .A3(new_n214_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n228_), .A2(new_n233_), .A3(KEYINPUT4), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n223_), .A2(new_n227_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n202_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n228_), .A2(new_n233_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n239_), .A2(new_n202_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G1gat), .B(G29gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT101), .B(G85gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT0), .B(G57gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n238_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n246_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G78gat), .B(G106gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G228gat), .A2(G233gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n255_));
  NAND3_X1  g054(.A1(new_n223_), .A2(KEYINPUT96), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT21), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(G197gat), .A2(G204gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G197gat), .A2(G204gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT21), .A3(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n262_), .A2(new_n263_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT97), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT97), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n256_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT96), .B1(new_n223_), .B2(new_n255_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n254_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n223_), .A2(KEYINPUT29), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT94), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n253_), .A4(new_n266_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT29), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n232_), .B2(new_n214_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n266_), .A2(new_n253_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT94), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n252_), .B1(new_n273_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT98), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n273_), .A2(new_n281_), .A3(new_n252_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n232_), .A2(new_n277_), .A3(new_n214_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT28), .ZN(new_n288_));
  XOR2_X1   g087(.A(G22gat), .B(G50gat), .Z(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  AND3_X1   g089(.A1(new_n273_), .A2(new_n281_), .A3(new_n252_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT93), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n291_), .A2(new_n282_), .A3(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n286_), .B(new_n290_), .C1(new_n293_), .C2(new_n284_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295_));
  XOR2_X1   g094(.A(G8gat), .B(G36gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT18), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G226gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT19), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT23), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT22), .B(G169gat), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n312_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT85), .ZN(new_n317_));
  INV_X1    g116(.A(G169gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(new_n314_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT26), .B(G190gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT25), .B(G183gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n319_), .A2(KEYINPUT24), .A3(new_n312_), .A4(new_n320_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n323_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT88), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT88), .B1(new_n304_), .B2(KEYINPUT23), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n316_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n333_), .A2(KEYINPUT99), .A3(new_n266_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT99), .B1(new_n333_), .B2(new_n266_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(KEYINPUT83), .B(G183gat), .Z(new_n337_));
  OAI22_X1  g136(.A1(new_n330_), .A2(new_n331_), .B1(new_n337_), .B2(G190gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n318_), .A2(KEYINPUT86), .A3(KEYINPUT22), .ZN(new_n339_));
  AND2_X1   g138(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n339_), .B(new_n314_), .C1(new_n318_), .C2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT87), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n341_), .A2(new_n342_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n338_), .B(new_n312_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n266_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT25), .ZN(new_n347_));
  INV_X1    g146(.A(G183gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(KEYINPUT84), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT83), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(G183gat), .ZN(new_n351_));
  NOR4_X1   g150(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT83), .A4(KEYINPUT84), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n324_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n353_), .A2(new_n308_), .A3(new_n323_), .A4(new_n327_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n345_), .A2(new_n346_), .A3(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n355_), .A2(KEYINPUT20), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n303_), .B1(new_n336_), .B2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT20), .B(new_n303_), .C1(new_n333_), .C2(new_n266_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n346_), .B1(new_n345_), .B2(new_n354_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n300_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n333_), .A2(new_n266_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT99), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n333_), .A2(KEYINPUT99), .A3(new_n266_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n364_), .A2(KEYINPUT20), .A3(new_n355_), .A4(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n360_), .B1(new_n366_), .B2(new_n302_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n299_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n361_), .A2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT20), .B1(new_n270_), .B2(new_n333_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n359_), .B1(new_n370_), .B2(KEYINPUT105), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT20), .ZN(new_n372_));
  INV_X1    g171(.A(new_n269_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n268_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n333_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n372_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT105), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n303_), .B1(new_n371_), .B2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n366_), .A2(new_n302_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n300_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n295_), .B1(new_n367_), .B2(new_n299_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n295_), .A2(new_n369_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n283_), .A2(KEYINPUT93), .A3(new_n285_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n290_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(KEYINPUT98), .ZN(new_n387_));
  AND4_X1   g186(.A1(new_n251_), .A2(new_n294_), .A3(new_n384_), .A4(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n249_), .A2(KEYINPUT33), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT33), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n390_), .B(new_n248_), .C1(new_n237_), .C2(new_n240_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n234_), .A2(new_n202_), .A3(new_n236_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n392_), .A2(KEYINPUT102), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n246_), .B1(new_n239_), .B2(new_n202_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n392_), .B2(KEYINPUT102), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n389_), .A2(new_n391_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT100), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n361_), .A2(new_n368_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n361_), .B2(new_n368_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n396_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT103), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n396_), .B(KEYINPUT103), .C1(new_n398_), .C2(new_n399_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n380_), .A2(new_n381_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n299_), .A2(KEYINPUT32), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(KEYINPUT104), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n367_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n250_), .A2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n402_), .A2(new_n403_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n294_), .A2(new_n387_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n388_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n345_), .A2(new_n354_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416_));
  INV_X1    g215(.A(G71gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G99gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n415_), .B(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G15gat), .B(G43gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT89), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT30), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(new_n227_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n426_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT106), .B1(new_n414_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT106), .ZN(new_n431_));
  INV_X1    g230(.A(new_n429_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n413_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n410_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n403_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n431_), .B(new_n432_), .C1(new_n435_), .C2(new_n388_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n384_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(new_n429_), .A3(new_n251_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n430_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT69), .ZN(new_n441_));
  INV_X1    g240(.A(G230gat), .ZN(new_n442_));
  INV_X1    g241(.A(G233gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G57gat), .B(G64gat), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n446_), .A2(KEYINPUT11), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(KEYINPUT11), .ZN(new_n448_));
  XOR2_X1   g247(.A(G71gat), .B(G78gat), .Z(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n448_), .A2(new_n449_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT7), .ZN(new_n454_));
  INV_X1    g253(.A(G99gat), .ZN(new_n455_));
  INV_X1    g254(.A(G106gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n457_), .A2(new_n460_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G85gat), .A2(G92gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT8), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT8), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n463_), .A2(new_n471_), .A3(new_n468_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT64), .B(G106gat), .ZN(new_n474_));
  OR2_X1    g273(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n467_), .A2(KEYINPUT9), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n460_), .A2(new_n461_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n466_), .A2(KEYINPUT9), .A3(new_n467_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT65), .B1(new_n473_), .B2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n463_), .A2(new_n471_), .A3(new_n468_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n471_), .B1(new_n463_), .B2(new_n468_), .ZN(new_n484_));
  OAI211_X1 g283(.A(KEYINPUT65), .B(new_n481_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n453_), .B1(new_n482_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n481_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT65), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n452_), .A3(new_n485_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n445_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT66), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n453_), .A2(KEYINPUT12), .A3(new_n488_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n452_), .B1(new_n490_), .B2(new_n485_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(KEYINPUT12), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n445_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n498_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n487_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n500_), .A2(new_n502_), .A3(KEYINPUT67), .A4(new_n495_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n493_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G120gat), .B(G148gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G176gat), .B(G204gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n493_), .A2(new_n499_), .A3(new_n503_), .A4(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(KEYINPUT13), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT13), .B1(new_n510_), .B2(new_n512_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n441_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT69), .A3(new_n513_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G169gat), .B(G197gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G1gat), .B(G8gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT76), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(G15gat), .A2(G22gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G15gat), .A2(G22gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G1gat), .A2(G8gat), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n530_), .A2(new_n531_), .B1(KEYINPUT14), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n529_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G29gat), .B(G36gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G43gat), .B(G50gat), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n536_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n534_), .B(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n537_), .A2(KEYINPUT15), .A3(new_n538_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT15), .B1(new_n537_), .B2(new_n538_), .ZN(new_n545_));
  OR3_X1    g344(.A1(new_n534_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n534_), .A2(new_n539_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n541_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n526_), .B1(new_n543_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n543_), .A2(new_n548_), .A3(new_n526_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(KEYINPUT81), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT81), .ZN(new_n553_));
  INV_X1    g352(.A(new_n551_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(new_n549_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT82), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(new_n555_), .A3(KEYINPUT82), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n520_), .A2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n440_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n452_), .B(new_n562_), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(new_n534_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT78), .ZN(new_n566_));
  XOR2_X1   g365(.A(G183gat), .B(G211gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n570_), .A2(new_n571_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n564_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n573_), .A2(new_n564_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT37), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT72), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT34), .Z(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n544_), .A2(new_n545_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n488_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n490_), .A2(new_n539_), .A3(new_n485_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n581_), .A2(new_n582_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT71), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n587_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(KEYINPUT71), .A3(new_n589_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n584_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n583_), .B1(new_n585_), .B2(new_n488_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n588_), .A2(new_n595_), .A3(new_n589_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(KEYINPUT36), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n579_), .B1(new_n594_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n601_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n588_), .A2(KEYINPUT71), .A3(new_n589_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT71), .B1(new_n588_), .B2(new_n589_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n587_), .ZN(new_n606_));
  OAI211_X1 g405(.A(KEYINPUT72), .B(new_n603_), .C1(new_n606_), .C2(new_n584_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n599_), .B(KEYINPUT36), .Z(new_n609_));
  INV_X1    g408(.A(new_n596_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n609_), .B1(new_n594_), .B2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n578_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n590_), .A2(new_n591_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n593_), .A3(new_n586_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n583_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT72), .B1(new_n616_), .B2(new_n603_), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n579_), .B(new_n601_), .C1(new_n615_), .C2(new_n583_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n578_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n609_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT73), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n594_), .B2(new_n610_), .ZN(new_n622_));
  OAI211_X1 g421(.A(KEYINPUT73), .B(new_n596_), .C1(new_n606_), .C2(new_n584_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n620_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n619_), .A2(new_n624_), .A3(KEYINPUT74), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT74), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT73), .B1(new_n616_), .B2(new_n596_), .ZN(new_n627_));
  AOI211_X1 g426(.A(new_n621_), .B(new_n610_), .C1(new_n615_), .C2(new_n583_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n609_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT37), .B1(new_n602_), .B2(new_n607_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n613_), .B1(new_n625_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT75), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT74), .B1(new_n619_), .B2(new_n624_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n629_), .A2(new_n626_), .A3(new_n630_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(KEYINPUT75), .A3(new_n613_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n577_), .B1(new_n634_), .B2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n561_), .A2(new_n639_), .ZN(new_n640_));
  OR3_X1    g439(.A1(new_n640_), .A2(G1gat), .A3(new_n251_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT38), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n629_), .A2(new_n608_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n440_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n552_), .A2(new_n555_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n520_), .A2(new_n577_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n251_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n641_), .A2(new_n642_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n643_), .A2(new_n650_), .A3(new_n651_), .ZN(G1324gat));
  NAND3_X1  g451(.A1(new_n645_), .A2(new_n437_), .A3(new_n648_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G8gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT39), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n384_), .A2(G8gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n561_), .A2(new_n639_), .A3(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT107), .Z(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n655_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  OAI21_X1  g461(.A(G15gat), .B1(new_n649_), .B2(new_n432_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n640_), .A2(G15gat), .A3(new_n432_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1326gat));
  OAI21_X1  g465(.A(G22gat), .B1(new_n649_), .B2(new_n413_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT42), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n413_), .A2(G22gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n640_), .B2(new_n669_), .ZN(G1327gat));
  NOR2_X1   g469(.A1(new_n644_), .A2(new_n576_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n561_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G29gat), .B1(new_n673_), .B2(new_n250_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n520_), .A2(new_n576_), .A3(new_n647_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT75), .B1(new_n637_), .B2(new_n613_), .ZN(new_n677_));
  AOI211_X1 g476(.A(new_n633_), .B(new_n612_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT109), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n634_), .A2(new_n680_), .A3(new_n638_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n676_), .B1(new_n682_), .B2(new_n440_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n634_), .A2(new_n638_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(KEYINPUT43), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(new_n440_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n675_), .C1(new_n683_), .C2(new_n686_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n687_), .A2(G29gat), .A3(new_n250_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n440_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n690_));
  AOI22_X1  g489(.A1(new_n690_), .A2(KEYINPUT43), .B1(new_n440_), .B2(new_n685_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n675_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n674_), .B1(new_n688_), .B2(new_n693_), .ZN(G1328gat));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n695_));
  INV_X1    g494(.A(G36gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n691_), .A2(new_n692_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n384_), .B1(new_n697_), .B2(KEYINPUT44), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n698_), .B2(new_n693_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n561_), .A2(new_n696_), .A3(new_n437_), .A4(new_n671_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n695_), .B1(new_n699_), .B2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n693_), .A2(new_n687_), .A3(new_n437_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(G36gat), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1329gat));
  NAND4_X1  g506(.A1(new_n693_), .A2(new_n687_), .A3(G43gat), .A4(new_n429_), .ZN(new_n708_));
  INV_X1    g507(.A(G43gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n672_), .B2(new_n432_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g511(.A(G50gat), .B1(new_n673_), .B2(new_n433_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n687_), .A2(G50gat), .A3(new_n433_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(new_n693_), .ZN(G1331gat));
  NAND3_X1  g514(.A1(new_n557_), .A2(new_n576_), .A3(new_n558_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n519_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n645_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n251_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n440_), .A2(new_n520_), .A3(new_n647_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(new_n639_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n251_), .A2(G57gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n721_), .A2(new_n725_), .A3(new_n437_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n718_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n437_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(G64gat), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G64gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n726_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT111), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n726_), .B(new_n734_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1333gat));
  NAND3_X1  g535(.A1(new_n721_), .A2(new_n417_), .A3(new_n429_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT49), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n727_), .A2(new_n429_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G71gat), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT49), .B(new_n417_), .C1(new_n727_), .C2(new_n429_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT112), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(new_n737_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1334gat));
  OAI21_X1  g545(.A(G78gat), .B1(new_n718_), .B2(new_n413_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT50), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n413_), .A2(G78gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n722_), .B2(new_n749_), .ZN(G1335gat));
  NOR3_X1   g549(.A1(new_n519_), .A2(new_n576_), .A3(new_n646_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n751_), .B1(new_n683_), .B2(new_n686_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n251_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n720_), .A2(new_n671_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n464_), .A3(new_n250_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1336gat));
  OAI21_X1  g555(.A(G92gat), .B1(new_n752_), .B2(new_n384_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n754_), .A2(new_n465_), .A3(new_n437_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n752_), .B2(new_n432_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n754_), .A2(new_n475_), .A3(new_n476_), .A4(new_n429_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n754_), .A2(new_n474_), .A3(new_n433_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n433_), .B(new_n751_), .C1(new_n683_), .C2(new_n686_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(G106gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G106gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT53), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n764_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1339gat));
  NAND2_X1  g572(.A1(new_n540_), .A2(new_n541_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT119), .B1(new_n774_), .B2(new_n525_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n546_), .A2(new_n547_), .A3(new_n542_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(KEYINPUT119), .A3(new_n525_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n554_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n512_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n503_), .A2(new_n499_), .A3(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n497_), .A2(new_n498_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT55), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n502_), .A2(new_n495_), .A3(new_n491_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n444_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n509_), .B1(new_n782_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT56), .B(new_n509_), .C1(new_n782_), .C2(new_n787_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n780_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT58), .B1(new_n792_), .B2(KEYINPUT120), .ZN(new_n793_));
  INV_X1    g592(.A(new_n792_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n634_), .A2(new_n638_), .A3(new_n793_), .A4(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n646_), .A2(new_n512_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT116), .B(new_n509_), .C1(new_n782_), .C2(new_n787_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(KEYINPUT55), .A2(new_n783_), .B1(new_n785_), .B2(new_n444_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n503_), .A2(new_n499_), .A3(new_n781_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n511_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(KEYINPUT116), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n802_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n791_), .A2(KEYINPUT118), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(new_n809_), .A3(KEYINPUT56), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n799_), .B1(new_n807_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n510_), .A2(new_n512_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n813_), .A2(new_n779_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT57), .B(new_n644_), .C1(new_n812_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n808_), .B(new_n810_), .C1(new_n802_), .C2(new_n806_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n799_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n814_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n644_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n798_), .A2(new_n815_), .A3(new_n821_), .A4(KEYINPUT121), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n798_), .A2(new_n815_), .A3(new_n821_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n576_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n716_), .A2(new_n515_), .A3(new_n514_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n826_), .B(new_n827_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT114), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n684_), .A2(new_n830_), .A3(new_n826_), .A4(new_n827_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n559_), .A2(new_n517_), .A3(new_n576_), .A4(new_n513_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n634_), .B2(new_n638_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n835_), .B2(new_n826_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n827_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n826_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(KEYINPUT115), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n822_), .A2(new_n825_), .B1(new_n832_), .B2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n432_), .A2(new_n251_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n438_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(KEYINPUT59), .ZN(new_n845_));
  INV_X1    g644(.A(new_n815_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n798_), .A2(new_n821_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n798_), .A2(new_n821_), .A3(KEYINPUT122), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n576_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n829_), .A2(new_n831_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n845_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n844_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n559_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n841_), .A2(new_n843_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n647_), .A2(G113gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n858_), .B2(new_n859_), .ZN(G1340gat));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n847_), .A2(new_n848_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(new_n815_), .A3(new_n850_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n863_), .A2(new_n577_), .B1(new_n832_), .B2(new_n840_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n845_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n520_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n823_), .A2(new_n824_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n868_), .A2(new_n577_), .A3(new_n822_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n835_), .A2(new_n833_), .A3(new_n826_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT115), .B1(new_n837_), .B2(new_n838_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n829_), .B(new_n831_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n869_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n843_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n867_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n861_), .B1(new_n866_), .B2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n844_), .A2(KEYINPUT123), .A3(new_n520_), .A4(new_n854_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(G120gat), .ZN(new_n878_));
  INV_X1    g677(.A(G120gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n519_), .B2(KEYINPUT60), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n857_), .B(new_n880_), .C1(KEYINPUT60), .C2(new_n879_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(G1341gat));
  OAI21_X1  g681(.A(G127gat), .B1(new_n855_), .B2(new_n577_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n577_), .A2(G127gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n858_), .B2(new_n884_), .ZN(G1342gat));
  OAI21_X1  g684(.A(G134gat), .B1(new_n855_), .B2(new_n684_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n644_), .A2(G134gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n858_), .B2(new_n887_), .ZN(G1343gat));
  NAND4_X1  g687(.A1(new_n433_), .A2(new_n432_), .A3(new_n250_), .A4(new_n384_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT124), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n873_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n647_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n519_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT125), .B(G148gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1345gat));
  OAI21_X1  g695(.A(KEYINPUT126), .B1(new_n891_), .B2(new_n577_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT126), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n873_), .A2(new_n898_), .A3(new_n576_), .A4(new_n890_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n897_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n897_), .B2(new_n899_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1346gat));
  INV_X1    g702(.A(G162gat), .ZN(new_n904_));
  INV_X1    g703(.A(new_n682_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n891_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n873_), .A2(new_n820_), .A3(new_n890_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n904_), .B2(new_n907_), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n384_), .A2(new_n250_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n432_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n413_), .B(new_n912_), .C1(new_n851_), .C2(new_n853_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n647_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n909_), .B1(new_n914_), .B2(new_n318_), .ZN(new_n915_));
  OAI211_X1 g714(.A(KEYINPUT62), .B(G169gat), .C1(new_n913_), .C2(new_n647_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n313_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(G1348gat));
  INV_X1    g717(.A(new_n913_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G176gat), .B1(new_n919_), .B2(new_n520_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n841_), .A2(new_n433_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n912_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n519_), .A2(new_n314_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n920_), .B1(new_n921_), .B2(new_n923_), .ZN(G1349gat));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n577_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n337_), .B1(new_n921_), .B2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n864_), .A2(new_n433_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n922_), .A2(new_n577_), .A3(new_n325_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n913_), .B2(new_n684_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n820_), .A2(new_n324_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n913_), .B2(new_n931_), .ZN(G1351gat));
  NAND3_X1  g731(.A1(new_n433_), .A2(new_n432_), .A3(new_n910_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n841_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n646_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g735(.A1(new_n841_), .A2(new_n519_), .A3(new_n933_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  XOR2_X1   g738(.A(KEYINPUT127), .B(G204gat), .Z(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n937_), .B2(new_n940_), .ZN(G1353gat));
  NAND2_X1  g740(.A1(new_n934_), .A2(new_n576_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  AND2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n942_), .A2(new_n943_), .A3(new_n944_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n942_), .A2(new_n943_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1354gat));
  INV_X1    g746(.A(G218gat), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n934_), .A2(new_n948_), .A3(new_n820_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n841_), .A2(new_n684_), .A3(new_n933_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n948_), .ZN(G1355gat));
endmodule


