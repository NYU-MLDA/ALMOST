//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT78), .B(G1gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n208_), .A2(G8gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n207_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n206_), .A2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(new_n204_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT80), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(KEYINPUT81), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n213_), .B(new_n204_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G229gat), .A3(G233gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT81), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n216_), .A2(new_n218_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G141gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G169gat), .B(G197gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n226_), .B(new_n227_), .Z(new_n228_));
  OR2_X1    g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n228_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G71gat), .B(G78gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(G57gat), .B(G64gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n234_), .B1(KEYINPUT11), .B2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT68), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n235_), .A2(KEYINPUT11), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240_));
  INV_X1    g039(.A(G99gat), .ZN(new_n241_));
  INV_X1    g040(.A(G106gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT7), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G99gat), .A2(G106gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT6), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n249_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n252_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n248_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G85gat), .B(G92gat), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n248_), .A2(new_n251_), .A3(new_n249_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n257_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT8), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n258_), .A2(KEYINPUT8), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(KEYINPUT9), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT10), .B(G99gat), .Z(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n242_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT64), .B(G92gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT9), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(G85gat), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n263_), .A2(new_n265_), .A3(new_n251_), .A4(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n239_), .B1(new_n262_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n259_), .A2(new_n261_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n253_), .B1(new_n252_), .B2(new_n251_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n260_), .B1(new_n275_), .B2(new_n248_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT8), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n274_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n237_), .B(new_n238_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n269_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n239_), .A2(KEYINPUT12), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n269_), .B(KEYINPUT70), .Z(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n262_), .A2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n280_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G230gat), .A2(G233gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OR3_X1    g086(.A1(new_n273_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n271_), .A2(new_n289_), .A3(new_n280_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n290_), .B(new_n287_), .C1(new_n289_), .C2(new_n280_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G120gat), .B(G148gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(G176gat), .B(G204gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n292_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n292_), .A2(new_n298_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n233_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n292_), .A2(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n292_), .A2(new_n298_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n301_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n231_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT99), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n301_), .A2(new_n305_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT73), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n301_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT99), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n231_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G8gat), .B(G36gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT18), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G64gat), .B(G92gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT19), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT95), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT21), .ZN(new_n326_));
  AND2_X1   g125(.A1(G197gat), .A2(G204gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G197gat), .A2(G204gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G197gat), .ZN(new_n330_));
  INV_X1    g129(.A(G204gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G197gat), .A2(G204gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT21), .A3(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n329_), .A2(new_n334_), .A3(KEYINPUT88), .A4(new_n335_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n329_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n336_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n342_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT25), .B(G183gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT26), .B(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT23), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(G183gat), .A3(G190gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT84), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT84), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n350_), .B2(KEYINPUT23), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n346_), .B(new_n349_), .C1(new_n354_), .C2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT22), .ZN(new_n358_));
  INV_X1    g157(.A(G169gat), .ZN(new_n359_));
  INV_X1    g158(.A(G176gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT92), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n351_), .A2(new_n353_), .ZN(new_n365_));
  INV_X1    g164(.A(G183gat), .ZN(new_n366_));
  INV_X1    g165(.A(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT92), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n361_), .A2(new_n370_), .A3(new_n362_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n364_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n357_), .A2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT20), .B1(new_n341_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT89), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n375_), .B(new_n336_), .C1(new_n337_), .C2(new_n339_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n329_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n378_));
  INV_X1    g177(.A(G218gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G211gat), .ZN(new_n380_));
  INV_X1    g179(.A(G211gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G218gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n327_), .A2(new_n328_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(KEYINPUT21), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n378_), .A2(new_n338_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n375_), .B1(new_n386_), .B2(new_n336_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n377_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n366_), .A2(KEYINPUT25), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(G183gat), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT82), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n366_), .B2(KEYINPUT25), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n392_), .A2(KEYINPUT83), .A3(new_n394_), .A4(new_n348_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n367_), .A2(KEYINPUT26), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT26), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G190gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n394_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n390_), .A2(G183gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n366_), .A2(KEYINPUT25), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n393_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n396_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n395_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n346_), .A2(new_n365_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n368_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n363_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n405_), .A2(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n325_), .A2(new_n374_), .B1(new_n388_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n357_), .A2(new_n372_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(new_n340_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT95), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n324_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n410_), .B1(new_n377_), .B2(new_n387_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n413_), .B1(new_n341_), .B2(new_n373_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n418_), .A2(new_n324_), .A3(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n321_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n340_), .A2(KEYINPUT89), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n408_), .A2(new_n409_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n406_), .B1(new_n395_), .B2(new_n404_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n422_), .B(new_n376_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n324_), .A3(new_n415_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n340_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n376_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(new_n410_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n320_), .B(new_n426_), .C1(new_n429_), .C2(new_n324_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n430_), .A2(KEYINPUT27), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n421_), .A2(new_n431_), .A3(KEYINPUT98), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n374_), .A2(new_n325_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(new_n416_), .A3(new_n425_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n323_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n420_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n320_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n430_), .A2(KEYINPUT27), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n433_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n426_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n324_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n321_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n430_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT27), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n432_), .A2(new_n440_), .A3(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G22gat), .B(G50gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G155gat), .A2(G162gat), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(KEYINPUT1), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G155gat), .A2(G162gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n451_), .B2(KEYINPUT1), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT85), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n450_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT1), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n455_), .B1(G155gat), .B2(G162gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(KEYINPUT85), .A3(new_n449_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G141gat), .A2(G148gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G141gat), .A2(G148gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT29), .ZN(new_n464_));
  INV_X1    g263(.A(new_n449_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n465_), .A2(new_n451_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT3), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n461_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT2), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n459_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n466_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n463_), .A2(new_n464_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT28), .ZN(new_n478_));
  INV_X1    g277(.A(new_n462_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n466_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n471_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n467_), .B(KEYINPUT86), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT28), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n464_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n448_), .B1(new_n478_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n478_), .A2(new_n487_), .A3(new_n448_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT91), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n492_));
  INV_X1    g291(.A(new_n490_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n488_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G78gat), .B(G106gat), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G233gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(G228gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(G228gat), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n497_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n464_), .B1(new_n463_), .B2(new_n476_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n341_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n504_), .B(KEYINPUT29), .C1(new_n480_), .C2(new_n484_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n502_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n502_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT29), .B1(new_n480_), .B2(new_n484_), .ZN(new_n510_));
  AND4_X1   g309(.A1(new_n509_), .A2(new_n422_), .A3(new_n510_), .A4(new_n376_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n496_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n340_), .B1(new_n510_), .B2(KEYINPUT90), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n509_), .B1(new_n514_), .B2(new_n506_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n515_), .A2(new_n511_), .A3(new_n495_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n491_), .B(new_n494_), .C1(new_n513_), .C2(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n493_), .A2(new_n488_), .A3(new_n492_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n508_), .A2(new_n512_), .A3(new_n496_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n495_), .B1(new_n515_), .B2(new_n511_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n447_), .A2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G71gat), .B(G99gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G43gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n410_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G127gat), .B(G134gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G113gat), .B(G120gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n526_), .B(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G227gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(G15gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT30), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT31), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(new_n536_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G1gat), .B(G29gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(G85gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT0), .B(G57gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  XOR2_X1   g343(.A(new_n527_), .B(new_n528_), .Z(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n456_), .A2(KEYINPUT85), .A3(new_n449_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT85), .B1(new_n456_), .B2(new_n449_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n450_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n476_), .B(new_n529_), .C1(new_n549_), .C2(new_n479_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n546_), .A2(new_n550_), .A3(KEYINPUT4), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT93), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT93), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n546_), .A2(new_n550_), .A3(new_n553_), .A4(KEYINPUT4), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G225gat), .A2(G233gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT94), .Z(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n546_), .B2(KEYINPUT4), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n546_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n550_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n557_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n544_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n558_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n544_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n566_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT97), .B1(new_n565_), .B2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n563_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n544_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT97), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n567_), .B1(new_n566_), .B2(new_n563_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n540_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n523_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT4), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n557_), .B1(new_n561_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n555_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n561_), .A2(new_n562_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n544_), .B1(new_n581_), .B2(new_n557_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n443_), .A3(new_n430_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT33), .B1(new_n570_), .B2(new_n544_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT33), .ZN(new_n586_));
  NOR4_X1   g385(.A1(new_n566_), .A2(new_n586_), .A3(new_n563_), .A4(new_n567_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n584_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n565_), .A2(new_n568_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n320_), .A2(KEYINPUT32), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n426_), .B(new_n590_), .C1(new_n429_), .C2(new_n324_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n420_), .B1(new_n323_), .B2(new_n435_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n591_), .B1(new_n592_), .B2(new_n590_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n522_), .B1(new_n588_), .B2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n522_), .B1(new_n569_), .B2(new_n574_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n595_), .A2(KEYINPUT96), .B1(new_n447_), .B2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n517_), .A2(new_n521_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n585_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n443_), .A2(new_n430_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n587_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .A4(new_n583_), .ZN(new_n602_));
  OAI221_X1 g401(.A(new_n591_), .B1(new_n592_), .B2(new_n590_), .C1(new_n565_), .C2(new_n568_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n598_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n597_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n577_), .B1(new_n607_), .B2(new_n539_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT34), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n262_), .A2(new_n204_), .A3(new_n270_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n205_), .B1(new_n278_), .B2(new_n282_), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT35), .B(new_n610_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n206_), .B1(new_n262_), .B2(new_n283_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n204_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n278_), .A2(new_n615_), .A3(new_n269_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n610_), .A2(KEYINPUT35), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n610_), .A2(KEYINPUT35), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n614_), .A2(new_n616_), .A3(new_n617_), .A4(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT36), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n623_), .A2(KEYINPUT36), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n613_), .A2(new_n626_), .A3(new_n619_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT100), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n608_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n279_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(new_n213_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G127gat), .B(G155gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G183gat), .B(G211gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT17), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n640_), .A2(new_n641_), .ZN(new_n643_));
  OR3_X1    g442(.A1(new_n635_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n635_), .A2(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n310_), .A2(new_n316_), .A3(new_n631_), .A4(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n575_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT101), .Z(new_n650_));
  INV_X1    g449(.A(KEYINPUT74), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n312_), .A2(KEYINPUT74), .A3(new_n313_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n231_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n608_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n624_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n613_), .B2(new_n619_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n627_), .B1(new_n658_), .B2(KEYINPUT75), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n620_), .A2(KEYINPUT75), .A3(new_n624_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT37), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT76), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT76), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n663_), .B(KEYINPUT37), .C1(new_n659_), .C2(new_n660_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT37), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n625_), .A2(new_n665_), .A3(new_n627_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT77), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT77), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n628_), .A2(new_n668_), .A3(new_n665_), .ZN(new_n669_));
  AOI22_X1  g468(.A1(new_n662_), .A2(new_n664_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n646_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n654_), .A2(new_n656_), .A3(new_n671_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n672_), .A2(new_n575_), .A3(new_n208_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT38), .Z(new_n674_));
  NAND2_X1  g473(.A1(new_n650_), .A2(new_n674_), .ZN(G1324gat));
  OAI21_X1  g474(.A(G8gat), .B1(new_n648_), .B2(new_n447_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT39), .ZN(new_n677_));
  OR3_X1    g476(.A1(new_n672_), .A2(G8gat), .A3(new_n447_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g479(.A1(new_n540_), .A2(new_n532_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n672_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G15gat), .B1(new_n648_), .B2(new_n539_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n685_));
  AOI21_X1  g484(.A(new_n682_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n684_), .B2(new_n685_), .ZN(G1326gat));
  OAI21_X1  g486(.A(G22gat), .B1(new_n648_), .B2(new_n522_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT42), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n522_), .A2(G22gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n672_), .B2(new_n690_), .ZN(G1327gat));
  NOR2_X1   g490(.A1(new_n647_), .A2(new_n629_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n314_), .A2(new_n656_), .A3(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT105), .ZN(new_n694_));
  INV_X1    g493(.A(new_n575_), .ZN(new_n695_));
  INV_X1    g494(.A(G29gat), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT106), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n310_), .A2(new_n316_), .A3(new_n646_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n310_), .A2(new_n316_), .A3(KEYINPUT103), .A4(new_n646_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n540_), .B1(new_n597_), .B2(new_n606_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n705_), .B(new_n670_), .C1(new_n706_), .C2(new_n577_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT104), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n575_), .A2(new_n598_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n432_), .A2(new_n440_), .A3(new_n446_), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n604_), .A2(new_n605_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n595_), .A2(KEYINPUT96), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n539_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n577_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n705_), .A4(new_n670_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n670_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n608_), .B2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n708_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n704_), .A2(KEYINPUT44), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT44), .B1(new_n704_), .B2(new_n720_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n722_), .A2(new_n575_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n699_), .B1(new_n724_), .B2(new_n696_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT107), .B(new_n699_), .C1(new_n724_), .C2(new_n696_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n693_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n693_), .A2(new_n730_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n447_), .A2(G36gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n735_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n694_), .B2(new_n733_), .ZN(new_n738_));
  OAI22_X1  g537(.A1(new_n736_), .A2(new_n738_), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n704_), .A2(new_n720_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n710_), .A3(new_n721_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n739_), .B1(new_n743_), .B2(G36gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT110), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n744_), .B(new_n746_), .ZN(G1329gat));
  NAND4_X1  g546(.A1(new_n742_), .A2(G43gat), .A3(new_n540_), .A4(new_n721_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n694_), .A2(new_n540_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(G43gat), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g550(.A1(new_n522_), .A2(G50gat), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT111), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n694_), .A2(new_n753_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n722_), .A2(new_n522_), .A3(new_n723_), .ZN(new_n755_));
  INV_X1    g554(.A(G50gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(G1331gat));
  INV_X1    g556(.A(new_n314_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n608_), .A2(new_n231_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n671_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(G57gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n695_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n231_), .A2(new_n646_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n652_), .A2(new_n653_), .A3(new_n631_), .A4(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G57gat), .B1(new_n764_), .B2(new_n575_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1332gat));
  INV_X1    g565(.A(G64gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n760_), .A2(new_n767_), .A3(new_n710_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n764_), .A2(new_n447_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(G64gat), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G64gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(G1333gat));
  INV_X1    g572(.A(G71gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n760_), .A2(new_n774_), .A3(new_n540_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G71gat), .B1(new_n764_), .B2(new_n539_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(KEYINPUT49), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(KEYINPUT49), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n777_), .B2(new_n778_), .ZN(G1334gat));
  NOR2_X1   g578(.A1(new_n522_), .A2(G78gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT113), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n760_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(G78gat), .B1(new_n764_), .B2(new_n522_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(KEYINPUT50), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT50), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n782_), .B1(new_n784_), .B2(new_n785_), .ZN(G1335gat));
  AND3_X1   g585(.A1(new_n652_), .A2(new_n653_), .A3(new_n692_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n759_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(G85gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n695_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n312_), .A2(new_n646_), .A3(new_n655_), .A4(new_n313_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n720_), .A2(KEYINPUT114), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n708_), .A2(new_n719_), .A3(new_n717_), .A4(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n792_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n796_), .A2(new_n695_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n791_), .B1(new_n797_), .B2(new_n790_), .ZN(G1336gat));
  AOI21_X1  g597(.A(G92gat), .B1(new_n789_), .B2(new_n710_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n710_), .A2(new_n266_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n796_), .B2(new_n800_), .ZN(G1337gat));
  AOI21_X1  g600(.A(new_n241_), .B1(new_n796_), .B2(new_n540_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n787_), .A2(new_n540_), .A3(new_n264_), .A4(new_n759_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT115), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n539_), .B(new_n792_), .C1(new_n793_), .C2(new_n795_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n806_), .B(new_n803_), .C1(new_n807_), .C2(new_n241_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(KEYINPUT51), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n796_), .A2(new_n540_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n804_), .B1(new_n811_), .B2(G99gat), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n810_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n809_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n805_), .A2(new_n810_), .A3(KEYINPUT51), .A4(new_n808_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1338gat));
  NOR2_X1   g619(.A1(new_n792_), .A2(new_n522_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n242_), .B1(new_n821_), .B2(new_n720_), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n822_), .B(KEYINPUT52), .Z(new_n823_));
  NAND2_X1  g622(.A1(new_n598_), .A2(new_n242_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n788_), .B2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n827_));
  INV_X1    g626(.A(G113gat), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n718_), .A2(new_n311_), .A3(new_n763_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n831_), .A2(KEYINPUT54), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(KEYINPUT54), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n273_), .A2(new_n285_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n287_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n288_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n837_), .A2(new_n836_), .A3(new_n287_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n298_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT120), .B1(new_n843_), .B2(KEYINPUT56), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n838_), .A2(new_n839_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n297_), .B1(new_n845_), .B2(new_n841_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n844_), .A2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT56), .B(new_n297_), .C1(new_n845_), .C2(new_n841_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n228_), .B1(new_n220_), .B2(new_n218_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n216_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n218_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n230_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n852_), .A2(KEYINPUT58), .A3(new_n303_), .A4(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n844_), .A2(new_n849_), .B1(KEYINPUT56), .B2(new_n843_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n303_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n861_), .A3(new_n670_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n851_), .A2(KEYINPUT119), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n655_), .A2(new_n299_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n843_), .A2(KEYINPUT56), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n851_), .A2(KEYINPUT119), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n863_), .B(new_n864_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n856_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n629_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(KEYINPUT57), .A3(new_n629_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n862_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n835_), .B1(new_n874_), .B2(new_n646_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n523_), .A2(new_n575_), .A3(new_n539_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n829_), .B1(new_n875_), .B2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n869_), .B2(new_n629_), .ZN(new_n879_));
  AOI211_X1 g678(.A(new_n871_), .B(new_n630_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n647_), .B1(new_n881_), .B2(new_n862_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT59), .B(new_n876_), .C1(new_n882_), .C2(new_n835_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n878_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n828_), .B1(new_n884_), .B2(new_n231_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n875_), .A2(new_n877_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n231_), .A2(new_n828_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n827_), .B1(new_n885_), .B2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n655_), .B1(new_n878_), .B2(new_n883_), .ZN(new_n891_));
  OAI221_X1 g690(.A(KEYINPUT121), .B1(new_n887_), .B2(new_n888_), .C1(new_n891_), .C2(new_n828_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1340gat));
  NOR2_X1   g692(.A1(new_n314_), .A2(KEYINPUT60), .ZN(new_n894_));
  MUX2_X1   g693(.A(new_n894_), .B(KEYINPUT60), .S(G120gat), .Z(new_n895_));
  NAND2_X1  g694(.A1(new_n886_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n654_), .B1(new_n878_), .B2(new_n883_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G120gat), .B1(new_n897_), .B2(new_n898_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n896_), .B1(new_n899_), .B2(new_n900_), .ZN(G1341gat));
  AOI21_X1  g700(.A(G127gat), .B1(new_n886_), .B2(new_n647_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n902_), .A2(KEYINPUT123), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(KEYINPUT123), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n647_), .A2(G127gat), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n903_), .A2(new_n904_), .B1(new_n884_), .B2(new_n905_), .ZN(G1342gat));
  INV_X1    g705(.A(G134gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n886_), .A2(new_n907_), .A3(new_n630_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n718_), .B1(new_n878_), .B2(new_n883_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n907_), .ZN(G1343gat));
  INV_X1    g709(.A(new_n875_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n540_), .A2(new_n522_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n911_), .A2(new_n695_), .A3(new_n447_), .A4(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n655_), .ZN(new_n914_));
  INV_X1    g713(.A(G141gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1344gat));
  NOR2_X1   g715(.A1(new_n913_), .A2(new_n654_), .ZN(new_n917_));
  INV_X1    g716(.A(G148gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1345gat));
  NOR2_X1   g718(.A1(new_n913_), .A2(new_n646_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT61), .B(G155gat), .Z(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1346gat));
  INV_X1    g721(.A(G162gat), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n913_), .A2(new_n923_), .A3(new_n718_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n913_), .B2(new_n629_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(KEYINPUT124), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n927_), .B(new_n923_), .C1(new_n913_), .C2(new_n629_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n924_), .B1(new_n926_), .B2(new_n928_), .ZN(G1347gat));
  NOR3_X1   g728(.A1(new_n576_), .A2(new_n447_), .A3(new_n598_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n875_), .A2(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(KEYINPUT22), .B(G169gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n932_), .A2(new_n231_), .A3(new_n933_), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n231_), .B(new_n930_), .C1(new_n882_), .C2(new_n835_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n359_), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n934_), .B1(new_n938_), .B2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  OAI211_X1 g741(.A(KEYINPUT126), .B(new_n934_), .C1(new_n938_), .C2(new_n939_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1348gat));
  INV_X1    g743(.A(new_n932_), .ZN(new_n945_));
  OAI21_X1  g744(.A(G176gat), .B1(new_n945_), .B2(new_n654_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n932_), .A2(new_n360_), .A3(new_n758_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1349gat));
  AOI21_X1  g747(.A(G183gat), .B1(new_n932_), .B2(new_n647_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n949_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n932_), .A2(new_n647_), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n950_), .B(new_n951_), .C1(new_n347_), .C2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(new_n347_), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT127), .B1(new_n954_), .B2(new_n949_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n953_), .A2(new_n955_), .ZN(G1350gat));
  OAI21_X1  g755(.A(G190gat), .B1(new_n945_), .B2(new_n718_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n932_), .A2(new_n348_), .A3(new_n630_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1351gat));
  NAND4_X1  g758(.A1(new_n911_), .A2(new_n575_), .A3(new_n710_), .A4(new_n912_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n960_), .A2(new_n655_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(new_n330_), .ZN(G1352gat));
  NOR2_X1   g761(.A1(new_n960_), .A2(new_n654_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(new_n331_), .ZN(G1353gat));
  NOR2_X1   g763(.A1(new_n960_), .A2(new_n646_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  AND2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n968_), .B1(new_n965_), .B2(new_n966_), .ZN(G1354gat));
  OAI21_X1  g768(.A(G218gat), .B1(new_n960_), .B2(new_n718_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n630_), .A2(new_n379_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n970_), .B1(new_n960_), .B2(new_n971_), .ZN(G1355gat));
endmodule


