//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT92), .B1(G155gat), .B2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR3_X1   g005(.A1(KEYINPUT92), .A2(G155gat), .A3(G162gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n204_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT91), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT91), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .A4(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n202_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT95), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT93), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT94), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n211_), .B(new_n221_), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n218_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n214_), .B1(new_n216_), .B2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G127gat), .B(G134gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G120gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT99), .B1(new_n224_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n215_), .A2(KEYINPUT95), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n215_), .A2(KEYINPUT95), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n218_), .A2(new_n220_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n229_), .B(new_n230_), .C1(new_n231_), .C2(new_n222_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT99), .ZN(new_n233_));
  INV_X1    g032(.A(new_n227_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .A4(new_n214_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n225_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(new_n226_), .ZN(new_n237_));
  MUX2_X1   g036(.A(new_n237_), .B(new_n227_), .S(KEYINPUT89), .Z(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n224_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n228_), .A2(new_n235_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT4), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G225gat), .A2(G233gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT0), .B(G57gat), .ZN(new_n247_));
  INV_X1    g046(.A(G85gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G1gat), .B(G29gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n240_), .A2(new_n242_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n246_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n251_), .B1(new_n246_), .B2(new_n252_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G169gat), .ZN(new_n256_));
  INV_X1    g055(.A(G176gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT97), .Z(new_n260_));
  NAND2_X1  g059(.A1(G183gat), .A2(G190gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(KEYINPUT23), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT87), .B(KEYINPUT23), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(new_n261_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n258_), .B(new_n260_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(KEYINPUT23), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n267_), .B1(new_n263_), .B2(new_n261_), .ZN(new_n268_));
  INV_X1    g067(.A(G169gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n257_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(KEYINPUT24), .A3(new_n259_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(KEYINPUT24), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT25), .B(G183gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G190gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n268_), .A2(new_n271_), .A3(new_n273_), .A4(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n266_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT21), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(KEYINPUT21), .ZN(new_n281_));
  XOR2_X1   g080(.A(G197gat), .B(G204gat), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n278_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n258_), .A2(new_n259_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n265_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(new_n268_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n271_), .ZN(new_n291_));
  INV_X1    g090(.A(G183gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT25), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT25), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(G183gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n295_), .A3(KEYINPUT84), .ZN(new_n296_));
  OR3_X1    g095(.A1(new_n294_), .A2(KEYINPUT84), .A3(G183gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G190gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT26), .B1(new_n299_), .B2(KEYINPUT85), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT26), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(G190gat), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n291_), .B1(new_n298_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n273_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n294_), .A2(KEYINPUT84), .A3(G183gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(new_n274_), .B2(KEYINPUT84), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n300_), .A2(new_n303_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n306_), .B(new_n271_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n264_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n290_), .B1(new_n307_), .B2(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(KEYINPUT20), .B(new_n286_), .C1(new_n314_), .C2(new_n285_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT19), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT20), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n314_), .B2(new_n285_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n278_), .A2(new_n285_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n318_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G8gat), .B(G36gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  NOR2_X1   g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n319_), .B2(new_n324_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT27), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n278_), .B(KEYINPUT101), .ZN(new_n336_));
  INV_X1    g135(.A(new_n285_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n318_), .B1(new_n338_), .B2(new_n321_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n315_), .A2(new_n317_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(new_n330_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT27), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n342_), .A2(new_n343_), .A3(new_n333_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n335_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G71gat), .B(G99gat), .ZN(new_n346_));
  INV_X1    g145(.A(G15gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G227gat), .ZN(new_n350_));
  INV_X1    g149(.A(G233gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n271_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n272_), .B1(new_n353_), .B2(KEYINPUT86), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n264_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n355_));
  AOI211_X1 g154(.A(new_n352_), .B(new_n289_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n352_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n310_), .B1(new_n297_), .B2(new_n296_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT86), .B1(new_n358_), .B2(new_n291_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n359_), .A2(new_n311_), .A3(new_n312_), .A4(new_n273_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n360_), .B2(new_n290_), .ZN(new_n361_));
  OAI21_X1  g160(.A(G43gat), .B1(new_n356_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT88), .B(KEYINPUT30), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n314_), .A2(new_n352_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n357_), .A3(new_n290_), .ZN(new_n365_));
  INV_X1    g164(.A(G43gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n362_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n363_), .B1(new_n362_), .B2(new_n367_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n349_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n363_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n356_), .A2(new_n361_), .A3(G43gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n366_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n362_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n348_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n370_), .A2(KEYINPUT90), .A3(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n238_), .B(KEYINPUT31), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n370_), .A2(new_n376_), .A3(KEYINPUT90), .A4(new_n378_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT96), .B(G22gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n337_), .B1(new_n224_), .B2(KEYINPUT29), .ZN(new_n386_));
  INV_X1    g185(.A(G50gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n224_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT28), .B1(new_n224_), .B2(KEYINPUT29), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(G228gat), .A3(G233gat), .A4(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n391_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(new_n389_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n388_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n388_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n385_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(new_n395_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n388_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n388_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(new_n384_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n398_), .A2(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n380_), .A2(new_n381_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n255_), .B(new_n345_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n380_), .A2(new_n381_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT100), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT33), .B1(new_n254_), .B2(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n241_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n240_), .A2(new_n243_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n410_), .B2(KEYINPUT33), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n251_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n410_), .A2(KEYINPUT33), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n246_), .A2(new_n252_), .A3(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n411_), .A2(new_n334_), .A3(new_n415_), .A4(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n325_), .A2(new_n419_), .ZN(new_n420_));
  OAI221_X1 g219(.A(new_n420_), .B1(new_n341_), .B2(new_n419_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n404_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n409_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n407_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT68), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT7), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G99gat), .A2(G106gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n426_), .B(new_n427_), .C1(G99gat), .C2(G106gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT69), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G99gat), .A2(G106gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n431_), .A2(KEYINPUT69), .A3(new_n432_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n435_), .A2(new_n438_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G85gat), .B(G92gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(KEYINPUT8), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT8), .ZN(new_n445_));
  INV_X1    g244(.A(new_n439_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT67), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n438_), .A2(new_n449_), .A3(new_n439_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n448_), .A2(new_n450_), .B1(new_n432_), .B2(new_n431_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n445_), .B1(new_n451_), .B2(new_n442_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n248_), .A2(KEYINPUT64), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT64), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G85gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n455_), .A3(G92gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT9), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT65), .ZN(new_n459_));
  OR2_X1    g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n456_), .A2(new_n461_), .A3(new_n457_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n463_), .B(KEYINPUT66), .Z(new_n464_));
  NAND4_X1  g263(.A1(new_n459_), .A2(new_n460_), .A3(new_n462_), .A4(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT10), .B(G99gat), .Z(new_n466_));
  INV_X1    g265(.A(G106gat), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n448_), .A2(new_n450_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n444_), .A2(new_n452_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT71), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n451_), .A2(new_n442_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n473_), .A2(new_n445_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(KEYINPUT71), .A3(new_n444_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G57gat), .B(G64gat), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n479_));
  XOR2_X1   g278(.A(G71gat), .B(G78gat), .Z(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n479_), .A2(new_n480_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT12), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n476_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n483_), .B(KEYINPUT70), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n470_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n484_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n487_), .A2(new_n470_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G230gat), .A2(G233gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n486_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT72), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n476_), .A2(new_n485_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT72), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n493_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n488_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n492_), .B1(new_n500_), .B2(new_n490_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G120gat), .B(G148gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(G204gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT5), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(new_n257_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n499_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT13), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT13), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n508_), .A2(new_n512_), .A3(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT73), .B(G43gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(G50gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(G29gat), .B(G36gat), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n516_), .B(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT15), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n516_), .B(new_n517_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT15), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT77), .B(G22gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(new_n347_), .ZN(new_n526_));
  INV_X1    g325(.A(G1gat), .ZN(new_n527_));
  INV_X1    g326(.A(G8gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G1gat), .B(G8gat), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n531_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n524_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n521_), .A3(new_n533_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n519_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n537_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(G229gat), .A3(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n269_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(G197gat), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(KEYINPUT82), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT82), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n549_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n548_), .A2(new_n550_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT83), .Z(new_n552_));
  AND3_X1   g351(.A1(new_n425_), .A2(new_n514_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n534_), .B(new_n554_), .Z(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT78), .Z(new_n556_));
  INV_X1    g355(.A(new_n483_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n555_), .B(KEYINPUT78), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n483_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G127gat), .B(G155gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n558_), .A2(new_n560_), .A3(KEYINPUT17), .A4(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n555_), .B(new_n487_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n565_), .B(KEYINPUT17), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT80), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT81), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT81), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n573_), .A3(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT74), .B(G134gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G162gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(KEYINPUT36), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n520_), .A2(new_n523_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n470_), .A2(new_n519_), .ZN(new_n587_));
  OAI211_X1 g386(.A(KEYINPUT35), .B(new_n584_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT71), .B1(new_n474_), .B2(new_n444_), .ZN(new_n589_));
  AND4_X1   g388(.A1(KEYINPUT71), .A2(new_n444_), .A3(new_n452_), .A4(new_n469_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n524_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n593_));
  INV_X1    g392(.A(new_n587_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .A4(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n582_), .B1(new_n588_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n581_), .A2(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n582_), .B(KEYINPUT75), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n598_), .A2(KEYINPUT37), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT76), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n588_), .A2(new_n595_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n582_), .ZN(new_n604_));
  AND4_X1   g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .A4(new_n597_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n602_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n600_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n601_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n576_), .A2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n553_), .A2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n255_), .B(KEYINPUT102), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n612_), .A2(new_n527_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT104), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n615_), .B1(new_n616_), .B2(KEYINPUT38), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n618_));
  INV_X1    g417(.A(new_n607_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n407_), .B2(new_n424_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n571_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n551_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n514_), .A4(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT103), .ZN(new_n624_));
  INV_X1    g423(.A(new_n255_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI221_X1 g425(.A(new_n617_), .B1(new_n618_), .B2(new_n615_), .C1(new_n527_), .C2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT105), .Z(G1324gat));
  OAI21_X1  g427(.A(G8gat), .B1(new_n623_), .B2(new_n345_), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT106), .B(KEYINPUT39), .Z(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n345_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n612_), .A2(new_n528_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n629_), .A2(new_n631_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT107), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT40), .ZN(G1325gat));
  AOI21_X1  g437(.A(new_n347_), .B1(new_n624_), .B2(new_n408_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT41), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n612_), .A2(new_n347_), .A3(new_n408_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1326gat));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n624_), .B2(new_n404_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT42), .Z(new_n645_));
  NAND3_X1  g444(.A1(new_n612_), .A2(new_n643_), .A3(new_n404_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(new_n514_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n648_), .A2(new_n575_), .A3(new_n551_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n425_), .B2(new_n610_), .ZN(new_n651_));
  AOI211_X1 g450(.A(KEYINPUT43), .B(new_n609_), .C1(new_n407_), .C2(new_n424_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n649_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n649_), .B(KEYINPUT44), .C1(new_n651_), .C2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G29gat), .B1(new_n657_), .B2(new_n613_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n553_), .A2(new_n576_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n619_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(G29gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n255_), .B2(new_n661_), .ZN(G1328gat));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n655_), .A2(new_n633_), .A3(new_n656_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT108), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n655_), .A2(new_n666_), .A3(new_n633_), .A4(new_n656_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(G36gat), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n660_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n345_), .A2(G36gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT45), .B1(new_n660_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n663_), .B1(new_n668_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n668_), .B2(new_n675_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT46), .ZN(new_n679_));
  OAI22_X1  g478(.A1(KEYINPUT110), .A2(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n668_), .A2(new_n675_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT109), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n677_), .A3(KEYINPUT46), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1329gat));
  NOR3_X1   g483(.A1(new_n657_), .A2(new_n366_), .A3(new_n409_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n669_), .A2(new_n408_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n366_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g487(.A(G50gat), .B1(new_n657_), .B2(new_n423_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n669_), .A2(new_n387_), .A3(new_n404_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1331gat));
  NAND2_X1  g490(.A1(new_n611_), .A2(new_n648_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n693_), .A2(KEYINPUT111), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n622_), .B1(new_n693_), .B2(KEYINPUT111), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(new_n425_), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G57gat), .B1(new_n696_), .B2(new_n614_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n552_), .ZN(new_n698_));
  AND4_X1   g497(.A1(new_n575_), .A2(new_n620_), .A3(new_n648_), .A4(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT112), .B(G57gat), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n255_), .A2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n699_), .B2(new_n701_), .ZN(G1332gat));
  INV_X1    g501(.A(G64gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n696_), .A2(new_n703_), .A3(new_n633_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n699_), .B2(new_n633_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT48), .Z(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1333gat));
  INV_X1    g506(.A(G71gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n696_), .A2(new_n708_), .A3(new_n408_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n699_), .B2(new_n408_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT49), .Z(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1334gat));
  INV_X1    g511(.A(G78gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n696_), .A2(new_n713_), .A3(new_n404_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n699_), .B2(new_n404_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT50), .Z(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1335gat));
  NOR3_X1   g516(.A1(new_n575_), .A2(new_n514_), .A3(new_n622_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n718_), .A2(new_n619_), .A3(new_n425_), .ZN(new_n719_));
  AOI21_X1  g518(.A(G85gat), .B1(new_n719_), .B2(new_n614_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n651_), .A2(new_n652_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(new_n718_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n625_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(G1336gat));
  AOI21_X1  g523(.A(G92gat), .B1(new_n719_), .B2(new_n633_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n633_), .A2(G92gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n722_), .B2(new_n726_), .ZN(G1337gat));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(KEYINPUT51), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n719_), .A2(new_n466_), .A3(new_n408_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT113), .Z(new_n731_));
  NAND2_X1  g530(.A1(new_n722_), .A2(new_n408_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G99gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n729_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n728_), .A2(KEYINPUT51), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(G1338gat));
  NAND3_X1  g535(.A1(new_n719_), .A2(new_n467_), .A3(new_n404_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n722_), .A2(new_n404_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G106gat), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT52), .B(new_n467_), .C1(new_n722_), .C2(new_n404_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g542(.A(G113gat), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT118), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT55), .B1(new_n495_), .B2(new_n498_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n490_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n496_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n492_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n496_), .A2(KEYINPUT55), .A3(new_n493_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT56), .B(new_n507_), .C1(new_n746_), .C2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n551_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n507_), .B1(new_n746_), .B2(new_n751_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n754_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n752_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n759_), .A3(new_n509_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n535_), .A2(new_n537_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n536_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n762_), .B2(new_n761_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n547_), .B1(new_n540_), .B2(new_n536_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n548_), .A2(new_n550_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT117), .B1(new_n764_), .B2(new_n765_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n510_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n619_), .B1(new_n760_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n745_), .B1(new_n773_), .B2(KEYINPUT57), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(KEYINPUT57), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  INV_X1    g575(.A(new_n509_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n758_), .B2(new_n752_), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n778_), .A2(new_n755_), .B1(new_n510_), .B2(new_n771_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT118), .B(new_n776_), .C1(new_n779_), .C2(new_n619_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n777_), .B1(new_n753_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n756_), .A2(new_n757_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT119), .A3(new_n752_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n784_), .A3(new_n771_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n782_), .A2(new_n784_), .A3(KEYINPUT58), .A4(new_n771_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n610_), .A3(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n774_), .A2(new_n775_), .A3(new_n780_), .A4(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n571_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n698_), .A2(new_n575_), .A3(new_n609_), .ZN(new_n792_));
  OR3_X1    g591(.A1(new_n792_), .A2(new_n648_), .A3(KEYINPUT54), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT54), .B1(new_n792_), .B2(new_n648_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n614_), .A2(new_n345_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n406_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n744_), .B1(new_n800_), .B2(new_n551_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT120), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n744_), .C1(new_n800_), .C2(new_n551_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n790_), .A2(new_n571_), .B1(new_n794_), .B2(new_n793_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n799_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT59), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n776_), .B1(new_n779_), .B2(new_n619_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n775_), .A2(new_n808_), .A3(new_n789_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n576_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n795_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n799_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n807_), .A2(G113gat), .A3(new_n552_), .A4(new_n813_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n802_), .A2(new_n804_), .A3(new_n814_), .ZN(G1340gat));
  AOI21_X1  g614(.A(new_n806_), .B1(new_n791_), .B2(new_n795_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n813_), .B(new_n648_), .C1(new_n816_), .C2(new_n812_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT122), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n807_), .A2(new_n819_), .A3(new_n648_), .A4(new_n813_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(G120gat), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(G120gat), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n822_), .A2(KEYINPUT60), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n514_), .B2(KEYINPUT60), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n816_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT121), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n821_), .A2(new_n826_), .ZN(G1341gat));
  INV_X1    g626(.A(G127gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n800_), .B2(new_n576_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT123), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n828_), .C1(new_n800_), .C2(new_n576_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n807_), .A2(G127gat), .A3(new_n621_), .A4(new_n813_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n830_), .A2(new_n832_), .A3(new_n833_), .ZN(G1342gat));
  AOI21_X1  g633(.A(G134gat), .B1(new_n816_), .B2(new_n619_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n807_), .A2(new_n610_), .A3(new_n813_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g636(.A(new_n405_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n797_), .A2(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT124), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n796_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT125), .B1(new_n805_), .B2(new_n840_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n551_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT126), .B(G141gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1344gat));
  AOI21_X1  g646(.A(new_n514_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n848_));
  INV_X1    g647(.A(G148gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1345gat));
  AOI21_X1  g649(.A(new_n576_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT61), .B(G155gat), .Z(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1346gat));
  NAND2_X1  g652(.A1(new_n843_), .A2(new_n844_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G162gat), .B1(new_n854_), .B2(new_n619_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n609_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(G162gat), .B2(new_n856_), .ZN(G1347gat));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n614_), .A2(new_n345_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n811_), .A2(new_n406_), .A3(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n551_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n858_), .B1(new_n861_), .B2(new_n269_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n256_), .ZN(new_n863_));
  OAI211_X1 g662(.A(KEYINPUT62), .B(G169gat), .C1(new_n860_), .C2(new_n551_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(G1348gat));
  INV_X1    g664(.A(new_n860_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G176gat), .B1(new_n866_), .B2(new_n648_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n805_), .A2(new_n404_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n859_), .A2(G176gat), .A3(new_n408_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n514_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n868_), .B2(new_n870_), .ZN(G1349gat));
  NOR3_X1   g670(.A1(new_n860_), .A2(new_n571_), .A3(new_n274_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n868_), .A2(new_n575_), .A3(new_n408_), .A4(new_n859_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n292_), .ZN(G1350gat));
  NAND3_X1  g673(.A1(new_n866_), .A2(new_n619_), .A3(new_n275_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G190gat), .B1(new_n860_), .B2(new_n609_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1351gat));
  NOR2_X1   g676(.A1(new_n805_), .A2(new_n625_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n838_), .A2(new_n345_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n622_), .A3(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n648_), .A3(new_n879_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT127), .B(G204gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1353gat));
  NAND3_X1  g683(.A1(new_n878_), .A2(new_n621_), .A3(new_n879_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT63), .B(G211gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n885_), .B2(new_n888_), .ZN(G1354gat));
  AND3_X1   g688(.A1(new_n878_), .A2(new_n619_), .A3(new_n879_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n878_), .A2(new_n610_), .A3(new_n879_), .ZN(new_n891_));
  MUX2_X1   g690(.A(new_n890_), .B(new_n891_), .S(G218gat), .Z(G1355gat));
endmodule


