//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT2), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n204_), .A3(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT85), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT83), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n202_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n210_), .A2(KEYINPUT1), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(KEYINPUT1), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT84), .ZN(new_n218_));
  AOI211_X1 g017(.A(new_n205_), .B(new_n214_), .C1(new_n216_), .C2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G127gat), .B(G134gat), .Z(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(G113gat), .ZN(new_n222_));
  INV_X1    g021(.A(G120gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n224_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n226_), .B1(new_n213_), .B2(new_n219_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(KEYINPUT4), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G225gat), .A2(G233gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT93), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT94), .B(KEYINPUT4), .Z(new_n231_));
  OR2_X1    g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT95), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n225_), .A2(new_n227_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n230_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n228_), .A2(new_n232_), .A3(KEYINPUT95), .A4(new_n230_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT0), .B(G57gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(G85gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(G1gat), .B(G29gat), .Z(new_n243_));
  XOR2_X1   g042(.A(new_n242_), .B(new_n243_), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n235_), .A2(new_n238_), .A3(new_n239_), .A4(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT20), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT23), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(G183gat), .B2(G190gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT90), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT22), .B(G169gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT89), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n253_), .B(new_n254_), .C1(G176gat), .C2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT25), .B(G183gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G169gat), .ZN(new_n261_));
  INV_X1    g060(.A(G176gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n263_), .A2(KEYINPUT24), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(KEYINPUT24), .A3(new_n254_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n260_), .A2(new_n251_), .A3(new_n264_), .A4(new_n265_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n257_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT21), .ZN(new_n268_));
  XOR2_X1   g067(.A(G211gat), .B(G218gat), .Z(new_n269_));
  INV_X1    g068(.A(G204gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(G197gat), .ZN(new_n271_));
  AOI211_X1 g070(.A(new_n268_), .B(new_n269_), .C1(KEYINPUT87), .C2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G197gat), .B(G204gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n268_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n249_), .B1(new_n267_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n255_), .A2(new_n262_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n252_), .A2(new_n254_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n266_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n277_), .B1(new_n276_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT19), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  OR3_X1    g085(.A1(new_n267_), .A2(KEYINPUT91), .A3(new_n276_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n249_), .B1(new_n276_), .B2(new_n281_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT91), .B1(new_n267_), .B2(new_n276_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n287_), .A2(new_n284_), .A3(new_n288_), .A4(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT32), .ZN(new_n292_));
  XOR2_X1   g091(.A(G8gat), .B(G36gat), .Z(new_n293_));
  XNOR2_X1  g092(.A(G64gat), .B(G92gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n291_), .B1(new_n292_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n282_), .A2(new_n284_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n287_), .A2(new_n285_), .A3(new_n288_), .A4(new_n289_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(KEYINPUT32), .A3(new_n297_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n248_), .A2(new_n299_), .A3(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n228_), .A2(new_n237_), .A3(new_n232_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n236_), .A2(new_n230_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n306_), .A2(KEYINPUT96), .A3(new_n244_), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT96), .B1(new_n306_), .B2(new_n244_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT97), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT33), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n247_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n291_), .B(new_n298_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n247_), .A2(new_n312_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n304_), .B1(new_n311_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT29), .B1(new_n213_), .B2(new_n219_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n276_), .ZN(new_n319_));
  INV_X1    g118(.A(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT86), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(G228gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(G228gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n320_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(new_n319_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G78gat), .B(G106gat), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OR3_X1    g130(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n331_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n213_), .A2(KEYINPUT29), .A3(new_n219_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G22gat), .B(G50gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT28), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n335_), .B(new_n337_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(KEYINPUT88), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n334_), .B(new_n340_), .Z(new_n341_));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT30), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n280_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G15gat), .B(G43gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n348_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n347_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n350_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n343_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n345_), .A2(new_n346_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n353_), .A2(new_n354_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n349_), .A2(new_n350_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(new_n342_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n357_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n224_), .B(KEYINPUT31), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n317_), .A2(new_n341_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n341_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n248_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n366_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n341_), .A3(new_n364_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n291_), .A2(new_n297_), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n375_), .B(KEYINPUT99), .Z(new_n376_));
  INV_X1    g175(.A(KEYINPUT98), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n302_), .B2(new_n298_), .ZN(new_n378_));
  AOI211_X1 g177(.A(KEYINPUT98), .B(new_n297_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(KEYINPUT27), .A3(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n381_), .B1(KEYINPUT27), .B2(new_n314_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n368_), .B1(new_n374_), .B2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(KEYINPUT77), .B(G1gat), .Z(new_n384_));
  INV_X1    g183(.A(G8gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT14), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G15gat), .B(G22gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G1gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G8gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n388_), .B(G1gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n385_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G50gat), .ZN(new_n395_));
  INV_X1    g194(.A(G29gat), .ZN(new_n396_));
  INV_X1    g195(.A(G36gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G43gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G29gat), .A2(G36gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n399_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n395_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(G50gat), .A3(new_n401_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n394_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n391_), .A2(new_n393_), .A3(new_n407_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G229gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT15), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n407_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n404_), .A2(new_n406_), .A3(KEYINPUT15), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n409_), .B(new_n412_), .C1(new_n394_), .C2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G113gat), .B(G141gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(new_n261_), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n423_), .B(G197gat), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(KEYINPUT80), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n414_), .B(new_n420_), .C1(KEYINPUT80), .C2(new_n425_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n430_));
  NOR2_X1   g229(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n431_));
  OAI22_X1  g230(.A1(new_n430_), .A2(new_n431_), .B1(G99gat), .B2(G106gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G99gat), .A2(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT6), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(G99gat), .A3(G106gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G99gat), .A2(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n432_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(G85gat), .A2(G92gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT8), .B1(new_n441_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT68), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n435_), .B1(G99gat), .B2(G106gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n433_), .A2(KEYINPUT6), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n434_), .A2(new_n436_), .A3(KEYINPUT68), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n438_), .B1(new_n453_), .B2(new_n439_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n440_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT69), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT69), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n432_), .A2(new_n457_), .A3(new_n440_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n452_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n445_), .A2(KEYINPUT8), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n446_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n462_));
  NOR2_X1   g261(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n442_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT65), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n444_), .B1(new_n443_), .B2(KEYINPUT9), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT65), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n467_), .B(new_n442_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT66), .ZN(new_n470_));
  XOR2_X1   g269(.A(KEYINPUT10), .B(G99gat), .Z(new_n471_));
  INV_X1    g270(.A(G106gat), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n471_), .A2(new_n472_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT66), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n465_), .A2(new_n474_), .A3(new_n466_), .A4(new_n468_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n461_), .A2(new_n476_), .A3(new_n408_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n461_), .A2(new_n476_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n478_), .A2(KEYINPUT72), .A3(new_n418_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT72), .B1(new_n478_), .B2(new_n418_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n477_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G232gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT34), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(KEYINPUT35), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n478_), .A2(new_n418_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT72), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n478_), .A2(KEYINPUT72), .A3(new_n418_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n483_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n491_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n489_), .A2(new_n493_), .A3(new_n494_), .A4(new_n477_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G190gat), .B(G218gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G134gat), .ZN(new_n497_));
  INV_X1    g296(.A(G162gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n501_), .B(KEYINPUT74), .Z(new_n502_));
  NAND3_X1  g301(.A1(new_n484_), .A2(new_n495_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT75), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n484_), .A2(new_n495_), .A3(KEYINPUT75), .A4(new_n502_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n484_), .A2(new_n495_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n499_), .B(KEYINPUT36), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(KEYINPUT76), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n505_), .A2(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT76), .A3(KEYINPUT37), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT13), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT71), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n517_), .A2(KEYINPUT71), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G230gat), .A2(G233gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n524_));
  XOR2_X1   g323(.A(G71gat), .B(G78gat), .Z(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n461_), .A2(new_n476_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n461_), .B2(new_n476_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n521_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G120gat), .B(G148gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n270_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT5), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(new_n262_), .ZN(new_n535_));
  AOI211_X1 g334(.A(KEYINPUT12), .B(new_n528_), .C1(new_n461_), .C2(new_n476_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n529_), .A2(new_n530_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(KEYINPUT12), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n531_), .B(new_n535_), .C1(new_n538_), .C2(new_n521_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n535_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n528_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n478_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n461_), .A2(new_n476_), .A3(new_n528_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(KEYINPUT12), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT12), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n530_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n521_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n531_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n540_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n539_), .A2(new_n549_), .A3(KEYINPUT70), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT70), .B1(new_n539_), .B2(new_n549_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n518_), .B(new_n519_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n544_), .A2(new_n546_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n520_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n535_), .B1(new_n555_), .B2(new_n531_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n547_), .A2(new_n548_), .A3(new_n540_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n553_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n539_), .A2(new_n549_), .A3(KEYINPUT70), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n558_), .A2(KEYINPUT71), .A3(new_n517_), .A4(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n394_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n528_), .B(KEYINPUT78), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT16), .B(G183gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G211gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(G127gat), .B(G155gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n562_), .A2(new_n564_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n562_), .B(new_n563_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n569_), .A2(new_n570_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n552_), .A2(new_n560_), .A3(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n516_), .A2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n429_), .B1(new_n578_), .B2(KEYINPUT79), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n383_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n578_), .A2(KEYINPUT79), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(new_n371_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n384_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n584_), .B2(new_n384_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT38), .ZN(new_n588_));
  OR3_X1    g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n552_), .A2(new_n560_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n427_), .A2(new_n428_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT101), .Z(new_n594_));
  INV_X1    g393(.A(new_n576_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n595_), .A2(new_n514_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n383_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G1gat), .B1(new_n598_), .B2(new_n371_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n588_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n589_), .A2(new_n599_), .A3(new_n600_), .ZN(G1324gat));
  NAND3_X1  g400(.A1(new_n582_), .A2(new_n385_), .A3(new_n382_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n383_), .A2(new_n594_), .A3(new_n382_), .A4(new_n596_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n603_), .A2(new_n604_), .A3(G8gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n603_), .B2(G8gat), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT102), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(KEYINPUT102), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n608_), .A2(KEYINPUT40), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT40), .B1(new_n608_), .B2(new_n609_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(G1325gat));
  INV_X1    g411(.A(G15gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n367_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n597_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n582_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n597_), .B2(new_n369_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT42), .Z(new_n621_));
  NAND2_X1  g420(.A1(new_n369_), .A2(new_n619_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT103), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n621_), .B1(new_n583_), .B2(new_n623_), .ZN(G1327gat));
  AND2_X1   g423(.A1(new_n383_), .A2(new_n514_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n593_), .A2(new_n576_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n396_), .A3(new_n248_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT43), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n383_), .A2(new_n630_), .A3(new_n516_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n383_), .B2(new_n516_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n594_), .B(new_n595_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT44), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n383_), .A2(new_n516_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT43), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n383_), .A2(new_n630_), .A3(new_n516_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n639_), .A2(KEYINPUT44), .A3(new_n594_), .A4(new_n595_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n635_), .A2(new_n640_), .A3(new_n248_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n641_), .A2(KEYINPUT104), .A3(G29gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT104), .B1(new_n641_), .B2(G29gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n629_), .B1(new_n642_), .B2(new_n643_), .ZN(G1328gat));
  NAND3_X1  g443(.A1(new_n635_), .A2(new_n640_), .A3(new_n382_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G36gat), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n625_), .A2(new_n397_), .A3(new_n382_), .A4(new_n626_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT45), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n646_), .A2(KEYINPUT46), .A3(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1329gat));
  NOR3_X1   g452(.A1(new_n627_), .A2(G43gat), .A3(new_n367_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n635_), .A2(new_n640_), .A3(new_n614_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(G43gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g456(.A(G50gat), .B1(new_n628_), .B2(new_n369_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n635_), .A2(new_n640_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n341_), .A2(new_n395_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n658_), .B1(new_n659_), .B2(new_n660_), .ZN(G1331gat));
  NOR2_X1   g460(.A1(new_n591_), .A2(new_n592_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n383_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n516_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n663_), .A2(new_n576_), .A3(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G57gat), .B1(new_n665_), .B2(new_n248_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n663_), .A2(new_n596_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(new_n248_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(G57gat), .B2(new_n668_), .ZN(G1332gat));
  INV_X1    g468(.A(G64gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n667_), .B2(new_n382_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT48), .Z(new_n672_));
  NAND3_X1  g471(.A1(new_n665_), .A2(new_n670_), .A3(new_n382_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1333gat));
  INV_X1    g473(.A(G71gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n667_), .B2(new_n614_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT49), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n665_), .A2(new_n675_), .A3(new_n614_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1334gat));
  INV_X1    g478(.A(G78gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n667_), .B2(new_n369_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT50), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n665_), .A2(new_n680_), .A3(new_n369_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1335gat));
  INV_X1    g483(.A(G85gat), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n662_), .A2(new_n595_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n625_), .A2(new_n686_), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n686_), .B1(new_n625_), .B2(new_n688_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n685_), .B1(new_n691_), .B2(new_n371_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n692_), .A2(KEYINPUT106), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(KEYINPUT106), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n687_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n371_), .A2(new_n685_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n693_), .A2(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(G1336gat));
  INV_X1    g496(.A(new_n691_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G92gat), .B1(new_n698_), .B2(new_n382_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n382_), .A2(G92gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n695_), .B2(new_n700_), .ZN(G1337gat));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n614_), .A2(new_n471_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n691_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(G99gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n695_), .B2(new_n614_), .ZN(new_n706_));
  OR3_X1    g505(.A1(new_n704_), .A2(KEYINPUT51), .A3(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT51), .B1(new_n704_), .B2(new_n706_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1338gat));
  NAND3_X1  g508(.A1(new_n698_), .A2(new_n472_), .A3(new_n369_), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT52), .B(new_n472_), .C1(new_n695_), .C2(new_n369_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT52), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n695_), .A2(new_n369_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(G106gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT53), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT53), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n710_), .B(new_n717_), .C1(new_n714_), .C2(new_n711_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1339gat));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n555_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT112), .B1(new_n547_), .B2(new_n721_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n547_), .A2(KEYINPUT55), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n538_), .A2(new_n521_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n723_), .A2(new_n724_), .A3(new_n725_), .A4(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(KEYINPUT56), .A3(new_n540_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT56), .B1(new_n727_), .B2(new_n540_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n592_), .B(new_n539_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n411_), .A2(new_n412_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n409_), .B(new_n413_), .C1(new_n394_), .C2(new_n419_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n424_), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n414_), .A2(new_n425_), .A3(new_n420_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n732_), .A2(KEYINPUT113), .A3(new_n733_), .A4(new_n424_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n739_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n514_), .B1(new_n731_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(KEYINPUT57), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT57), .ZN(new_n745_));
  INV_X1    g544(.A(new_n514_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n592_), .A2(new_n539_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n730_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n728_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n749_), .B2(new_n740_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n745_), .B1(new_n750_), .B2(KEYINPUT114), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n744_), .A2(new_n751_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n730_), .A2(KEYINPUT115), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n730_), .A2(KEYINPUT115), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n728_), .A3(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n739_), .A2(new_n557_), .ZN(new_n756_));
  OR2_X1    g555(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT117), .B1(KEYINPUT116), .B2(KEYINPUT58), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n759_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .A4(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n516_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n752_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n595_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n552_), .A2(new_n560_), .A3(new_n576_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n766_), .A2(new_n429_), .A3(new_n515_), .A4(new_n513_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT54), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT109), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n770_), .A3(KEYINPUT54), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n516_), .A2(new_n592_), .A3(new_n577_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(KEYINPUT108), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n767_), .B2(KEYINPUT54), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n772_), .A2(new_n778_), .A3(KEYINPUT110), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT110), .B1(new_n772_), .B2(new_n778_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n765_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n382_), .A2(new_n371_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n781_), .A2(new_n341_), .A3(new_n614_), .A4(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G113gat), .B1(new_n785_), .B2(new_n592_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(KEYINPUT59), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n784_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n429_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n790_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g590(.A(KEYINPUT60), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n784_), .B1(new_n792_), .B2(G120gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n223_), .B1(new_n591_), .B2(KEYINPUT60), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n793_), .A2(KEYINPUT118), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT118), .B1(new_n793_), .B2(new_n794_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n591_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n797_));
  OAI22_X1  g596(.A1(new_n795_), .A2(new_n796_), .B1(new_n797_), .B2(new_n223_), .ZN(G1341gat));
  AOI21_X1  g597(.A(G127gat), .B1(new_n785_), .B2(new_n576_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n787_), .A2(new_n789_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n576_), .A2(G127gat), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT119), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n799_), .B1(new_n800_), .B2(new_n802_), .ZN(G1342gat));
  AOI21_X1  g602(.A(G134gat), .B1(new_n785_), .B2(new_n514_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n664_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(G134gat), .ZN(G1343gat));
  NAND3_X1  g605(.A1(new_n781_), .A2(new_n369_), .A3(new_n367_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n807_), .A2(new_n782_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(new_n429_), .ZN(new_n809_));
  INV_X1    g608(.A(G141gat), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(G1344gat));
  NOR2_X1   g610(.A1(new_n808_), .A2(new_n591_), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT120), .B(G148gat), .Z(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(G1345gat));
  NOR2_X1   g613(.A1(new_n808_), .A2(new_n595_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(G155gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n815_), .B(new_n817_), .ZN(G1346gat));
  NOR3_X1   g617(.A1(new_n808_), .A2(new_n498_), .A3(new_n664_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n808_), .A2(new_n746_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n498_), .B2(new_n820_), .ZN(G1347gat));
  AOI21_X1  g620(.A(KEYINPUT108), .B1(new_n773_), .B2(new_n774_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n767_), .A2(new_n776_), .A3(KEYINPUT54), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n767_), .A2(new_n770_), .A3(KEYINPUT54), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n770_), .B1(new_n767_), .B2(KEYINPUT54), .ZN(new_n825_));
  OAI22_X1  g624(.A1(new_n822_), .A2(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n772_), .A2(new_n778_), .A3(KEYINPUT110), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n369_), .B1(new_n830_), .B2(new_n765_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n382_), .A2(new_n371_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n367_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n592_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n834_), .A2(new_n835_), .A3(G169gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n834_), .B2(G169gat), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n576_), .B1(new_n752_), .B2(new_n763_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n833_), .ZN(new_n842_));
  NOR4_X1   g641(.A1(new_n841_), .A2(KEYINPUT122), .A3(new_n369_), .A4(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n839_), .A2(new_n843_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n429_), .A2(new_n256_), .ZN(new_n845_));
  OAI22_X1  g644(.A1(new_n836_), .A2(new_n837_), .B1(new_n844_), .B2(new_n845_), .ZN(G1348gat));
  NAND3_X1  g645(.A1(new_n781_), .A2(new_n341_), .A3(new_n833_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n847_), .A2(new_n262_), .A3(new_n591_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(KEYINPUT122), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n831_), .A2(new_n838_), .A3(new_n833_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n591_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT123), .B1(new_n851_), .B2(G176gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n590_), .B1(new_n839_), .B2(new_n843_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n262_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n848_), .B1(new_n852_), .B2(new_n855_), .ZN(G1349gat));
  NOR3_X1   g655(.A1(new_n844_), .A2(new_n258_), .A3(new_n595_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n847_), .A2(new_n595_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(G183gat), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1350gat));
  OAI21_X1  g659(.A(G190gat), .B1(new_n844_), .B2(new_n664_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n514_), .A2(new_n259_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n844_), .B2(new_n862_), .ZN(G1351gat));
  INV_X1    g662(.A(new_n832_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n781_), .A2(new_n369_), .A3(new_n367_), .A4(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n592_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g667(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n865_), .A2(new_n591_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n870_), .B2(new_n869_), .ZN(G1353gat));
  AOI21_X1  g672(.A(new_n595_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT125), .B1(new_n865_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n865_), .A2(KEYINPUT125), .A3(new_n875_), .ZN(new_n878_));
  OAI22_X1  g677(.A1(new_n877_), .A2(new_n878_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n878_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n881_), .A3(new_n876_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1354gat));
  NAND2_X1  g682(.A1(new_n516_), .A2(G218gat), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(KEYINPUT126), .Z(new_n885_));
  NAND2_X1  g684(.A1(new_n866_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(G218gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n865_), .B2(new_n746_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT127), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n886_), .A2(new_n891_), .A3(new_n888_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1355gat));
endmodule


