//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n597_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT8), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT64), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  AND2_X1   g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n206_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G85gat), .B(G92gat), .Z(new_n215_));
  AOI21_X1  g014(.A(new_n204_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n204_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n212_), .A2(new_n213_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n207_), .A2(KEYINPUT64), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT65), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n206_), .B1(new_n219_), .B2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n217_), .B1(new_n226_), .B2(KEYINPUT66), .ZN(new_n227_));
  INV_X1    g026(.A(new_n206_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n218_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n223_), .A2(KEYINPUT65), .A3(new_n224_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n216_), .B1(new_n227_), .B2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n219_), .A2(new_n225_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT10), .B(G99gat), .ZN(new_n238_));
  OAI221_X1 g037(.A(new_n236_), .B1(KEYINPUT9), .B2(new_n237_), .C1(G106gat), .C2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n235_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n203_), .B1(new_n234_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n216_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n204_), .B(new_n215_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n226_), .A2(KEYINPUT66), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n240_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(KEYINPUT67), .A3(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G57gat), .B(G64gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G71gat), .B(G78gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(KEYINPUT11), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n248_), .A2(KEYINPUT11), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(new_n249_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n248_), .A2(KEYINPUT11), .ZN(new_n253_));
  OAI211_X1 g052(.A(KEYINPUT12), .B(new_n250_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n241_), .A2(new_n247_), .A3(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n227_), .A2(new_n233_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n240_), .B1(new_n258_), .B2(new_n242_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n250_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n257_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n256_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n259_), .A2(new_n260_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n245_), .A2(new_n260_), .A3(new_n246_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n262_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT5), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G176gat), .B(G204gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n264_), .A2(new_n267_), .A3(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT69), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n264_), .A2(new_n267_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n271_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(KEYINPUT70), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT70), .B1(new_n274_), .B2(new_n276_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n202_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n276_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n277_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n280_), .A2(new_n284_), .A3(KEYINPUT71), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n290_), .A2(KEYINPUT72), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(KEYINPUT72), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT85), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT25), .B(G183gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT26), .B(G190gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT23), .ZN(new_n299_));
  OR2_X1    g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n300_), .A2(KEYINPUT24), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(KEYINPUT24), .A3(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n297_), .A2(new_n299_), .A3(new_n301_), .A4(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n299_), .B1(G183gat), .B2(G190gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT84), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT22), .B(G169gat), .ZN(new_n307_));
  INV_X1    g106(.A(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n302_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT83), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n304_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G71gat), .B(G99gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(G43gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n312_), .B(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G227gat), .A2(G233gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(G15gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT30), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n318_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n294_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n294_), .A3(new_n320_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G127gat), .B(G134gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G113gat), .B(G120gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT31), .Z(new_n327_));
  NAND3_X1  g126(.A1(new_n322_), .A2(new_n323_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n327_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n321_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G197gat), .B(G204gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT21), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT92), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G211gat), .B(G218gat), .Z(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n334_), .B2(new_n333_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n333_), .B(KEYINPUT93), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n338_), .A2(KEYINPUT21), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n310_), .A2(KEYINPUT96), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n305_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n310_), .A2(KEYINPUT96), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n304_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n349_), .B(KEYINPUT20), .C1(new_n344_), .C2(new_n312_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT19), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n340_), .A2(new_n343_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n348_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n352_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n312_), .A2(new_n344_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n353_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT18), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G64gat), .B(G92gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n353_), .A2(new_n365_), .A3(new_n360_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G85gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT0), .B(G57gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT3), .ZN(new_n379_));
  INV_X1    g178(.A(G141gat), .ZN(new_n380_));
  INV_X1    g179(.A(G148gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n377_), .B(new_n379_), .C1(KEYINPUT2), .C2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G155gat), .B(G162gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT88), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G155gat), .ZN(new_n390_));
  INV_X1    g189(.A(G162gat), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n390_), .A2(new_n391_), .A3(KEYINPUT1), .ZN(new_n392_));
  NOR2_X1   g191(.A1(G155gat), .A2(G162gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT1), .B1(new_n390_), .B2(new_n391_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n396_), .A2(new_n382_), .A3(new_n378_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n389_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n326_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n397_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n326_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n374_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT98), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(KEYINPUT98), .B(new_n374_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n405_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT97), .B1(new_n400_), .B2(KEYINPUT4), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT97), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n399_), .A2(new_n412_), .A3(new_n413_), .A4(new_n326_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n400_), .A2(KEYINPUT4), .A3(new_n403_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n408_), .B(new_n409_), .C1(new_n410_), .C2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n410_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n404_), .A2(new_n405_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n374_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n369_), .B(new_n417_), .C1(new_n420_), .C2(KEYINPUT33), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n420_), .A2(KEYINPUT33), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n418_), .A2(new_n374_), .A3(new_n419_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(new_n420_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n365_), .A2(KEYINPUT32), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n353_), .A2(new_n360_), .A3(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n350_), .A2(new_n352_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n358_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n429_), .B2(new_n425_), .ZN(new_n430_));
  OAI22_X1  g229(.A1(new_n421_), .A2(new_n422_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G22gat), .B(G50gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT91), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT89), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n401_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n401_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n436_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n443_), .A2(new_n439_), .A3(new_n435_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n433_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n435_), .B1(new_n443_), .B2(new_n439_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n440_), .A2(new_n441_), .A3(new_n436_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(new_n432_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n355_), .B1(new_n399_), .B2(KEYINPUT29), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G228gat), .A2(G233gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n450_), .A2(new_n451_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G78gat), .B(G106gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OAI22_X1  g255(.A1(new_n453_), .A2(new_n454_), .B1(KEYINPUT94), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n454_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n456_), .A2(KEYINPUT94), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n452_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n449_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT95), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT95), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n449_), .A2(new_n461_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n449_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n450_), .B(new_n451_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(new_n455_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n463_), .A2(new_n465_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n431_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n468_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n449_), .A2(new_n461_), .A3(new_n464_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n464_), .B1(new_n449_), .B2(new_n461_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n366_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n475_), .A2(KEYINPUT27), .A3(new_n368_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT27), .B1(new_n367_), .B2(new_n368_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n478_), .A3(new_n424_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n332_), .B1(new_n470_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n332_), .A2(new_n424_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n471_), .B(new_n478_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT99), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n463_), .A2(new_n465_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n485_), .A2(KEYINPUT99), .A3(new_n471_), .A4(new_n478_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n481_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n480_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  INV_X1    g288(.A(G1gat), .ZN(new_n490_));
  INV_X1    g289(.A(G8gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT14), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G1gat), .B(G8gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  NAND2_X1  g294(.A1(G231gat), .A2(G233gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(new_n260_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G127gat), .B(G155gat), .Z(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G183gat), .B(G211gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n503_), .A2(KEYINPUT17), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(KEYINPUT17), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n498_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n506_), .B1(new_n504_), .B2(new_n498_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(KEYINPUT80), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(KEYINPUT80), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G29gat), .B(G36gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT15), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n241_), .A2(new_n247_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n259_), .A2(new_n514_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n520_), .A2(new_n517_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n523_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n516_), .A2(new_n521_), .A3(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G190gat), .B(G218gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT74), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G134gat), .B(G162gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n532_), .B(KEYINPUT75), .Z(new_n533_));
  NAND3_X1  g332(.A1(new_n524_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n534_), .A2(KEYINPUT76), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n530_), .B(new_n531_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT77), .ZN(new_n537_));
  INV_X1    g336(.A(new_n526_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n525_), .B1(new_n516_), .B2(new_n521_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT78), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT78), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n542_), .B(new_n537_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n534_), .A2(KEYINPUT76), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n535_), .A2(new_n541_), .A3(new_n543_), .A4(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT37), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n540_), .A2(new_n534_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT37), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n495_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n515_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT82), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n495_), .A2(new_n514_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT81), .B1(new_n495_), .B2(new_n514_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n495_), .A2(new_n514_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n554_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G169gat), .B(G197gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n556_), .A2(new_n561_), .A3(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n565_), .B1(new_n556_), .B2(new_n561_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR4_X1   g368(.A1(new_n488_), .A2(new_n511_), .A3(new_n550_), .A4(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n293_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n424_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n490_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT38), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n289_), .A2(new_n569_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n547_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n488_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n510_), .A3(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(G1gat), .B1(new_n580_), .B2(new_n424_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n575_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n576_), .A2(new_n581_), .A3(new_n582_), .ZN(G1324gat));
  OAI21_X1  g382(.A(G8gat), .B1(new_n580_), .B2(new_n478_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT39), .ZN(new_n585_));
  INV_X1    g384(.A(new_n478_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n572_), .A2(new_n491_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(G1325gat));
  OAI21_X1  g389(.A(G15gat), .B1(new_n580_), .B2(new_n331_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT41), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n571_), .A2(G15gat), .A3(new_n331_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(G1326gat));
  OAI21_X1  g393(.A(G22gat), .B1(new_n580_), .B2(new_n469_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT42), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n469_), .A2(G22gat), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n596_), .B1(new_n571_), .B2(new_n597_), .ZN(G1327gat));
  NOR2_X1   g397(.A1(new_n488_), .A2(new_n547_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n577_), .A2(new_n511_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(G29gat), .B1(new_n601_), .B2(new_n573_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n550_), .B1(new_n480_), .B2(new_n487_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT43), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT43), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n550_), .B(new_n605_), .C1(new_n480_), .C2(new_n487_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n510_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(new_n577_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT44), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n609_), .A2(G29gat), .A3(new_n573_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n608_), .A2(KEYINPUT44), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n602_), .B1(new_n610_), .B2(new_n612_), .ZN(G1328gat));
  NOR3_X1   g412(.A1(new_n600_), .A2(G36gat), .A3(new_n478_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT45), .Z(new_n615_));
  NAND2_X1  g414(.A1(new_n609_), .A2(new_n586_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G36gat), .B1(new_n616_), .B2(new_n611_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT101), .B(KEYINPUT46), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n618_), .B(new_n620_), .ZN(G1329gat));
  AOI21_X1  g420(.A(G43gat), .B1(new_n601_), .B2(new_n332_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT102), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n612_), .A2(G43gat), .A3(new_n332_), .A4(new_n609_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(G1330gat));
  NAND2_X1  g426(.A1(new_n609_), .A2(new_n474_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G50gat), .B1(new_n628_), .B2(new_n611_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n469_), .A2(G50gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT104), .Z(new_n631_));
  OAI21_X1  g430(.A(new_n629_), .B1(new_n600_), .B2(new_n631_), .ZN(G1331gat));
  INV_X1    g431(.A(G57gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n579_), .A2(new_n510_), .A3(new_n569_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n293_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n633_), .B1(new_n635_), .B2(new_n573_), .ZN(new_n636_));
  NOR4_X1   g435(.A1(new_n488_), .A2(new_n511_), .A3(new_n550_), .A4(new_n568_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n289_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(G57gat), .A3(new_n424_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n636_), .A2(new_n639_), .ZN(G1332gat));
  OR3_X1    g439(.A1(new_n638_), .A2(G64gat), .A3(new_n478_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n635_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G64gat), .B1(new_n642_), .B2(new_n478_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(KEYINPUT48), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(KEYINPUT48), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n644_), .B2(new_n645_), .ZN(G1333gat));
  OR3_X1    g445(.A1(new_n638_), .A2(G71gat), .A3(new_n331_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n634_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n291_), .A2(new_n292_), .A3(new_n332_), .A4(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT49), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(G71gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n649_), .B2(G71gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n647_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT105), .Z(G1334gat));
  OR3_X1    g453(.A1(new_n638_), .A2(G78gat), .A3(new_n469_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G78gat), .B1(new_n642_), .B2(new_n469_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n656_), .A2(KEYINPUT50), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(KEYINPUT50), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(G1335gat));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n510_), .A2(new_n568_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n599_), .A2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n660_), .B1(new_n293_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n662_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n291_), .A2(KEYINPUT106), .A3(new_n292_), .A4(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G85gat), .B1(new_n666_), .B2(new_n573_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n604_), .A2(KEYINPUT107), .A3(new_n606_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n661_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT107), .B1(new_n604_), .B2(new_n606_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT108), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n604_), .A2(new_n606_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n670_), .A4(new_n668_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n673_), .A2(new_n678_), .A3(KEYINPUT109), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT109), .B1(new_n673_), .B2(new_n678_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n573_), .A2(G85gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n667_), .B1(new_n681_), .B2(new_n682_), .ZN(G1336gat));
  INV_X1    g482(.A(KEYINPUT110), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n586_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G92gat), .ZN(new_n686_));
  INV_X1    g485(.A(G92gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n586_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n684_), .B1(new_n686_), .B2(new_n690_), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT110), .B(new_n689_), .C1(new_n685_), .C2(G92gat), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1337gat));
  INV_X1    g492(.A(new_n238_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n666_), .A2(new_n694_), .A3(new_n332_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n673_), .A2(new_n678_), .A3(new_n332_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G99gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g498(.A(G106gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n666_), .A2(new_n700_), .A3(new_n474_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n674_), .A2(new_n474_), .A3(new_n670_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT52), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n702_), .B(G106gat), .C1(KEYINPUT111), .C2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(KEYINPUT111), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n701_), .A2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g507(.A(KEYINPUT117), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n511_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n710_), .A2(new_n280_), .A3(new_n284_), .A4(new_n569_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(KEYINPUT113), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n711_), .A2(new_n713_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT113), .B1(new_n711_), .B2(new_n713_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n274_), .A2(new_n568_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT114), .ZN(new_n720_));
  INV_X1    g519(.A(new_n266_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n256_), .A2(new_n721_), .A3(new_n261_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n264_), .A2(KEYINPUT55), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT55), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n256_), .A2(new_n261_), .A3(new_n263_), .A4(new_n724_), .ZN(new_n725_));
  AOI221_X4 g524(.A(new_n720_), .B1(new_n722_), .B2(new_n262_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n725_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n722_), .A2(new_n262_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT114), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n271_), .B1(new_n726_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT56), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(KEYINPUT56), .B(new_n271_), .C1(new_n726_), .C2(new_n729_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n719_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n553_), .A2(new_n560_), .A3(new_n555_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n564_), .B1(new_n559_), .B2(new_n554_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n566_), .A2(KEYINPUT115), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT115), .B1(new_n566_), .B2(new_n737_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n283_), .B2(new_n277_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n547_), .B1(new_n734_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT57), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT57), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(new_n547_), .C1(new_n734_), .C2(new_n741_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n274_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n740_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n727_), .A2(new_n728_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n720_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n727_), .A2(KEYINPUT114), .A3(new_n728_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT56), .B1(new_n751_), .B2(new_n271_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n733_), .ZN(new_n753_));
  OAI211_X1 g552(.A(KEYINPUT58), .B(new_n747_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n747_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT58), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n549_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n743_), .A2(new_n745_), .B1(new_n754_), .B2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n510_), .B1(new_n758_), .B2(KEYINPUT116), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n754_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n719_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n762_));
  OAI22_X1  g561(.A1(new_n278_), .A2(new_n279_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n744_), .B1(new_n764_), .B2(new_n547_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n745_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n760_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n718_), .B1(new_n759_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n484_), .A2(new_n486_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n573_), .A3(new_n332_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n709_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  OR3_X1    g572(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n774_));
  OAI211_X1 g573(.A(KEYINPUT116), .B(new_n760_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n511_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n758_), .A2(KEYINPUT116), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n774_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n772_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(KEYINPUT117), .A3(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n773_), .A2(new_n568_), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(G113gat), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT118), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n785_), .A3(new_n782_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n772_), .A2(KEYINPUT59), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n767_), .A2(new_n511_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n774_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n778_), .A2(new_n779_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(KEYINPUT59), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n569_), .A2(new_n782_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n784_), .A2(new_n786_), .B1(new_n791_), .B2(new_n792_), .ZN(G1340gat));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794_));
  INV_X1    g593(.A(G120gat), .ZN(new_n795_));
  INV_X1    g594(.A(new_n293_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n791_), .B2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n290_), .A2(KEYINPUT60), .ZN(new_n798_));
  MUX2_X1   g597(.A(KEYINPUT60), .B(new_n798_), .S(new_n795_), .Z(new_n799_));
  NAND3_X1  g598(.A1(new_n773_), .A2(new_n780_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n794_), .B1(new_n797_), .B2(new_n801_), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n789_), .B(new_n293_), .C1(new_n790_), .C2(KEYINPUT59), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT119), .B(new_n800_), .C1(new_n803_), .C2(new_n795_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1341gat));
  AND2_X1   g604(.A1(new_n773_), .A2(new_n780_), .ZN(new_n806_));
  AOI21_X1  g605(.A(G127gat), .B1(new_n806_), .B2(new_n510_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n510_), .A2(G127gat), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT120), .Z(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n791_), .B2(new_n809_), .ZN(G1342gat));
  INV_X1    g609(.A(G134gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n806_), .A2(new_n811_), .A3(new_n578_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n791_), .A2(new_n550_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n811_), .ZN(G1343gat));
  NOR4_X1   g613(.A1(new_n469_), .A2(new_n332_), .A3(new_n586_), .A4(new_n424_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n778_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(new_n569_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(new_n380_), .ZN(G1344gat));
  NOR2_X1   g617(.A1(new_n816_), .A2(new_n293_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(new_n381_), .ZN(G1345gat));
  NOR2_X1   g619(.A1(new_n816_), .A2(new_n511_), .ZN(new_n821_));
  XOR2_X1   g620(.A(KEYINPUT61), .B(G155gat), .Z(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1346gat));
  OAI21_X1  g622(.A(G162gat), .B1(new_n816_), .B2(new_n549_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n578_), .A2(new_n391_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n816_), .B2(new_n825_), .ZN(G1347gat));
  NAND2_X1  g625(.A1(new_n586_), .A2(new_n424_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(new_n331_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT121), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n469_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n758_), .A2(new_n510_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n568_), .B(new_n831_), .C1(new_n832_), .C2(new_n718_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G169gat), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n837_));
  INV_X1    g636(.A(new_n307_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n836_), .B(new_n837_), .C1(new_n838_), .C2(new_n833_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1348gat));
  AOI21_X1  g640(.A(new_n830_), .B1(new_n774_), .B2(new_n788_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G176gat), .B1(new_n842_), .B2(new_n289_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT123), .B1(new_n770_), .B2(new_n474_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n778_), .A2(new_n845_), .A3(new_n469_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n796_), .A2(G176gat), .A3(new_n829_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT124), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n851_), .A3(new_n848_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n843_), .B1(new_n850_), .B2(new_n852_), .ZN(G1349gat));
  NOR2_X1   g652(.A1(new_n511_), .A2(new_n295_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n842_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n829_), .A2(new_n510_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n857_), .B2(G183gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT125), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n860_), .B(new_n855_), .C1(new_n857_), .C2(G183gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1350gat));
  NAND2_X1  g661(.A1(new_n842_), .A2(new_n550_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G190gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n578_), .A2(new_n296_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT126), .Z(new_n866_));
  NAND2_X1  g665(.A1(new_n842_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(G1351gat));
  NOR4_X1   g667(.A1(new_n770_), .A2(new_n469_), .A3(new_n332_), .A4(new_n827_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n568_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n796_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g672(.A(new_n511_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n869_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n875_), .B(new_n876_), .Z(G1354gat));
  INV_X1    g676(.A(G218gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n869_), .A2(new_n878_), .A3(new_n578_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n869_), .A2(new_n550_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n878_), .ZN(G1355gat));
endmodule


