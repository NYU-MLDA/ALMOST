//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n583_, new_n584_, new_n585_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G85gat), .B(G92gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR3_X1   g010(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n209_), .B1(new_n213_), .B2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT8), .B1(new_n219_), .B2(KEYINPUT68), .ZN(new_n220_));
  INV_X1    g019(.A(new_n209_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n215_), .A2(new_n217_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n210_), .ZN(new_n227_));
  OAI211_X1 g026(.A(KEYINPUT68), .B(new_n221_), .C1(new_n222_), .C2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT69), .B1(new_n220_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n219_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n232_), .B(new_n221_), .C1(new_n222_), .C2(new_n227_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT67), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n221_), .B1(new_n222_), .B2(new_n227_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(KEYINPUT8), .A4(new_n228_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n230_), .A2(new_n236_), .A3(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G29gat), .B(G36gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G43gat), .B(G50gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT10), .B(G99gat), .Z(new_n246_));
  AOI21_X1  g045(.A(new_n222_), .B1(new_n225_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT9), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT65), .B(G85gat), .Z(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT66), .B(G92gat), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(KEYINPUT64), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n248_), .B1(G85gat), .B2(G92gat), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n248_), .A2(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G85gat), .A2(G92gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n247_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n242_), .A2(new_n245_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT74), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n203_), .A2(new_n205_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT75), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n207_), .B2(new_n206_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n242_), .A2(new_n258_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n245_), .B(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n263_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n208_), .B1(new_n260_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n260_), .A2(new_n208_), .A3(new_n267_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G190gat), .B(G218gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G134gat), .B(G162gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT36), .Z(new_n274_));
  NAND3_X1  g073(.A1(new_n269_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT37), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n273_), .A2(KEYINPUT36), .ZN(new_n279_));
  INV_X1    g078(.A(new_n270_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(new_n268_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n275_), .A3(KEYINPUT37), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G64gat), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n288_));
  XOR2_X1   g087(.A(G71gat), .B(G78gat), .Z(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n288_), .A2(new_n289_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G231gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT78), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(G15gat), .A2(G22gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G15gat), .A2(G22gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G1gat), .A2(G8gat), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n298_), .A2(new_n299_), .B1(KEYINPUT14), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n297_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n294_), .B(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G127gat), .B(G155gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G183gat), .B(G211gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT17), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n303_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT80), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n308_), .A2(new_n309_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n303_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n285_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G230gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n241_), .A2(new_n235_), .A3(new_n233_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n232_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n240_), .B1(new_n321_), .B2(new_n228_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n292_), .B(new_n258_), .C1(new_n320_), .C2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n292_), .B1(new_n242_), .B2(new_n258_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n319_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT70), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT12), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n323_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n328_), .A2(KEYINPUT12), .ZN(new_n331_));
  INV_X1    g130(.A(new_n292_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n264_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n331_), .ZN(new_n334_));
  AOI211_X1 g133(.A(new_n292_), .B(new_n334_), .C1(new_n242_), .C2(new_n258_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n330_), .B(new_n318_), .C1(new_n333_), .C2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G120gat), .B(G148gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT5), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G176gat), .B(G204gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  OR3_X1    g140(.A1(new_n327_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n341_), .B1(new_n327_), .B2(new_n337_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT13), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n317_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G197gat), .B(G204gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT21), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n347_), .A2(new_n348_), .ZN(new_n352_));
  MUX2_X1   g151(.A(new_n351_), .B(new_n350_), .S(new_n352_), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT95), .ZN(new_n354_));
  OR2_X1    g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G155gat), .B(G162gat), .Z(new_n359_));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT90), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  OR3_X1    g162(.A1(new_n355_), .A2(KEYINPUT91), .A3(KEYINPUT3), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(new_n355_), .B2(KEYINPUT91), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n357_), .A2(KEYINPUT92), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT2), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n359_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n363_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n354_), .B1(KEYINPUT29), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(KEYINPUT93), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n353_), .B(KEYINPUT94), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(KEYINPUT29), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n373_), .ZN(new_n376_));
  OAI22_X1  g175(.A1(new_n371_), .A2(new_n373_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G78gat), .B(G106gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT96), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n377_), .B(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n370_), .A2(KEYINPUT29), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT28), .ZN(new_n382_));
  XOR2_X1   g181(.A(G22gat), .B(G50gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n384_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G71gat), .B(G99gat), .ZN(new_n388_));
  INV_X1    g187(.A(G43gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT88), .B(G15gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OR3_X1    g199(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G183gat), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n403_), .A2(KEYINPUT83), .A3(KEYINPUT25), .ZN(new_n404_));
  INV_X1    g203(.A(G190gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT26), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n404_), .B1(KEYINPUT84), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT25), .B1(new_n403_), .B2(KEYINPUT83), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT26), .B(G190gat), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n407_), .B(new_n408_), .C1(KEYINPUT84), .C2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n396_), .A2(KEYINPUT85), .A3(new_n397_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT23), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(G183gat), .A3(G190gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT86), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT23), .B1(new_n403_), .B2(new_n405_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n402_), .A2(new_n410_), .A3(new_n411_), .A4(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(G176gat), .B1(KEYINPUT87), .B2(KEYINPUT22), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G169gat), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n415_), .A2(new_n413_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n425_), .A2(KEYINPUT89), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(KEYINPUT89), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n394_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n426_), .B2(new_n394_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G127gat), .B(G134gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G113gat), .B(G120gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n432_), .B(KEYINPUT31), .Z(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n429_), .A2(new_n434_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT106), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT22), .B(G169gat), .ZN(new_n440_));
  INV_X1    g239(.A(G176gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n414_), .A2(new_n415_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n397_), .B(new_n442_), .C1(new_n443_), .C2(new_n421_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT99), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT25), .B(G183gat), .Z(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT98), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n409_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n420_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n449_), .A2(new_n398_), .A3(new_n401_), .A4(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n446_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n353_), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n453_), .B(KEYINPUT100), .Z(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT20), .B1(new_n374_), .B2(new_n423_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G226gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT19), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n452_), .A2(new_n353_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n374_), .B2(new_n423_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n462_), .A2(KEYINPUT97), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(KEYINPUT97), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n460_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n457_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n459_), .A2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G8gat), .B(G36gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(G64gat), .B(G92gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT32), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n439_), .B1(new_n468_), .B2(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n459_), .A2(KEYINPUT106), .A3(new_n467_), .A4(new_n474_), .ZN(new_n477_));
  AOI211_X1 g276(.A(KEYINPUT4), .B(new_n432_), .C1(new_n363_), .C2(new_n369_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n370_), .B(new_n432_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(KEYINPUT4), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G225gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT102), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n480_), .A2(new_n482_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G1gat), .B(G29gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G85gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT0), .B(G57gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n354_), .A2(new_n451_), .A3(new_n444_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n492_), .B(KEYINPUT20), .C1(new_n374_), .C2(new_n423_), .ZN(new_n493_));
  MUX2_X1   g292(.A(new_n493_), .B(new_n465_), .S(new_n466_), .Z(new_n494_));
  AOI21_X1  g293(.A(new_n491_), .B1(new_n494_), .B2(new_n475_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n476_), .A2(new_n477_), .A3(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n459_), .A2(new_n473_), .A3(new_n467_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n473_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n468_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n483_), .A2(KEYINPUT33), .A3(new_n487_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT103), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT104), .B(KEYINPUT33), .Z(new_n502_));
  INV_X1    g301(.A(new_n479_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n503_), .A2(KEYINPUT105), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(KEYINPUT105), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n482_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n487_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n489_), .A2(new_n502_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  AND4_X1   g307(.A1(new_n497_), .A2(new_n499_), .A3(new_n501_), .A4(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n387_), .B(new_n438_), .C1(new_n496_), .C2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n387_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n438_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n437_), .A2(new_n387_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n490_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n499_), .A2(new_n497_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT107), .B(KEYINPUT27), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n494_), .A2(new_n498_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n497_), .A2(new_n518_), .A3(KEYINPUT27), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n510_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n302_), .B(new_n245_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(G229gat), .A3(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n302_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n266_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n302_), .A2(new_n245_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G229gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT81), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n523_), .A2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G113gat), .B(G141gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT82), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n530_), .A2(new_n533_), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n521_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT108), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT108), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n521_), .A2(new_n540_), .A3(new_n537_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n346_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n490_), .B(KEYINPUT109), .Z(new_n544_));
  OR3_X1    g343(.A1(new_n543_), .A2(G1gat), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT38), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n345_), .A2(new_n537_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT110), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n277_), .A2(new_n282_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(new_n316_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n521_), .A3(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(G1gat), .B1(new_n552_), .B2(new_n491_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n545_), .A2(new_n546_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(new_n553_), .A3(new_n554_), .ZN(G1324gat));
  NAND2_X1  g354(.A1(new_n517_), .A2(new_n519_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(G8gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n542_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT111), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT111), .B1(new_n542_), .B2(new_n558_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(G8gat), .B1(new_n552_), .B2(new_n557_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT112), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT39), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n563_), .A2(new_n569_), .A3(KEYINPUT40), .A4(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT40), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n569_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(G1325gat));
  OAI21_X1  g375(.A(G15gat), .B1(new_n552_), .B2(new_n438_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT113), .B(KEYINPUT41), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n438_), .A2(G15gat), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n579_), .B(new_n580_), .C1(new_n543_), .C2(new_n581_), .ZN(G1326gat));
  OAI21_X1  g381(.A(G22gat), .B1(new_n552_), .B2(new_n387_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT42), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n387_), .A2(G22gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n584_), .B1(new_n543_), .B2(new_n585_), .ZN(G1327gat));
  NAND2_X1  g385(.A1(new_n539_), .A2(new_n541_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n550_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(new_n315_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n589_), .A2(new_n345_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(G29gat), .B1(new_n592_), .B2(new_n490_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT44), .ZN(new_n594_));
  INV_X1    g393(.A(new_n285_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n510_), .B2(new_n520_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT43), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n549_), .A2(new_n316_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT43), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n596_), .B(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n601_), .A2(KEYINPUT44), .A3(new_n316_), .A4(new_n549_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n544_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n604_), .A2(G29gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n593_), .B1(new_n603_), .B2(new_n605_), .ZN(G1328gat));
  NAND3_X1  g405(.A1(new_n599_), .A2(new_n602_), .A3(new_n556_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(G36gat), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n557_), .A2(G36gat), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n587_), .A2(new_n590_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT45), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT46), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n608_), .A2(new_n611_), .A3(KEYINPUT46), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1329gat));
  NAND4_X1  g415(.A1(new_n599_), .A2(new_n602_), .A3(G43gat), .A4(new_n437_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n389_), .B1(new_n591_), .B2(new_n438_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g419(.A(G50gat), .B1(new_n592_), .B2(new_n511_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n511_), .A2(G50gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n603_), .B2(new_n622_), .ZN(G1331gat));
  NOR2_X1   g422(.A1(new_n345_), .A2(new_n537_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n521_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(new_n551_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G57gat), .B1(new_n627_), .B2(new_n491_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n625_), .A2(new_n317_), .ZN(new_n629_));
  INV_X1    g428(.A(G57gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n604_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(G1332gat));
  INV_X1    g431(.A(G64gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n626_), .B2(new_n556_), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n629_), .A2(new_n633_), .A3(new_n556_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1333gat));
  INV_X1    g437(.A(G71gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n626_), .B2(new_n437_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT49), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n629_), .A2(new_n639_), .A3(new_n437_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1334gat));
  NOR2_X1   g442(.A1(new_n387_), .A2(G78gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT115), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n629_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n626_), .A2(new_n511_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT50), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n647_), .A2(new_n648_), .A3(G78gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n647_), .B2(G78gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT116), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(G1335gat));
  AND2_X1   g452(.A1(new_n625_), .A2(new_n589_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G85gat), .B1(new_n654_), .B2(new_n604_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n624_), .A2(new_n316_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n597_), .A2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n490_), .A2(new_n249_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(G1336gat));
  AOI21_X1  g458(.A(G92gat), .B1(new_n654_), .B2(new_n556_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n556_), .A2(new_n250_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n657_), .B2(new_n661_), .ZN(G1337gat));
  AOI21_X1  g461(.A(new_n224_), .B1(new_n657_), .B2(new_n437_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n437_), .A2(new_n246_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n654_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT51), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(G1338gat));
  NAND3_X1  g466(.A1(new_n654_), .A2(new_n225_), .A3(new_n511_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n601_), .A2(new_n511_), .A3(new_n316_), .A4(new_n624_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT52), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(new_n670_), .A3(G106gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(G106gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT53), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT53), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n675_), .B(new_n668_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1339gat));
  NOR2_X1   g476(.A1(new_n556_), .A2(new_n544_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n513_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n330_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n319_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(KEYINPUT55), .A3(new_n336_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n333_), .A2(new_n335_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT55), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n318_), .A4(new_n330_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT117), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT117), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n683_), .A2(new_n689_), .A3(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT56), .B1(new_n691_), .B2(new_n341_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n683_), .A2(new_n689_), .A3(new_n686_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n689_), .B1(new_n683_), .B2(new_n686_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT56), .B(new_n341_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n537_), .B(new_n342_), .C1(new_n692_), .C2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n528_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n525_), .A2(new_n526_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n533_), .B1(new_n522_), .B2(new_n528_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n530_), .A2(new_n533_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n344_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n550_), .B1(new_n697_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n342_), .A2(new_n701_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT58), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n595_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n341_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT56), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n704_), .B1(new_n711_), .B2(new_n695_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT58), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n703_), .A2(KEYINPUT57), .B1(new_n708_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n537_), .A2(new_n342_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n711_), .B2(new_n695_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n702_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n588_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT118), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT118), .B(new_n588_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n714_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n316_), .ZN(new_n725_));
  OR3_X1    g524(.A1(new_n346_), .A2(KEYINPUT54), .A3(new_n537_), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT54), .B1(new_n346_), .B2(new_n537_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n680_), .B1(new_n725_), .B2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G113gat), .B1(new_n729_), .B2(new_n537_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(KEYINPUT120), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT121), .B1(new_n724_), .B2(new_n316_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT121), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n733_), .B(new_n315_), .C1(new_n714_), .C2(new_n723_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n728_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n680_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT59), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n735_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n315_), .B1(new_n714_), .B2(new_n723_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n728_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n736_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT59), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n740_), .A2(G113gat), .A3(new_n537_), .A4(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n730_), .A2(KEYINPUT120), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n731_), .A2(new_n745_), .A3(new_n746_), .ZN(G1340gat));
  INV_X1    g546(.A(KEYINPUT123), .ZN(new_n748_));
  INV_X1    g547(.A(G120gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n345_), .B1(new_n743_), .B2(KEYINPUT59), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n740_), .B2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n345_), .A2(KEYINPUT60), .ZN(new_n752_));
  MUX2_X1   g551(.A(KEYINPUT60), .B(new_n752_), .S(new_n749_), .Z(new_n753_));
  OAI211_X1 g552(.A(new_n736_), .B(new_n753_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT122), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n748_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n713_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n285_), .B1(new_n712_), .B2(KEYINPUT58), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n757_), .A2(new_n758_), .B1(new_n718_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n722_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n721_), .B2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n733_), .B1(new_n763_), .B2(new_n315_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n741_), .A2(KEYINPUT121), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n738_), .B1(new_n766_), .B2(new_n728_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n345_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n729_), .B2(new_n737_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G120gat), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT122), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n754_), .B(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(KEYINPUT123), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n756_), .A2(new_n773_), .ZN(G1341gat));
  NAND2_X1  g573(.A1(new_n740_), .A2(new_n744_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G127gat), .B1(new_n775_), .B2(new_n316_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n316_), .A2(G127gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n743_), .B2(new_n777_), .ZN(G1342gat));
  OAI21_X1  g577(.A(G134gat), .B1(new_n775_), .B2(new_n595_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n588_), .A2(G134gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n743_), .B2(new_n780_), .ZN(G1343gat));
  NOR2_X1   g580(.A1(new_n741_), .A2(new_n742_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(new_n512_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n678_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n537_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(KEYINPUT124), .B(G141gat), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(G1344gat));
  NOR2_X1   g587(.A1(new_n784_), .A2(new_n345_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT125), .B(G148gat), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1345gat));
  NOR2_X1   g590(.A1(new_n784_), .A2(new_n316_), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT61), .B(G155gat), .Z(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1346gat));
  OAI21_X1  g593(.A(G162gat), .B1(new_n784_), .B2(new_n595_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n588_), .A2(G162gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n784_), .B2(new_n796_), .ZN(G1347gat));
  NOR2_X1   g596(.A1(new_n557_), .A2(new_n604_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n735_), .A2(new_n679_), .A3(new_n537_), .A4(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G169gat), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT62), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n742_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n798_), .A2(new_n679_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n440_), .A3(new_n537_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n799_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n802_), .A2(new_n806_), .A3(new_n807_), .ZN(G1348gat));
  AOI21_X1  g607(.A(G176gat), .B1(new_n805_), .B2(new_n768_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n782_), .A2(new_n511_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n798_), .A2(new_n437_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n811_), .A2(new_n441_), .A3(new_n345_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n809_), .B1(new_n810_), .B2(new_n812_), .ZN(G1349gat));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n316_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G183gat), .B1(new_n816_), .B2(KEYINPUT126), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT126), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n316_), .A2(new_n448_), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n817_), .A2(new_n819_), .B1(new_n805_), .B2(new_n820_), .ZN(G1350gat));
  NAND3_X1  g620(.A1(new_n805_), .A2(new_n409_), .A3(new_n550_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n803_), .A2(new_n595_), .A3(new_n804_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n405_), .ZN(G1351gat));
  NOR2_X1   g623(.A1(new_n557_), .A2(new_n490_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n783_), .A2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n785_), .ZN(new_n827_));
  INV_X1    g626(.A(G197gat), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(G1352gat));
  INV_X1    g628(.A(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n768_), .A3(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT127), .B(G204gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n826_), .B2(new_n345_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1353gat));
  XOR2_X1   g634(.A(KEYINPUT63), .B(G211gat), .Z(new_n836_));
  NAND3_X1  g635(.A1(new_n830_), .A2(new_n315_), .A3(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n826_), .B2(new_n316_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1354gat));
  OAI21_X1  g639(.A(G218gat), .B1(new_n826_), .B2(new_n595_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n588_), .A2(G218gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n826_), .B2(new_n842_), .ZN(G1355gat));
endmodule


