//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_;
  INV_X1    g000(.A(G134gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G127gat), .ZN(new_n203_));
  INV_X1    g002(.A(G127gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G134gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G120gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G113gat), .ZN(new_n208_));
  INV_X1    g007(.A(G113gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G120gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n203_), .A2(new_n205_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G227gat), .A2(G233gat), .ZN(new_n215_));
  INV_X1    g014(.A(G15gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G71gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n215_), .B(G15gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(G71gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(G99gat), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT81), .B(G43gat), .Z(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(G71gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n217_), .A2(new_n218_), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n222_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n224_), .B1(new_n222_), .B2(new_n228_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT25), .B(G183gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G169gat), .ZN(new_n240_));
  INV_X1    g039(.A(G176gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n242_), .A2(KEYINPUT24), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G169gat), .A2(G176gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(KEYINPUT24), .A3(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n234_), .A2(new_n239_), .A3(new_n243_), .A4(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(G183gat), .A2(G190gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n237_), .A2(new_n247_), .A3(new_n238_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n244_), .ZN(new_n249_));
  AND2_X1   g048(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G169gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n249_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n248_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n240_), .A2(KEYINPUT22), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT22), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G169gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n257_), .A2(new_n258_), .A3(new_n260_), .A4(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n244_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(KEYINPUT80), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT30), .B(new_n246_), .C1(new_n256_), .C2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(KEYINPUT80), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n254_), .A2(new_n255_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n248_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT30), .B1(new_n269_), .B2(new_n246_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT82), .B1(new_n266_), .B2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n246_), .B1(new_n256_), .B2(new_n264_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT30), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT82), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n265_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n231_), .B1(new_n271_), .B2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n276_), .A2(new_n231_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT31), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n231_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n274_), .A2(new_n275_), .A3(new_n265_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n275_), .B1(new_n274_), .B2(new_n265_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n276_), .A2(new_n231_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT83), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n279_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n279_), .B2(new_n286_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n214_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n277_), .A2(new_n278_), .A3(KEYINPUT31), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n284_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT83), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n212_), .A2(new_n213_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n279_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n297_));
  INV_X1    g096(.A(G141gat), .ZN(new_n298_));
  INV_X1    g097(.A(G148gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n300_), .A2(new_n303_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(KEYINPUT1), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT1), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(G155gat), .A3(G162gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n313_), .A3(new_n307_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G141gat), .B(G148gat), .Z(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n294_), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n306_), .A2(new_n309_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n214_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n320_), .A3(KEYINPUT92), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT92), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n322_), .A3(new_n214_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(KEYINPUT4), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G1gat), .B(G29gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT93), .B(G85gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT0), .B(G57gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n329_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n330_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n335_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n328_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n336_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n290_), .A2(new_n296_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n319_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT84), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G22gat), .B(G50gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT28), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n347_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT86), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(KEYINPUT21), .ZN(new_n352_));
  INV_X1    g151(.A(G197gat), .ZN(new_n353_));
  INV_X1    g152(.A(G204gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT85), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT85), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G204gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n353_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(G197gat), .A2(G204gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n352_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(KEYINPUT86), .A2(G197gat), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n362_));
  AOI21_X1  g161(.A(G204gat), .B1(new_n353_), .B2(KEYINPUT86), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT21), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G211gat), .B(G218gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n367_), .A2(KEYINPUT21), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n358_), .A2(new_n359_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT87), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n366_), .A2(new_n370_), .A3(KEYINPUT87), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G228gat), .A2(G233gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n319_), .B2(new_n345_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n363_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT85), .B(G204gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n361_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n367_), .B1(new_n383_), .B2(KEYINPUT21), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n384_), .A2(new_n360_), .B1(new_n369_), .B2(new_n368_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n319_), .A2(new_n345_), .ZN(new_n386_));
  OAI211_X1 g185(.A(G228gat), .B(G233gat), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n378_), .A2(new_n380_), .A3(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n366_), .A2(KEYINPUT87), .A3(new_n370_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT87), .B1(new_n366_), .B2(new_n370_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n376_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n386_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n375_), .B1(new_n392_), .B2(new_n371_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n379_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  AND4_X1   g193(.A1(KEYINPUT88), .A2(new_n350_), .A3(new_n388_), .A4(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT88), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n388_), .A2(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n397_), .A2(new_n350_), .B1(new_n394_), .B2(new_n388_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n373_), .A2(new_n374_), .A3(new_n272_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT89), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n244_), .B(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n262_), .A3(new_n248_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n404_), .A2(new_n262_), .A3(new_n248_), .A4(KEYINPUT90), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n246_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT91), .B1(new_n371_), .B2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n407_), .A2(new_n246_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT91), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n411_), .A2(new_n385_), .A3(new_n412_), .A4(new_n408_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n402_), .A2(KEYINPUT20), .A3(new_n410_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G226gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT19), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n414_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G8gat), .B(G36gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT18), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(new_n421_), .Z(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n272_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT20), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n371_), .B2(new_n409_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n416_), .A3(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n418_), .A2(new_n423_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n423_), .B1(new_n418_), .B2(new_n428_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n401_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n389_), .A2(new_n390_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n426_), .B1(new_n432_), .B2(new_n272_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n413_), .A2(new_n410_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n416_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n425_), .A2(new_n416_), .A3(new_n427_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n422_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n246_), .A2(new_n405_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT95), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT95), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n246_), .A2(new_n440_), .A3(new_n405_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n385_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n402_), .A2(KEYINPUT20), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n416_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n425_), .A2(new_n417_), .A3(new_n427_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n423_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n437_), .A2(new_n447_), .A3(KEYINPUT27), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n400_), .A2(new_n431_), .A3(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n344_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT94), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n436_), .B1(new_n417_), .B2(new_n414_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n422_), .A2(KEYINPUT32), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n451_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n446_), .A2(new_n454_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n456_));
  OAI211_X1 g255(.A(KEYINPUT94), .B(new_n453_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n328_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n459_));
  AOI211_X1 g258(.A(new_n335_), .B(new_n459_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT33), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n461_), .B2(new_n338_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n330_), .A2(KEYINPUT33), .A3(new_n335_), .A4(new_n337_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n418_), .A2(new_n423_), .A3(new_n428_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n437_), .A4(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n458_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n400_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n431_), .A2(new_n448_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n399_), .A2(new_n343_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT96), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n395_), .A2(new_n342_), .A3(new_n398_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT96), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n471_), .A2(new_n431_), .A3(new_n472_), .A4(new_n448_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n290_), .A2(new_n296_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n450_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT68), .ZN(new_n477_));
  NOR2_X1   g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n480_), .B2(KEYINPUT9), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT65), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(new_n479_), .ZN(new_n484_));
  AND2_X1   g283(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n485_));
  NOR2_X1   g284(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n482_), .B(new_n479_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n481_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G106gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT6), .B1(new_n227_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(G99gat), .A3(G106gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT10), .B(G99gat), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n490_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n489_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n500_));
  XOR2_X1   g299(.A(G71gat), .B(G78gat), .Z(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n500_), .A2(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT8), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n494_), .A2(KEYINPUT66), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT66), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n491_), .A2(new_n507_), .A3(new_n493_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT7), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n480_), .A2(new_n478_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n505_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n505_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n514_), .B1(new_n494_), .B2(new_n510_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n497_), .B(new_n504_), .C1(new_n513_), .C2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT67), .ZN(new_n517_));
  INV_X1    g316(.A(G230gat), .ZN(new_n518_));
  INV_X1    g317(.A(G233gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n497_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT12), .ZN(new_n524_));
  INV_X1    g323(.A(new_n504_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n524_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n522_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n517_), .B1(new_n516_), .B2(new_n521_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n477_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n523_), .A2(new_n525_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n516_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n520_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(KEYINPUT12), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n529_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n536_), .A2(KEYINPUT68), .A3(new_n537_), .A4(new_n522_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n530_), .A2(new_n533_), .A3(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G120gat), .B(G148gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G176gat), .B(G204gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n530_), .A2(new_n533_), .A3(new_n538_), .A4(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n548_), .A2(KEYINPUT13), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(KEYINPUT13), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G169gat), .B(G197gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n552_), .B(new_n553_), .Z(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G15gat), .B(G22gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G1gat), .A2(G8gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT14), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G1gat), .B(G8gat), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n560_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G43gat), .B(G50gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G29gat), .B(G36gat), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT70), .ZN(new_n567_));
  INV_X1    g366(.A(G36gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(G29gat), .ZN(new_n569_));
  INV_X1    g368(.A(G29gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(G36gat), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n569_), .A2(new_n571_), .A3(KEYINPUT70), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n565_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n571_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT70), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n566_), .A2(KEYINPUT70), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n564_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n573_), .A2(KEYINPUT15), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT15), .B1(new_n573_), .B2(new_n578_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n563_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n561_), .A2(new_n573_), .A3(new_n562_), .A4(new_n578_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT77), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n582_), .A2(KEYINPUT77), .A3(new_n583_), .A4(new_n584_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n573_), .A2(new_n578_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n563_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n584_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n583_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT76), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT76), .ZN(new_n595_));
  AOI211_X1 g394(.A(new_n595_), .B(new_n583_), .C1(new_n591_), .C2(new_n584_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n589_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n555_), .B1(new_n588_), .B2(new_n597_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n594_), .A2(new_n596_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n599_), .A2(new_n587_), .A3(new_n589_), .A4(new_n554_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT78), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT78), .B(new_n555_), .C1(new_n588_), .C2(new_n597_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n476_), .A2(new_n551_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT34), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT35), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(KEYINPUT72), .ZN(new_n611_));
  OR3_X1    g410(.A1(new_n523_), .A2(KEYINPUT71), .A3(new_n590_), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT71), .B1(new_n523_), .B2(new_n590_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n580_), .A2(new_n581_), .ZN(new_n615_));
  AOI22_X1  g414(.A1(new_n615_), .A2(new_n523_), .B1(new_n609_), .B2(new_n608_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n611_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n610_), .A2(KEYINPUT72), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT73), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G134gat), .B(G162gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT36), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT74), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n614_), .A2(KEYINPUT72), .A3(new_n610_), .A4(new_n616_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n620_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n624_), .A2(KEYINPUT36), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n620_), .B2(new_n627_), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT37), .B1(new_n628_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n620_), .A2(new_n627_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n629_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT37), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n620_), .A2(new_n627_), .A3(new_n625_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n504_), .B(new_n563_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(G127gat), .B(G155gat), .Z(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT16), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT17), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n642_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n646_), .A2(new_n647_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(new_n642_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT75), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n639_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n605_), .A2(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(G1gat), .A3(new_n343_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT97), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT38), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(KEYINPUT38), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n474_), .A2(new_n475_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n450_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n634_), .A2(new_n636_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT98), .Z(new_n663_));
  AND2_X1   g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n551_), .A2(new_n604_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n652_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n664_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G1gat), .B1(new_n669_), .B2(new_n343_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n657_), .A2(new_n658_), .A3(new_n670_), .ZN(G1324gat));
  INV_X1    g470(.A(new_n468_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n654_), .A2(G8gat), .A3(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n664_), .A2(new_n468_), .A3(new_n668_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(G8gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n675_), .B1(new_n674_), .B2(G8gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT39), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n678_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT39), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(new_n681_), .A3(new_n676_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n673_), .B1(new_n679_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n683_), .B(new_n685_), .ZN(G1325gat));
  INV_X1    g485(.A(new_n669_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n475_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n689_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT41), .B1(new_n689_), .B2(G15gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n216_), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n690_), .A2(new_n691_), .B1(new_n654_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n687_), .A2(new_n399_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(G22gat), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n696_), .B2(G22gat), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n400_), .A2(G22gat), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT103), .Z(new_n701_));
  OAI22_X1  g500(.A1(new_n698_), .A2(new_n699_), .B1(new_n654_), .B2(new_n701_), .ZN(G1327gat));
  NOR2_X1   g501(.A1(new_n666_), .A2(new_n662_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n661_), .A2(new_n703_), .A3(new_n665_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n570_), .A3(new_n342_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n476_), .B2(new_n638_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n471_), .A2(new_n431_), .A3(new_n448_), .ZN(new_n710_));
  AOI22_X1  g509(.A1(new_n400_), .A2(new_n466_), .B1(new_n710_), .B2(KEYINPUT96), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n688_), .B1(new_n711_), .B2(new_n473_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n709_), .B(new_n639_), .C1(new_n712_), .C2(new_n450_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n708_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n665_), .A2(new_n652_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n707_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n708_), .A2(new_n713_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n717_), .A2(KEYINPUT44), .A3(new_n652_), .A4(new_n665_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n342_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n721_), .A2(KEYINPUT104), .A3(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT104), .B1(new_n721_), .B2(G29gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n706_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  OAI21_X1  g523(.A(G36gat), .B1(new_n719_), .B2(new_n672_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n672_), .A2(G36gat), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n704_), .A2(KEYINPUT105), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT105), .B1(new_n704_), .B2(new_n727_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(KEYINPUT45), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT45), .B1(new_n728_), .B2(new_n729_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT106), .B1(new_n725_), .B2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(KEYINPUT46), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT106), .B(new_n735_), .C1(new_n725_), .C2(new_n732_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1329gat));
  AOI21_X1  g536(.A(G43gat), .B1(new_n705_), .B2(new_n688_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT107), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n688_), .A2(G43gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n719_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g541(.A(G50gat), .B1(new_n705_), .B2(new_n399_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n399_), .A2(G50gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n720_), .B2(new_n744_), .ZN(G1331gat));
  NAND4_X1  g544(.A1(new_n664_), .A2(new_n666_), .A3(new_n551_), .A4(new_n604_), .ZN(new_n746_));
  INV_X1    g545(.A(G57gat), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n343_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT108), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(KEYINPUT108), .ZN(new_n751_));
  INV_X1    g550(.A(new_n551_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n602_), .A2(new_n603_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n476_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n653_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G57gat), .B1(new_n756_), .B2(new_n342_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n750_), .A2(new_n751_), .A3(new_n757_), .ZN(G1332gat));
  OAI21_X1  g557(.A(G64gat), .B1(new_n746_), .B2(new_n672_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT48), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n672_), .A2(G64gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n755_), .B2(new_n761_), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n746_), .B2(new_n475_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT49), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n756_), .A2(new_n218_), .A3(new_n688_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1334gat));
  OAI21_X1  g565(.A(G78gat), .B1(new_n746_), .B2(new_n400_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT50), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n400_), .A2(G78gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n755_), .B2(new_n769_), .ZN(G1335gat));
  AND2_X1   g569(.A1(new_n754_), .A2(new_n703_), .ZN(new_n771_));
  AOI21_X1  g570(.A(G85gat), .B1(new_n771_), .B2(new_n342_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT109), .Z(new_n773_));
  AND3_X1   g572(.A1(new_n708_), .A2(new_n713_), .A3(KEYINPUT110), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT110), .B1(new_n708_), .B2(new_n713_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n666_), .A2(new_n753_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n551_), .A2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(G85gat), .A3(new_n342_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n773_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT111), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n773_), .A2(new_n783_), .A3(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1336gat));
  INV_X1    g584(.A(G92gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n779_), .B2(new_n468_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n771_), .A2(new_n786_), .A3(new_n468_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1337gat));
  INV_X1    g588(.A(new_n778_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n688_), .B(new_n790_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G99gat), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n771_), .A2(new_n495_), .A3(new_n688_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n795_), .A2(KEYINPUT113), .A3(KEYINPUT51), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n793_), .B1(G99gat), .B2(new_n791_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n795_), .B2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT51), .B1(new_n798_), .B2(KEYINPUT113), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT114), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n792_), .A2(KEYINPUT113), .A3(new_n794_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n792_), .A2(new_n794_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT112), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n804_), .A2(new_n806_), .A3(new_n807_), .A4(new_n797_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n801_), .A2(new_n808_), .ZN(G1338gat));
  NAND2_X1  g608(.A1(new_n790_), .A2(new_n399_), .ZN(new_n810_));
  OAI21_X1  g609(.A(G106gat), .B1(new_n714_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT52), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n771_), .A2(new_n490_), .A3(new_n399_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g614(.A1(new_n475_), .A2(new_n449_), .A3(new_n343_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT116), .B1(new_n753_), .B2(new_n547_), .ZN(new_n819_));
  AND4_X1   g618(.A1(KEYINPUT116), .A2(new_n547_), .A3(new_n603_), .A4(new_n602_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n530_), .A2(new_n822_), .A3(new_n538_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n536_), .A2(KEYINPUT55), .A3(new_n537_), .A4(new_n522_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n516_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n520_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n545_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n828_), .A2(KEYINPUT56), .A3(new_n545_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n582_), .A2(new_n593_), .A3(new_n584_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n554_), .B1(new_n592_), .B2(new_n583_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n600_), .A2(new_n836_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n821_), .A2(new_n833_), .B1(new_n548_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n662_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n818_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n820_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842_));
  INV_X1    g641(.A(new_n547_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n604_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT56), .B1(new_n828_), .B2(new_n545_), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n830_), .B(new_n544_), .C1(new_n823_), .C2(new_n827_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n841_), .B(new_n844_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n548_), .A2(new_n837_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(KEYINPUT57), .A3(new_n662_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n547_), .A2(new_n837_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n639_), .B(new_n851_), .C1(new_n853_), .C2(KEYINPUT58), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(KEYINPUT58), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n852_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n851_), .B1(new_n860_), .B2(new_n639_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n840_), .B(new_n850_), .C1(new_n856_), .C2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT118), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n639_), .B1(new_n853_), .B2(KEYINPUT58), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT117), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n855_), .A3(new_n854_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n840_), .A4(new_n850_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n863_), .A2(new_n652_), .A3(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n652_), .A2(new_n753_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT115), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n638_), .A3(new_n752_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(KEYINPUT54), .Z(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n817_), .B1(new_n869_), .B2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n209_), .A3(new_n753_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n817_), .A2(KEYINPUT59), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n862_), .A2(new_n652_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n873_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n753_), .B(new_n879_), .C1(new_n875_), .C2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n876_), .B1(new_n882_), .B2(new_n209_), .ZN(G1340gat));
  OAI21_X1  g682(.A(new_n207_), .B1(new_n752_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n875_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n207_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n551_), .B(new_n879_), .C1(new_n875_), .C2(new_n880_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n887_), .B2(new_n207_), .ZN(G1341gat));
  AOI21_X1  g687(.A(new_n666_), .B1(new_n862_), .B2(KEYINPUT118), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n873_), .B1(new_n889_), .B2(new_n868_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n890_), .A2(new_n652_), .A3(new_n817_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT119), .B1(new_n891_), .B2(G127gat), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n869_), .A2(new_n874_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n816_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n893_), .B(new_n204_), .C1(new_n895_), .C2(new_n652_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n878_), .A2(new_n873_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n895_), .A2(KEYINPUT59), .B1(new_n897_), .B2(new_n877_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n652_), .A2(new_n204_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n892_), .A2(new_n896_), .B1(new_n898_), .B2(new_n899_), .ZN(G1342gat));
  OR3_X1    g699(.A1(new_n895_), .A2(G134gat), .A3(new_n663_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n639_), .B(new_n879_), .C1(new_n875_), .C2(new_n880_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n903_), .B2(new_n202_), .ZN(G1343gat));
  NAND4_X1  g703(.A1(new_n475_), .A2(new_n672_), .A3(new_n399_), .A4(new_n342_), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(KEYINPUT120), .Z(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n869_), .B2(new_n874_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n753_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n551_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT121), .B(G148gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1345gat));
  XNOR2_X1  g712(.A(KEYINPUT61), .B(G155gat), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n908_), .B2(new_n666_), .ZN(new_n917_));
  NOR4_X1   g716(.A1(new_n890_), .A2(KEYINPUT122), .A3(new_n652_), .A4(new_n907_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n915_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n894_), .A2(new_n666_), .A3(new_n906_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT122), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n908_), .A2(new_n916_), .A3(new_n666_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n921_), .A2(new_n922_), .A3(new_n914_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n919_), .A2(new_n923_), .ZN(G1346gat));
  INV_X1    g723(.A(new_n908_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G162gat), .B1(new_n925_), .B2(new_n638_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n663_), .A2(G162gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n925_), .B2(new_n927_), .ZN(G1347gat));
  INV_X1    g727(.A(new_n344_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n468_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n399_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n753_), .B(new_n931_), .C1(new_n878_), .C2(new_n873_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n240_), .B1(new_n933_), .B2(KEYINPUT62), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n935_), .A2(KEYINPUT123), .A3(new_n936_), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n932_), .B(new_n934_), .C1(new_n933_), .C2(KEYINPUT62), .ZN(new_n938_));
  INV_X1    g737(.A(new_n253_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n937_), .B(new_n938_), .C1(new_n939_), .C2(new_n932_), .ZN(G1348gat));
  NAND3_X1  g739(.A1(new_n897_), .A2(new_n551_), .A3(new_n931_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n890_), .A2(new_n399_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n752_), .A2(new_n930_), .A3(new_n241_), .ZN(new_n943_));
  AOI22_X1  g742(.A1(new_n941_), .A2(new_n252_), .B1(new_n942_), .B2(new_n943_), .ZN(G1349gat));
  NAND2_X1  g743(.A1(new_n897_), .A2(new_n931_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n945_), .A2(new_n652_), .A3(new_n232_), .ZN(new_n946_));
  INV_X1    g745(.A(G183gat), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n942_), .A2(new_n666_), .A3(new_n468_), .A4(new_n929_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n946_), .B1(new_n947_), .B2(new_n948_), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n945_), .B2(new_n638_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n233_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n663_), .A2(new_n951_), .ZN(new_n952_));
  XOR2_X1   g751(.A(new_n952_), .B(KEYINPUT124), .Z(new_n953_));
  OAI21_X1  g752(.A(new_n950_), .B1(new_n945_), .B2(new_n953_), .ZN(G1351gat));
  NOR3_X1   g753(.A1(new_n688_), .A2(new_n672_), .A3(new_n469_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n894_), .A2(new_n955_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n956_), .A2(new_n604_), .A3(new_n957_), .ZN(new_n958_));
  AND2_X1   g757(.A1(new_n894_), .A2(new_n955_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(new_n753_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(KEYINPUT125), .B(G197gat), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n958_), .B1(new_n960_), .B2(new_n961_), .ZN(G1352gat));
  AOI21_X1  g761(.A(G204gat), .B1(new_n959_), .B2(new_n551_), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n956_), .A2(new_n382_), .A3(new_n752_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1353gat));
  AOI21_X1  g764(.A(new_n652_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n959_), .A2(new_n966_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n968_));
  XOR2_X1   g767(.A(new_n968_), .B(KEYINPUT126), .Z(new_n969_));
  XOR2_X1   g768(.A(new_n969_), .B(KEYINPUT127), .Z(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n967_), .A2(new_n971_), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n959_), .A2(new_n966_), .A3(new_n970_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(G1354gat));
  OAI21_X1  g773(.A(G218gat), .B1(new_n956_), .B2(new_n638_), .ZN(new_n975_));
  OR2_X1    g774(.A1(new_n663_), .A2(G218gat), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n975_), .B1(new_n956_), .B2(new_n976_), .ZN(G1355gat));
endmodule


