//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n959_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n980_, new_n981_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n989_, new_n990_, new_n992_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1003_, new_n1004_, new_n1005_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT20), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n207_), .B(KEYINPUT92), .Z(new_n208_));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209_));
  AND2_X1   g008(.A1(new_n209_), .A2(KEYINPUT21), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n209_), .B1(new_n212_), .B2(new_n207_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n207_), .A2(new_n212_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT91), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT91), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n207_), .A2(new_n216_), .A3(new_n212_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n213_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT80), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT82), .B(G176gat), .Z(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT22), .B(G169gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G183gat), .A3(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(G183gat), .B2(G190gat), .ZN(new_n229_));
  OAI22_X1  g028(.A1(new_n228_), .A2(new_n229_), .B1(G183gat), .B2(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT25), .B(G183gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OR3_X1    g033(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n234_), .B(new_n235_), .C1(new_n222_), .C2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n229_), .A2(KEYINPUT81), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n229_), .A2(KEYINPUT81), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n228_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n231_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n206_), .B1(new_n219_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G226gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT19), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G183gat), .A2(G190gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n225_), .B1(new_n240_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G183gat), .ZN(new_n248_));
  INV_X1    g047(.A(G190gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT23), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n236_), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n250_), .A2(new_n227_), .B1(new_n251_), .B2(new_n220_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT95), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT95), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n252_), .A2(new_n255_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n247_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n242_), .B(new_n245_), .C1(new_n219_), .C2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n214_), .B(KEYINPUT91), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n259_), .A2(new_n213_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n237_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n238_), .A2(new_n239_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n227_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n261_), .A2(new_n263_), .B1(new_n230_), .B2(new_n225_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n206_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n257_), .A2(new_n219_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n205_), .B(new_n258_), .C1(new_n267_), .C2(new_n245_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT99), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n260_), .A2(new_n247_), .A3(new_n253_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n242_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n244_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(new_n245_), .A3(new_n266_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n205_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n269_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  AOI211_X1 g075(.A(KEYINPUT99), .B(new_n205_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n277_));
  OAI211_X1 g076(.A(KEYINPUT27), .B(new_n268_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(KEYINPUT20), .B(new_n245_), .C1(new_n260_), .C2(new_n264_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n257_), .A2(new_n219_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n245_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n275_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n268_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT27), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(KEYINPUT1), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n289_), .B2(KEYINPUT1), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT86), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n288_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n291_), .B2(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n293_), .A2(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n287_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT88), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  OAI22_X1  g104(.A1(KEYINPUT87), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n299_), .A2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n308_), .B(new_n310_), .C1(KEYINPUT2), .C2(new_n298_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n305_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n301_), .A2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G127gat), .B(G134gat), .Z(new_n314_));
  XOR2_X1   g113(.A(G113gat), .B(G120gat), .Z(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n293_), .A2(new_n300_), .B1(new_n305_), .B2(new_n311_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n316_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n320_), .A3(KEYINPUT4), .ZN(new_n321_));
  OR3_X1    g120(.A1(new_n318_), .A2(new_n319_), .A3(KEYINPUT4), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT96), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G57gat), .B(G85gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n325_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n326_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n331_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n325_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n337_), .B2(new_n332_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n278_), .A2(new_n286_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n219_), .B1(new_n318_), .B2(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(KEYINPUT90), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(KEYINPUT90), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(G228gat), .A4(G233gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n346_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G228gat), .A2(G233gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G22gat), .B(G50gat), .Z(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n301_), .A2(new_n343_), .A3(new_n312_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT28), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT28), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n318_), .A2(new_n355_), .A3(new_n343_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT89), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n352_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n356_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT89), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n351_), .A3(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT93), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT94), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n360_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n366_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n347_), .B(new_n350_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n316_), .B(KEYINPUT31), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374_));
  INV_X1    g173(.A(G15gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G71gat), .ZN(new_n377_));
  INV_X1    g176(.A(G99gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT83), .B(G43gat), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n379_), .B(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n264_), .A2(KEYINPUT30), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n241_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT84), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(new_n388_), .A3(new_n385_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n382_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n382_), .A2(new_n389_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n373_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n382_), .A2(new_n389_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n387_), .A2(new_n389_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n393_), .B(new_n372_), .C1(new_n394_), .C2(new_n382_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n358_), .A2(new_n359_), .A3(new_n352_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n351_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n367_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n350_), .A2(new_n347_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n360_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n371_), .A2(new_n396_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n396_), .B1(new_n371_), .B2(new_n402_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n342_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n326_), .A2(new_n333_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT33), .B1(new_n406_), .B2(new_n335_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n317_), .A2(new_n320_), .A3(new_n325_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n331_), .B(new_n408_), .C1(new_n323_), .C2(new_n325_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n268_), .A2(new_n283_), .A3(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n407_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT98), .B1(new_n338_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT98), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n406_), .A2(new_n414_), .A3(KEYINPUT33), .A4(new_n335_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n281_), .A2(new_n282_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n339_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n392_), .A2(new_n395_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n400_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(new_n424_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n405_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT69), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT65), .ZN(new_n431_));
  AND2_X1   g230(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(G85gat), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(G85gat), .A2(G92gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT9), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G99gat), .A2(G106gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT10), .B(G99gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G106gat), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n444_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n431_), .B1(new_n439_), .B2(new_n448_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n434_), .A2(new_n435_), .B1(KEYINPUT9), .B2(new_n437_), .ZN(new_n450_));
  AND3_X1   g249(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n453_), .B1(G106gat), .B2(new_n445_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n450_), .A2(new_n454_), .A3(KEYINPUT65), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT8), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT67), .B1(new_n451_), .B2(new_n452_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n442_), .A2(new_n458_), .A3(new_n443_), .ZN(new_n459_));
  AND2_X1   g258(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n460_));
  NOR2_X1   g259(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n461_));
  OAI22_X1  g260(.A1(new_n460_), .A2(new_n461_), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n378_), .A3(new_n447_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n457_), .A2(new_n459_), .A3(new_n462_), .A4(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n437_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n456_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n456_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n462_), .A2(new_n464_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n469_), .B1(new_n470_), .B2(new_n453_), .ZN(new_n471_));
  OAI22_X1  g270(.A1(new_n449_), .A2(new_n455_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G57gat), .B(G64gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G71gat), .B(G78gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(KEYINPUT11), .ZN(new_n475_));
  XOR2_X1   g274(.A(G71gat), .B(G78gat), .Z(new_n476_));
  INV_X1    g275(.A(G64gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(G57gat), .ZN(new_n478_));
  INV_X1    g277(.A(G57gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(G64gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n480_), .A3(KEYINPUT11), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n473_), .A2(KEYINPUT11), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n475_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT68), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n478_), .A2(new_n480_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT11), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n481_), .A3(new_n476_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n475_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n430_), .B1(new_n472_), .B2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n485_), .A2(new_n491_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n465_), .A2(new_n467_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT8), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n462_), .A2(new_n464_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n456_), .B(new_n467_), .C1(new_n497_), .C2(new_n444_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n439_), .A2(new_n448_), .A3(new_n431_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT65), .B1(new_n450_), .B2(new_n454_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n494_), .A2(new_n499_), .A3(KEYINPUT69), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n472_), .A2(new_n492_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n493_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(G230gat), .A2(G233gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT12), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n496_), .A2(new_n498_), .B1(new_n501_), .B2(new_n500_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n508_), .B1(new_n509_), .B2(new_n494_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n506_), .B1(new_n509_), .B2(new_n494_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n489_), .A2(KEYINPUT12), .A3(new_n475_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n472_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G120gat), .B(G148gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT5), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G176gat), .B(G204gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n507_), .A2(new_n515_), .A3(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(KEYINPUT70), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT13), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n507_), .A2(new_n515_), .A3(new_n519_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT13), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n504_), .A2(new_n508_), .B1(new_n472_), .B2(new_n513_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n506_), .A2(new_n505_), .B1(new_n526_), .B2(new_n511_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n524_), .B(new_n525_), .C1(new_n527_), .C2(new_n521_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT79), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G29gat), .B(G36gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G43gat), .B(G50gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G29gat), .B(G36gat), .Z(new_n535_));
  XOR2_X1   g334(.A(G43gat), .B(G50gat), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G1gat), .A2(G8gat), .ZN(new_n539_));
  INV_X1    g338(.A(G1gat), .ZN(new_n540_));
  INV_X1    g339(.A(G8gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(KEYINPUT14), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n538_), .A2(new_n539_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n538_), .A2(new_n543_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n534_), .B(new_n537_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n537_), .A2(new_n534_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n538_), .A2(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n542_), .A2(new_n539_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(new_n551_), .A3(new_n544_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT15), .ZN(new_n557_));
  INV_X1    g356(.A(new_n534_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n532_), .A2(new_n533_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n551_), .A2(new_n544_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n537_), .A2(KEYINPUT15), .A3(new_n534_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G113gat), .B(G141gat), .Z(new_n565_));
  XOR2_X1   g364(.A(G169gat), .B(G197gat), .Z(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  NAND3_X1  g366(.A1(new_n556_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n567_), .B1(new_n556_), .B2(new_n564_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI211_X1 g371(.A(new_n569_), .B(new_n567_), .C1(new_n556_), .C2(new_n564_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n531_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n556_), .A2(new_n564_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n567_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(new_n569_), .A3(new_n568_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n573_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(KEYINPUT79), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n530_), .A2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n429_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G134gat), .B(G162gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n587_), .A2(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n560_), .A2(new_n562_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT72), .B1(new_n509_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT72), .ZN(new_n594_));
  INV_X1    g393(.A(new_n592_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n472_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n593_), .A2(new_n596_), .B1(new_n548_), .B2(new_n509_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT34), .Z(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT73), .B1(new_n597_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n509_), .A2(new_n548_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n472_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n594_), .B1(new_n472_), .B2(new_n595_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n603_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT73), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n599_), .A2(new_n600_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n602_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT75), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n599_), .A2(new_n600_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n608_), .B2(KEYINPUT74), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(KEYINPUT74), .B2(new_n608_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n597_), .A2(new_n611_), .A3(new_n614_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n603_), .B(new_n614_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT75), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  AOI211_X1 g417(.A(new_n590_), .B(new_n591_), .C1(new_n610_), .C2(new_n618_), .ZN(new_n619_));
  AND4_X1   g418(.A1(new_n588_), .A2(new_n610_), .A3(new_n618_), .A4(new_n587_), .ZN(new_n620_));
  OAI22_X1  g419(.A1(new_n619_), .A2(new_n620_), .B1(KEYINPUT76), .B2(KEYINPUT37), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n610_), .A2(new_n618_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n591_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n589_), .A3(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n610_), .A2(new_n618_), .A3(new_n588_), .A4(new_n587_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n621_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n561_), .A2(new_n630_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n551_), .A2(G231gat), .A3(G233gat), .A4(new_n544_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n492_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n561_), .A2(new_n630_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n485_), .A2(new_n635_), .A3(new_n632_), .A4(new_n491_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G183gat), .B(G211gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(G127gat), .A2(G155gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(G127gat), .A2(G155gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(KEYINPUT16), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT16), .B1(new_n639_), .B2(new_n640_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n638_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n643_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n641_), .A3(new_n637_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT17), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n644_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n634_), .A2(new_n636_), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n484_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n635_), .A2(new_n632_), .A3(new_n475_), .A4(new_n489_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(new_n649_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n651_), .A2(KEYINPUT77), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT77), .B1(new_n651_), .B2(new_n654_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n629_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n584_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n540_), .A3(new_n339_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT38), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n371_), .A2(new_n396_), .A3(new_n402_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n341_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n424_), .A2(new_n371_), .A3(new_n402_), .ZN(new_n667_));
  AOI22_X1  g466(.A1(new_n411_), .A2(new_n416_), .B1(new_n339_), .B2(new_n421_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n619_), .A2(new_n620_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n572_), .A2(new_n573_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n529_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT100), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(new_n657_), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT101), .ZN(new_n677_));
  OAI21_X1  g476(.A(G1gat), .B1(new_n677_), .B2(new_n340_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n663_), .A2(new_n678_), .ZN(G1324gat));
  NAND2_X1  g478(.A1(new_n278_), .A2(new_n286_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G8gat), .B1(new_n676_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT39), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n661_), .A2(new_n541_), .A3(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT40), .Z(G1325gat));
  NOR2_X1   g485(.A1(new_n677_), .A2(new_n424_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT102), .B1(new_n687_), .B2(new_n375_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n689_), .B(G15gat), .C1(new_n677_), .C2(new_n424_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n661_), .A2(new_n375_), .A3(new_n396_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n688_), .A2(KEYINPUT41), .A3(new_n690_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n693_), .A2(new_n694_), .A3(new_n695_), .ZN(G1326gat));
  OAI21_X1  g495(.A(G22gat), .B1(new_n677_), .B2(new_n427_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT42), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n427_), .A2(G22gat), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT103), .Z(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n660_), .B2(new_n700_), .ZN(G1327gat));
  NAND2_X1  g500(.A1(new_n624_), .A2(new_n625_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n657_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n583_), .B(new_n703_), .C1(new_n666_), .C2(new_n669_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n429_), .A2(KEYINPUT105), .A3(new_n583_), .A4(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G29gat), .B1(new_n709_), .B2(new_n339_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n670_), .B2(new_n628_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n429_), .A2(new_n629_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n675_), .A2(new_n658_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n712_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n711_), .B(new_n717_), .C1(new_n713_), .C2(new_n715_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n339_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n710_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n681_), .A2(G36gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n706_), .A2(new_n707_), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n670_), .A2(KEYINPUT43), .A3(new_n628_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n714_), .B1(new_n429_), .B2(new_n629_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n711_), .B1(new_n732_), .B2(new_n717_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n716_), .A2(new_n718_), .A3(new_n712_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n680_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n729_), .B1(new_n735_), .B2(G36gat), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n724_), .B(new_n725_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n727_), .B(KEYINPUT45), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n719_), .A2(new_n720_), .A3(new_n681_), .ZN(new_n740_));
  INV_X1    g539(.A(G36gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT107), .B1(new_n742_), .B2(KEYINPUT106), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT46), .B1(new_n736_), .B2(new_n724_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n738_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(G1329gat));
  NAND3_X1  g545(.A1(new_n721_), .A2(G43gat), .A3(new_n396_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n708_), .A2(new_n424_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(G43gat), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g549(.A(new_n427_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G50gat), .B1(new_n709_), .B2(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n751_), .A2(G50gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n721_), .B2(new_n753_), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n529_), .A2(new_n673_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n429_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n659_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(KEYINPUT108), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n339_), .B1(new_n757_), .B2(KEYINPUT108), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n479_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n574_), .A2(new_n657_), .A3(new_n580_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n672_), .A2(new_n530_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n339_), .A2(G57gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT109), .Z(G1332gat));
  OAI21_X1  g565(.A(G64gat), .B1(new_n763_), .B2(new_n681_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n680_), .A2(new_n477_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n757_), .B2(new_n770_), .ZN(G1333gat));
  OAI21_X1  g570(.A(G71gat), .B1(new_n763_), .B2(new_n424_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT49), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n424_), .A2(G71gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n757_), .B2(new_n774_), .ZN(G1334gat));
  OAI21_X1  g574(.A(G78gat), .B1(new_n763_), .B2(new_n427_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT50), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n427_), .A2(G78gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n757_), .B2(new_n778_), .ZN(G1335gat));
  NAND2_X1  g578(.A1(new_n756_), .A2(new_n703_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(G85gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n339_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n716_), .A2(new_n658_), .A3(new_n755_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(new_n339_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n785_), .B2(new_n782_), .ZN(G1336gat));
  AOI21_X1  g585(.A(G92gat), .B1(new_n781_), .B2(new_n680_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n432_), .A2(new_n433_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n681_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n784_), .B2(new_n789_), .ZN(G1337gat));
  NAND2_X1  g589(.A1(new_n396_), .A2(new_n446_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792_));
  OAI22_X1  g591(.A1(new_n780_), .A2(new_n791_), .B1(KEYINPUT111), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n784_), .A2(new_n396_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(G99gat), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(KEYINPUT111), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n795_), .B(new_n796_), .Z(G1338gat));
  NAND3_X1  g596(.A1(new_n781_), .A2(new_n447_), .A3(new_n751_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n447_), .B1(new_n784_), .B2(new_n751_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n799_), .A2(new_n800_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT53), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n798_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1339gat));
  NOR2_X1   g606(.A1(new_n680_), .A2(new_n340_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n665_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(KEYINPUT59), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n515_), .A2(KEYINPUT55), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n526_), .A2(new_n816_), .A3(new_n511_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n510_), .B(new_n514_), .C1(new_n472_), .C2(new_n492_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n815_), .A2(new_n817_), .B1(new_n506_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n814_), .B1(new_n819_), .B2(new_n521_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n521_), .A2(new_n814_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT114), .B1(new_n819_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n818_), .A2(new_n506_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n816_), .B1(new_n526_), .B2(new_n511_), .ZN(new_n825_));
  AND4_X1   g624(.A1(new_n816_), .A2(new_n510_), .A3(new_n511_), .A4(new_n514_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n821_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n820_), .A2(new_n823_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n673_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n520_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n553_), .A2(new_n554_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n563_), .A2(new_n552_), .A3(new_n555_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n576_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n836_), .A2(new_n568_), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT115), .B(new_n837_), .C1(new_n520_), .C2(new_n522_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n524_), .B1(new_n527_), .B2(new_n521_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT115), .B1(new_n840_), .B2(new_n837_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n833_), .A2(new_n842_), .ZN(new_n843_));
  AND4_X1   g642(.A1(new_n813_), .A2(new_n843_), .A3(KEYINPUT57), .A4(new_n702_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n671_), .B1(new_n833_), .B2(new_n842_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n813_), .B1(new_n845_), .B2(KEYINPUT57), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n827_), .A2(new_n821_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n820_), .A2(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n524_), .A2(new_n837_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n851_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n524_), .A2(new_n837_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n855_), .B1(new_n820_), .B2(new_n848_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT58), .B1(new_n856_), .B2(KEYINPUT117), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n629_), .A2(new_n854_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n845_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n837_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n838_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n866_), .A2(KEYINPUT116), .A3(new_n671_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n858_), .B1(new_n861_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n847_), .B1(KEYINPUT119), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT116), .B1(new_n866_), .B2(new_n671_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n843_), .A2(new_n860_), .A3(new_n702_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n859_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n858_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n657_), .B1(new_n869_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n627_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n529_), .B2(new_n762_), .ZN(new_n880_));
  AOI211_X1 g679(.A(KEYINPUT112), .B(new_n761_), .C1(new_n523_), .C2(new_n528_), .ZN(new_n881_));
  OAI22_X1  g680(.A1(new_n876_), .A2(new_n878_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT113), .B1(new_n882_), .B2(KEYINPUT54), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n880_), .A2(new_n881_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT113), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .A4(new_n628_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n882_), .A2(KEYINPUT54), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n883_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n812_), .B1(new_n875_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n658_), .B1(new_n868_), .B2(new_n847_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n889_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n811_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n890_), .B1(new_n891_), .B2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G113gat), .B1(new_n895_), .B2(new_n582_), .ZN(new_n896_));
  AND4_X1   g695(.A1(new_n627_), .A2(new_n854_), .A3(new_n857_), .A4(new_n621_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n843_), .A2(new_n702_), .ZN(new_n898_));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n898_), .B2(KEYINPUT116), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n899_), .B2(new_n871_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT118), .B1(new_n898_), .B2(new_n859_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n845_), .A2(new_n813_), .A3(KEYINPUT57), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n657_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n810_), .B1(new_n904_), .B2(new_n889_), .ZN(new_n905_));
  OR3_X1    g704(.A1(new_n905_), .A2(G113gat), .A3(new_n831_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n896_), .A2(new_n906_), .ZN(G1340gat));
  INV_X1    g706(.A(G120gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n529_), .B1(new_n905_), .B2(KEYINPUT59), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n890_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n908_), .A2(KEYINPUT60), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n529_), .A2(KEYINPUT60), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n908_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n911_), .B1(new_n894_), .B2(new_n914_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n872_), .B(new_n858_), .C1(new_n846_), .C2(new_n844_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n889_), .B1(new_n916_), .B2(new_n658_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n914_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n917_), .A2(KEYINPUT120), .A3(new_n811_), .A4(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n915_), .A2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT121), .B1(new_n910_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n812_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n868_), .A2(KEYINPUT119), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(new_n903_), .A3(new_n874_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n658_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n922_), .B1(new_n925_), .B2(new_n893_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n530_), .B1(new_n894_), .B2(new_n891_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G120gat), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT120), .B1(new_n905_), .B2(new_n918_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n894_), .A2(new_n911_), .A3(new_n914_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n928_), .A2(new_n929_), .A3(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n921_), .A2(new_n933_), .ZN(G1341gat));
  OAI21_X1  g733(.A(G127gat), .B1(new_n895_), .B2(new_n658_), .ZN(new_n935_));
  OR3_X1    g734(.A1(new_n905_), .A2(G127gat), .A3(new_n658_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1342gat));
  OAI21_X1  g736(.A(G134gat), .B1(new_n895_), .B2(new_n628_), .ZN(new_n938_));
  OR3_X1    g737(.A1(new_n905_), .A2(G134gat), .A3(new_n702_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1343gat));
  NOR3_X1   g739(.A1(new_n917_), .A2(new_n664_), .A3(new_n809_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n673_), .ZN(new_n942_));
  XOR2_X1   g741(.A(KEYINPUT122), .B(G141gat), .Z(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1344gat));
  NAND2_X1  g743(.A1(new_n941_), .A2(new_n530_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n947_), .B1(new_n941_), .B2(new_n657_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n941_), .A2(new_n947_), .A3(new_n657_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(KEYINPUT61), .B(G155gat), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n949_), .A2(new_n950_), .A3(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n951_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n892_), .A2(new_n893_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n404_), .ZN(new_n955_));
  NOR4_X1   g754(.A1(new_n955_), .A2(KEYINPUT123), .A3(new_n658_), .A4(new_n809_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n953_), .B1(new_n956_), .B2(new_n948_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n952_), .A2(new_n957_), .ZN(G1346gat));
  INV_X1    g757(.A(new_n941_), .ZN(new_n959_));
  OR3_X1    g758(.A1(new_n959_), .A2(G162gat), .A3(new_n702_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G162gat), .B1(new_n959_), .B2(new_n628_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1347gat));
  NOR2_X1   g761(.A1(new_n681_), .A2(new_n339_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n963_), .A2(new_n396_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(new_n751_), .ZN(new_n965_));
  OAI211_X1 g764(.A(new_n673_), .B(new_n965_), .C1(new_n875_), .C2(new_n889_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(G169gat), .ZN(new_n967_));
  XNOR2_X1  g766(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  AOI211_X1 g768(.A(new_n751_), .B(new_n964_), .C1(new_n925_), .C2(new_n893_), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n970_), .A2(new_n224_), .A3(new_n673_), .ZN(new_n971_));
  INV_X1    g770(.A(new_n968_), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n966_), .A2(G169gat), .A3(new_n972_), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n969_), .A2(new_n971_), .A3(new_n973_), .ZN(G1348gat));
  NAND2_X1  g773(.A1(new_n970_), .A2(new_n530_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n917_), .A2(new_n751_), .ZN(new_n976_));
  INV_X1    g775(.A(G176gat), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n964_), .A2(new_n977_), .A3(new_n529_), .ZN(new_n978_));
  AOI22_X1  g777(.A1(new_n975_), .A2(new_n223_), .B1(new_n976_), .B2(new_n978_), .ZN(G1349gat));
  NOR2_X1   g778(.A1(new_n658_), .A2(new_n232_), .ZN(new_n980_));
  NAND4_X1  g779(.A1(new_n976_), .A2(new_n396_), .A3(new_n657_), .A4(new_n963_), .ZN(new_n981_));
  AOI22_X1  g780(.A1(new_n970_), .A2(new_n980_), .B1(new_n981_), .B2(new_n248_), .ZN(G1350gat));
  NAND3_X1  g781(.A1(new_n970_), .A2(new_n233_), .A3(new_n671_), .ZN(new_n983_));
  OAI211_X1 g782(.A(new_n629_), .B(new_n965_), .C1(new_n875_), .C2(new_n889_), .ZN(new_n984_));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n985_));
  AND3_X1   g784(.A1(new_n984_), .A2(new_n985_), .A3(G190gat), .ZN(new_n986_));
  AOI21_X1  g785(.A(new_n985_), .B1(new_n984_), .B2(G190gat), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n983_), .B1(new_n986_), .B2(new_n987_), .ZN(G1351gat));
  NOR4_X1   g787(.A1(new_n917_), .A2(new_n339_), .A3(new_n664_), .A4(new_n681_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n989_), .A2(new_n673_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(new_n990_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g790(.A1(new_n989_), .A2(new_n530_), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n992_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g792(.A1(new_n954_), .A2(new_n404_), .A3(new_n657_), .A4(new_n963_), .ZN(new_n994_));
  XNOR2_X1  g793(.A(KEYINPUT63), .B(G211gat), .ZN(new_n995_));
  NOR2_X1   g794(.A1(new_n994_), .A2(new_n995_), .ZN(new_n996_));
  INV_X1    g795(.A(KEYINPUT63), .ZN(new_n997_));
  INV_X1    g796(.A(G211gat), .ZN(new_n998_));
  NAND3_X1  g797(.A1(new_n994_), .A2(new_n997_), .A3(new_n998_), .ZN(new_n999_));
  OR2_X1    g798(.A1(new_n999_), .A2(KEYINPUT126), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n999_), .A2(KEYINPUT126), .ZN(new_n1001_));
  AOI21_X1  g800(.A(new_n996_), .B1(new_n1000_), .B2(new_n1001_), .ZN(G1354gat));
  AOI21_X1  g801(.A(G218gat), .B1(new_n989_), .B2(new_n671_), .ZN(new_n1003_));
  NAND2_X1  g802(.A1(new_n629_), .A2(G218gat), .ZN(new_n1004_));
  XNOR2_X1  g803(.A(new_n1004_), .B(KEYINPUT127), .ZN(new_n1005_));
  AOI21_X1  g804(.A(new_n1003_), .B1(new_n989_), .B2(new_n1005_), .ZN(G1355gat));
endmodule


