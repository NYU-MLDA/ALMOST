//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT25), .B(G183gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n210_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n207_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(KEYINPUT78), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G169gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT22), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT79), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT79), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n225_), .A3(KEYINPUT22), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n211_), .A2(KEYINPUT22), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n224_), .A2(new_n212_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n209_), .B2(new_n208_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n230_), .B1(new_n209_), .B2(new_n208_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n231_), .A2(new_n214_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n218_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G197gat), .B(G204gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT21), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G197gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT21), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT85), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n243_), .B2(new_n235_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT86), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n240_), .A2(G204gat), .ZN(new_n246_));
  INV_X1    g045(.A(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G197gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n248_), .A3(new_n237_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n236_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n244_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G218gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G211gat), .ZN(new_n253_));
  INV_X1    g052(.A(G211gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G218gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n237_), .B2(new_n235_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n246_), .A2(new_n248_), .A3(new_n243_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT21), .A3(new_n241_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT86), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n239_), .B1(new_n251_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT87), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n245_), .B1(new_n244_), .B2(new_n250_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n259_), .A3(KEYINPUT86), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n238_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT87), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n234_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT91), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G226gat), .A2(G233gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT19), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n207_), .A2(new_n217_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n263_), .A2(new_n264_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n266_), .B1(new_n275_), .B2(new_n239_), .ZN(new_n276_));
  AOI211_X1 g075(.A(KEYINPUT87), .B(new_n238_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n274_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT91), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(KEYINPUT20), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n217_), .A2(new_n205_), .ZN(new_n281_));
  XOR2_X1   g080(.A(KEYINPUT22), .B(G169gat), .Z(new_n282_));
  OAI211_X1 g081(.A(new_n231_), .B(new_n214_), .C1(G176gat), .C2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n261_), .A2(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n270_), .A2(new_n273_), .A3(new_n280_), .A4(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n261_), .A2(new_n284_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(new_n269_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n262_), .A2(new_n267_), .A3(new_n234_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n272_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT95), .ZN(new_n293_));
  XOR2_X1   g092(.A(G8gat), .B(G36gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(G64gat), .B(G92gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  NAND3_X1  g097(.A1(new_n292_), .A2(new_n293_), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n270_), .A2(new_n285_), .A3(new_n280_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n272_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n298_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n290_), .A2(new_n272_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n301_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n299_), .A2(KEYINPUT27), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n293_), .B1(new_n292_), .B2(new_n298_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT96), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n303_), .B1(new_n300_), .B2(new_n272_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(new_n302_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT96), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n309_), .A2(new_n312_), .A3(new_n313_), .A4(new_n299_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n311_), .A2(new_n302_), .ZN(new_n316_));
  AOI211_X1 g115(.A(new_n298_), .B(new_n303_), .C1(new_n300_), .C2(new_n272_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n310_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G22gat), .B(G50gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT3), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT2), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n326_), .B1(new_n328_), .B2(KEYINPUT1), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT83), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT83), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n333_), .B(new_n326_), .C1(new_n328_), .C2(KEYINPUT1), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n327_), .A2(new_n335_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n332_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT82), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n321_), .A2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n323_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n330_), .B1(new_n337_), .B2(new_n342_), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n343_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n331_), .A2(KEYINPUT83), .B1(new_n335_), .B2(new_n327_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n342_), .B1(new_n346_), .B2(new_n334_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n329_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n345_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n320_), .B1(new_n344_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT28), .B1(new_n343_), .B2(KEYINPUT29), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n345_), .A3(new_n351_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n319_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n343_), .B2(KEYINPUT29), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n262_), .A2(new_n359_), .A3(new_n267_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n350_), .A2(new_n351_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(new_n361_), .B2(new_n265_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT88), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n360_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n357_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT89), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n357_), .B(new_n370_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT90), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n353_), .A2(new_n356_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n360_), .A2(new_n362_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(new_n363_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n372_), .A2(new_n373_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n373_), .B1(new_n372_), .B2(new_n379_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G127gat), .B(G134gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G113gat), .B(G120gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n383_), .A2(new_n384_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n382_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n383_), .A2(new_n384_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(KEYINPUT81), .A3(new_n385_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT31), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G71gat), .B(G99gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(G15gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT30), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n234_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT80), .B(G43gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n274_), .B(new_n398_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n400_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n394_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n404_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n393_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n392_), .B(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G85gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n390_), .B(new_n388_), .C1(new_n347_), .C2(new_n349_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n389_), .A2(new_n385_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n330_), .B(new_n419_), .C1(new_n337_), .C2(new_n342_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n417_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT4), .B1(new_n391_), .B2(new_n343_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n416_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n388_), .A2(new_n390_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n350_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n386_), .A2(new_n387_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n347_), .A2(new_n430_), .A3(new_n349_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT4), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n418_), .A2(new_n417_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n425_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n426_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n415_), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n427_), .A2(new_n436_), .A3(KEYINPUT93), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT93), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n434_), .A2(new_n438_), .A3(new_n415_), .A4(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n411_), .A2(new_n440_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n380_), .A2(new_n381_), .A3(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n315_), .A2(new_n318_), .A3(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n437_), .A2(new_n439_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n302_), .A2(KEYINPUT32), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n301_), .A2(new_n304_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n445_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n292_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT94), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n311_), .A2(new_n302_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n415_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT33), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n429_), .A2(new_n431_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n416_), .B1(new_n455_), .B2(new_n425_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n423_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n454_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n453_), .B1(new_n452_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n451_), .A2(new_n305_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT94), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .A4(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n450_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n380_), .A2(new_n381_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n308_), .A2(new_n314_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n318_), .B(new_n440_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n443_), .B1(new_n469_), .B2(new_n410_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G232gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT6), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G85gat), .B(G92gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n483_));
  NAND2_X1  g282(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n480_), .A2(new_n482_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT66), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n476_), .B1(new_n486_), .B2(new_n479_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n479_), .A2(new_n486_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n481_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT67), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT8), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n489_), .A2(KEYINPUT67), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n485_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n482_), .A2(KEYINPUT9), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT10), .B(G99gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT64), .B(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G85gat), .ZN(new_n498_));
  INV_X1    g297(.A(G92gat), .ZN(new_n499_));
  OR3_X1    g298(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT9), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n494_), .A2(new_n497_), .A3(new_n479_), .A4(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n493_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G29gat), .B(G36gat), .Z(new_n503_));
  XOR2_X1   g302(.A(G43gat), .B(G50gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT15), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n505_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n502_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n473_), .B1(new_n511_), .B2(KEYINPUT70), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n510_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n517_), .A2(KEYINPUT70), .A3(new_n507_), .A4(new_n473_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n513_), .A2(new_n514_), .A3(new_n516_), .A4(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G190gat), .B(G218gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G134gat), .B(G162gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT36), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT71), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n518_), .A2(new_n516_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT72), .B1(new_n512_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n519_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n512_), .A2(new_n525_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n522_), .A2(KEYINPUT36), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n470_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G230gat), .A2(G233gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G57gat), .B(G64gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G71gat), .B(G78gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n536_), .A2(new_n538_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n493_), .A2(new_n543_), .A3(new_n501_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n493_), .B2(new_n501_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n534_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G120gat), .B(G148gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT5), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G176gat), .B(G204gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI211_X1 g350(.A(KEYINPUT12), .B(new_n543_), .C1(new_n493_), .C2(new_n501_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n544_), .A2(new_n545_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(new_n553_), .B2(KEYINPUT12), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n546_), .B(new_n551_), .C1(new_n554_), .C2(new_n534_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n543_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n502_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n493_), .A2(new_n543_), .A3(new_n501_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(KEYINPUT12), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n552_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n534_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n546_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n550_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n555_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  OAI211_X1 g364(.A(KEYINPUT68), .B(new_n550_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT13), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n568_), .A2(KEYINPUT69), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n568_), .A2(KEYINPUT69), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n567_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G15gat), .B(G22gat), .ZN(new_n574_));
  INV_X1    g373(.A(G8gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G1gat), .B(G8gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n506_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT75), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n509_), .A2(new_n579_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n509_), .B(new_n579_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT74), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n586_), .B2(new_n583_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G113gat), .B(G141gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT76), .ZN(new_n589_));
  XOR2_X1   g388(.A(G169gat), .B(G197gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n587_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n565_), .A2(KEYINPUT69), .A3(new_n568_), .A4(new_n566_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n573_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT97), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n573_), .A2(new_n597_), .A3(new_n593_), .A4(new_n594_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT16), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT73), .B1(new_n602_), .B2(KEYINPUT17), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n579_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(new_n556_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n602_), .A2(KEYINPUT17), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(new_n606_), .B2(new_n556_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n532_), .A2(new_n596_), .A3(new_n598_), .A4(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT98), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n202_), .B1(new_n612_), .B2(new_n444_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n470_), .A2(new_n592_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n513_), .A2(new_n516_), .A3(new_n518_), .A4(new_n524_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n531_), .B2(KEYINPUT37), .ZN(new_n619_));
  INV_X1    g418(.A(new_n610_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n573_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n594_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n614_), .A2(new_n621_), .A3(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n625_), .A2(G1gat), .A3(new_n440_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT38), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n613_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT99), .ZN(G1324gat));
  NAND2_X1  g428(.A1(new_n315_), .A2(new_n318_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G8gat), .B1(new_n611_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT39), .ZN(new_n633_));
  INV_X1    g432(.A(new_n625_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n575_), .A3(new_n630_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g436(.A(new_n396_), .B1(new_n612_), .B2(new_n411_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT41), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(new_n396_), .A3(new_n411_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n465_), .B(KEYINPUT100), .Z(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n612_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT42), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n634_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1327gat));
  NAND2_X1  g447(.A1(new_n527_), .A2(new_n530_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n649_), .A2(new_n615_), .B1(new_n617_), .B2(new_n616_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT43), .B1(new_n470_), .B2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n315_), .A2(new_n318_), .A3(new_n442_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n468_), .ZN(new_n653_));
  AOI22_X1  g452(.A1(new_n653_), .A2(new_n315_), .B1(new_n465_), .B2(new_n464_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n652_), .B1(new_n654_), .B2(new_n411_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n619_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n651_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n596_), .A2(new_n598_), .A3(new_n620_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n658_), .A2(KEYINPUT44), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT101), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n651_), .B2(new_n657_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n664_), .A3(KEYINPUT44), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n470_), .A2(KEYINPUT43), .A3(new_n650_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n656_), .B1(new_n655_), .B2(new_n619_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n660_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n666_), .A2(G29gat), .A3(new_n444_), .A4(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(G29gat), .ZN(new_n673_));
  INV_X1    g472(.A(new_n624_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n649_), .A2(new_n610_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n614_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n673_), .B1(new_n678_), .B2(new_n440_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n672_), .A2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT102), .Z(G1328gat));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(KEYINPUT105), .B2(KEYINPUT46), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n630_), .B1(new_n663_), .B2(KEYINPUT44), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n662_), .B2(new_n665_), .ZN(new_n686_));
  INV_X1    g485(.A(G36gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n631_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n689_));
  AND4_X1   g488(.A1(new_n664_), .A2(new_n658_), .A3(KEYINPUT44), .A4(new_n660_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n664_), .B1(new_n663_), .B2(KEYINPUT44), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n689_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(KEYINPUT103), .A3(G36gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n688_), .A2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n677_), .A2(new_n687_), .A3(new_n630_), .A4(new_n614_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n682_), .A2(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n683_), .B1(new_n694_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n683_), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n702_), .B(new_n699_), .C1(new_n688_), .C2(new_n693_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1329gat));
  AND2_X1   g503(.A1(new_n411_), .A2(G43gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n666_), .A2(new_n671_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n666_), .A2(KEYINPUT107), .A3(new_n671_), .A4(new_n705_), .ZN(new_n709_));
  XOR2_X1   g508(.A(KEYINPUT108), .B(G43gat), .Z(new_n710_));
  OAI21_X1  g509(.A(new_n710_), .B1(new_n678_), .B2(new_n410_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n708_), .A2(new_n709_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT47), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n708_), .A2(new_n709_), .A3(new_n714_), .A4(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1330gat));
  INV_X1    g515(.A(new_n465_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n666_), .A2(G50gat), .A3(new_n717_), .A4(new_n671_), .ZN(new_n718_));
  INV_X1    g517(.A(G50gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n678_), .B2(new_n643_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT109), .Z(G1331gat));
  NOR3_X1   g521(.A1(new_n624_), .A2(new_n593_), .A3(new_n620_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n532_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n440_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n470_), .A2(new_n593_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n674_), .A3(new_n621_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n440_), .A2(G57gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(G1332gat));
  OR3_X1    g528(.A1(new_n727_), .A2(G64gat), .A3(new_n631_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G64gat), .B1(new_n724_), .B2(new_n631_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(KEYINPUT48), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(KEYINPUT48), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n730_), .B1(new_n732_), .B2(new_n733_), .ZN(G1333gat));
  OR3_X1    g533(.A1(new_n727_), .A2(G71gat), .A3(new_n410_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n724_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n411_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT49), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(G71gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G71gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n739_), .B2(new_n740_), .ZN(G1334gat));
  OAI21_X1  g540(.A(G78gat), .B1(new_n724_), .B2(new_n643_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(KEYINPUT50), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(KEYINPUT50), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n643_), .A2(G78gat), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT110), .Z(new_n746_));
  OAI22_X1  g545(.A1(new_n743_), .A2(new_n744_), .B1(new_n727_), .B2(new_n746_), .ZN(G1335gat));
  NAND3_X1  g546(.A1(new_n726_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT111), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(KEYINPUT111), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n498_), .A3(new_n444_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n593_), .A2(new_n610_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n674_), .A2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n667_), .A2(new_n668_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n757_), .A2(KEYINPUT112), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(KEYINPUT112), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n756_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(new_n444_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n754_), .B1(new_n761_), .B2(new_n498_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT113), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n754_), .C1(new_n761_), .C2(new_n498_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1336gat));
  NAND3_X1  g565(.A1(new_n753_), .A2(new_n499_), .A3(new_n630_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n760_), .A2(new_n630_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n499_), .ZN(G1337gat));
  NAND3_X1  g568(.A1(new_n753_), .A2(new_n495_), .A3(new_n411_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n760_), .A2(new_n411_), .ZN(new_n771_));
  INV_X1    g570(.A(G99gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT51), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n770_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n753_), .A2(new_n496_), .A3(new_n717_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n658_), .A2(new_n674_), .A3(new_n717_), .A4(new_n755_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781_));
  OAI21_X1  g580(.A(G106gat), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n781_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n779_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n784_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n786_), .A2(new_n782_), .A3(KEYINPUT52), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n778_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n790_), .B(new_n778_), .C1(new_n785_), .C2(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1339gat));
  NOR2_X1   g591(.A1(new_n593_), .A2(new_n620_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n573_), .A2(new_n793_), .A3(new_n594_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT115), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n650_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT54), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n554_), .A2(new_n534_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  OR3_X1    g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n561_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n551_), .B1(new_n561_), .B2(new_n799_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n593_), .A2(KEYINPUT116), .A3(new_n555_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT116), .B1(new_n593_), .B2(new_n555_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n806_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n583_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n581_), .A2(new_n582_), .A3(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n812_), .B(new_n591_), .C1(new_n586_), .C2(new_n811_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n587_), .B2(new_n591_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n567_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n649_), .C1(new_n810_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n806_), .B2(new_n809_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n531_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n555_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n820_), .A2(new_n814_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT58), .B1(new_n822_), .B2(KEYINPUT117), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n619_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n822_), .A2(KEYINPUT117), .A3(KEYINPUT58), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n816_), .B(new_n819_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n620_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n797_), .A2(new_n827_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n630_), .A2(new_n440_), .A3(new_n410_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n465_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n593_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n717_), .B1(new_n797_), .B2(new_n827_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(KEYINPUT59), .A3(new_n829_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(G113gat), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n592_), .A2(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT118), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n832_), .B1(new_n837_), .B2(new_n840_), .ZN(G1340gat));
  INV_X1    g640(.A(G120gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n624_), .B2(KEYINPUT60), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n831_), .B(new_n843_), .C1(KEYINPUT60), .C2(new_n842_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n624_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n842_), .ZN(G1341gat));
  AOI21_X1  g645(.A(G127gat), .B1(new_n831_), .B2(new_n610_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT119), .B(G127gat), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n610_), .A2(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT120), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n847_), .B1(new_n837_), .B2(new_n850_), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n831_), .A2(new_n852_), .A3(new_n531_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n650_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n852_), .ZN(G1343gat));
  NOR4_X1   g654(.A1(new_n630_), .A2(new_n440_), .A3(new_n465_), .A4(new_n411_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT121), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n828_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n593_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n674_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g662(.A1(new_n858_), .A2(new_n620_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT61), .B(G155gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  OR3_X1    g665(.A1(new_n858_), .A2(G162gat), .A3(new_n649_), .ZN(new_n867_));
  OAI21_X1  g666(.A(G162gat), .B1(new_n858_), .B2(new_n650_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1347gat));
  AOI21_X1  g668(.A(new_n211_), .B1(KEYINPUT122), .B2(KEYINPUT62), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n631_), .A2(new_n441_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n871_), .A2(new_n643_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n828_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n870_), .B1(new_n873_), .B2(new_n592_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI221_X1 g675(.A(new_n870_), .B1(KEYINPUT122), .B2(KEYINPUT62), .C1(new_n873_), .C2(new_n592_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n873_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n593_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n876_), .B(new_n877_), .C1(new_n282_), .C2(new_n879_), .ZN(G1348gat));
  AOI21_X1  g679(.A(G176gat), .B1(new_n878_), .B2(new_n674_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n835_), .A2(new_n871_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n624_), .A2(new_n212_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(G1349gat));
  AOI21_X1  g683(.A(G183gat), .B1(new_n882_), .B2(new_n610_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n873_), .A2(new_n620_), .A3(new_n203_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n873_), .B2(new_n650_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n531_), .A2(new_n204_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n873_), .B2(new_n889_), .ZN(G1351gat));
  NOR4_X1   g689(.A1(new_n631_), .A2(new_n444_), .A3(new_n465_), .A4(new_n411_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n828_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n240_), .A2(KEYINPUT123), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(new_n593_), .A3(new_n894_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT123), .B(G197gat), .Z(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n892_), .B2(new_n592_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1352gat));
  NOR2_X1   g697(.A1(new_n892_), .A2(new_n624_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n247_), .ZN(G1353gat));
  AOI21_X1  g699(.A(new_n620_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT124), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT125), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n893_), .A2(new_n902_), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n893_), .A2(new_n902_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n903_), .B(KEYINPUT125), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(G1354gat));
  NAND3_X1  g707(.A1(new_n828_), .A2(new_n619_), .A3(new_n891_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n909_), .A2(G218gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n531_), .A2(new_n252_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n892_), .A2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT126), .B1(new_n910_), .B2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n909_), .A2(G218gat), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n914_), .B(new_n915_), .C1(new_n892_), .C2(new_n911_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n916_), .ZN(G1355gat));
endmodule


