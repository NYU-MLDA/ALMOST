//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n842_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_;
  NOR2_X1   g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n202_), .B1(new_n205_), .B2(KEYINPUT9), .ZN(new_n206_));
  INV_X1    g005(.A(new_n205_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT9), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n207_), .A2(KEYINPUT66), .A3(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT66), .B1(new_n207_), .B2(new_n208_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT10), .B(G99gat), .Z(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n211_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT7), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n221_), .B(new_n222_), .C1(G99gat), .C2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n224_), .B(new_n218_), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n226_), .A2(new_n216_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n205_), .A2(new_n202_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT8), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT68), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(KEYINPUT68), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n226_), .A2(KEYINPUT70), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n213_), .A2(new_n215_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n216_), .A2(KEYINPUT69), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n223_), .A2(new_n225_), .A3(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n235_), .A2(new_n237_), .A3(new_n238_), .A4(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n229_), .B1(new_n241_), .B2(new_n228_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n234_), .B1(new_n242_), .B2(KEYINPUT71), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n244_));
  AOI211_X1 g043(.A(new_n244_), .B(new_n229_), .C1(new_n241_), .C2(new_n228_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n220_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT72), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(KEYINPUT72), .B(new_n220_), .C1(new_n243_), .C2(new_n245_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G64gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n251_));
  XOR2_X1   g050(.A(G71gat), .B(G78gat), .Z(new_n252_));
  AND2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(KEYINPUT11), .B2(new_n250_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n251_), .A2(new_n252_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT12), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n248_), .A2(new_n249_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n246_), .A2(new_n257_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n256_), .B(new_n220_), .C1(new_n243_), .C2(new_n245_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G230gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(KEYINPUT73), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT73), .B1(new_n264_), .B2(new_n267_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n260_), .B(new_n263_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n261_), .A2(new_n264_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n267_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G120gat), .B(G148gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT5), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G176gat), .B(G204gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  OR2_X1    g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n279_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT13), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(KEYINPUT13), .A3(new_n281_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n286_), .A2(KEYINPUT74), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(KEYINPUT74), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G29gat), .B(G36gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G43gat), .B(G50gat), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n291_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT15), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296_));
  INV_X1    g095(.A(G1gat), .ZN(new_n297_));
  INV_X1    g096(.A(G8gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT14), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G1gat), .B(G8gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n294_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(new_n302_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G229gat), .A2(G233gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n304_), .B(new_n302_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n306_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G113gat), .B(G141gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G169gat), .B(G197gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  NAND3_X1  g112(.A1(new_n307_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT79), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n307_), .A2(new_n310_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT80), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT80), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n315_), .A2(new_n320_), .A3(new_n317_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n289_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  OR3_X1    g123(.A1(new_n324_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT84), .B1(new_n324_), .B2(KEYINPUT23), .ZN(new_n326_));
  INV_X1    g125(.A(new_n324_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n325_), .B(new_n326_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT82), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  OR3_X1    g133(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT25), .B(G183gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT81), .B1(new_n337_), .B2(G190gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(G190gat), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n336_), .B(new_n338_), .C1(new_n339_), .C2(KEYINPUT81), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n329_), .A2(new_n334_), .A3(new_n335_), .A4(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT86), .B(G176gat), .ZN(new_n342_));
  INV_X1    g141(.A(G169gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT85), .B1(new_n343_), .B2(KEYINPUT22), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT22), .B(G169gat), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n342_), .B(new_n344_), .C1(new_n345_), .C2(KEYINPUT85), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n324_), .A2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n328_), .B2(new_n324_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n346_), .B(new_n331_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n341_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT88), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n352_), .B(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G71gat), .B(G99gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(G15gat), .B(G43gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(KEYINPUT87), .B(KEYINPUT30), .Z(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n355_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT89), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G127gat), .B(G134gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(G113gat), .B(G120gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT31), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n361_), .A2(new_n362_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n363_), .A2(new_n369_), .A3(new_n367_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G22gat), .B(G50gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G197gat), .B(G204gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT21), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n376_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G211gat), .B(G218gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  OR3_X1    g179(.A1(new_n375_), .A2(new_n379_), .A3(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT3), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G141gat), .A2(G148gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT2), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(KEYINPUT1), .B2(new_n388_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(KEYINPUT1), .B2(new_n388_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n383_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(new_n385_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n382_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(G228gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(G228gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n399_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n398_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n404_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n382_), .B(new_n407_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT90), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n406_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT92), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n396_), .A2(new_n397_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT28), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n405_), .A2(new_n408_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n406_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT92), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n417_), .A2(KEYINPUT90), .A3(new_n418_), .A4(new_n409_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n412_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n414_), .B1(new_n412_), .B2(new_n419_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n374_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n422_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n373_), .A3(new_n420_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n391_), .A2(new_n395_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(new_n366_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(new_n431_), .A3(new_n366_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n429_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n430_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G1gat), .B(G29gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G57gat), .B(G85gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n440_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n380_), .A2(new_n381_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(new_n351_), .A3(new_n341_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n330_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n335_), .B1(new_n446_), .B2(new_n332_), .ZN(new_n447_));
  AOI211_X1 g246(.A(new_n447_), .B(new_n349_), .C1(new_n336_), .C2(new_n339_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n342_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n345_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n331_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n350_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n329_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n448_), .A2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n445_), .B(KEYINPUT20), .C1(new_n454_), .C2(new_n444_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G226gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT19), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n444_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n457_), .B1(new_n352_), .B2(new_n382_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT20), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G8gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT18), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G64gat), .B(G92gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT32), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT96), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n443_), .B1(new_n462_), .B2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n455_), .A2(new_n457_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n459_), .A2(KEYINPUT20), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n471_), .A2(KEYINPUT97), .B1(new_n382_), .B2(new_n352_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(KEYINPUT97), .B2(new_n471_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n470_), .B1(new_n473_), .B2(new_n457_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT98), .B1(new_n474_), .B2(new_n467_), .ZN(new_n475_));
  OR3_X1    g274(.A1(new_n474_), .A2(KEYINPUT98), .A3(new_n467_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n469_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n441_), .A2(new_n478_), .ZN(new_n479_));
  OR3_X1    g278(.A1(new_n435_), .A2(new_n478_), .A3(new_n440_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n440_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n481_), .A2(KEYINPUT95), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(KEYINPUT95), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n482_), .B(new_n483_), .C1(new_n434_), .C2(new_n433_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n479_), .A2(new_n480_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n466_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n462_), .A2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n487_), .A2(KEYINPUT93), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(KEYINPUT93), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n462_), .A2(new_n486_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n426_), .B1(new_n477_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n423_), .A2(new_n425_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n466_), .B(KEYINPUT99), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n474_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT27), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n487_), .A2(new_n497_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n496_), .A2(new_n498_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n443_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n494_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n372_), .B1(new_n493_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT100), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n426_), .A2(new_n503_), .A3(new_n499_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n496_), .A2(new_n498_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n491_), .A2(new_n497_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT100), .B1(new_n494_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n371_), .A2(new_n443_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n502_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n323_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n248_), .A2(new_n295_), .A3(new_n249_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G232gat), .A2(G233gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT34), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(KEYINPUT35), .ZN(new_n516_));
  INV_X1    g315(.A(new_n220_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n241_), .A2(new_n228_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT8), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n233_), .B1(new_n519_), .B2(new_n244_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n245_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n517_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n516_), .B1(new_n522_), .B2(new_n294_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n515_), .A2(KEYINPUT35), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n513_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n524_), .B1(new_n513_), .B2(new_n523_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G190gat), .B(G218gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(G134gat), .B(G162gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n531_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT75), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT76), .B1(new_n527_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT76), .ZN(new_n538_));
  NOR4_X1   g337(.A1(new_n525_), .A2(new_n526_), .A3(new_n538_), .A4(new_n535_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n533_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n533_), .B(KEYINPUT37), .C1(new_n537_), .C2(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G127gat), .B(G155gat), .Z(new_n545_));
  XNOR2_X1  g344(.A(G183gat), .B(G211gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT17), .Z(new_n550_));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n302_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(new_n257_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT78), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n549_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(KEYINPUT17), .A3(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(new_n555_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n544_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n512_), .A2(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n563_), .A2(G1gat), .A3(new_n500_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n564_), .A2(KEYINPUT38), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(KEYINPUT38), .ZN(new_n566_));
  INV_X1    g365(.A(new_n540_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n511_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n560_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(new_n323_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n297_), .B1(new_n570_), .B2(new_n443_), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n565_), .A2(new_n566_), .A3(new_n571_), .ZN(G1324gat));
  INV_X1    g371(.A(KEYINPUT39), .ZN(new_n573_));
  OAI21_X1  g372(.A(G8gat), .B1(new_n573_), .B2(KEYINPUT101), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n570_), .B2(new_n507_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n573_), .A2(KEYINPUT101), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n563_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n298_), .A3(new_n507_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT40), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(G1325gat));
  NOR3_X1   g381(.A1(new_n563_), .A2(G15gat), .A3(new_n371_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT102), .ZN(new_n584_));
  INV_X1    g383(.A(G15gat), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n570_), .B2(new_n372_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT41), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n587_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n588_), .A3(new_n589_), .ZN(G1326gat));
  INV_X1    g389(.A(G22gat), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n570_), .B2(new_n494_), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n578_), .A2(new_n591_), .A3(new_n494_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(G1327gat));
  NOR2_X1   g395(.A1(new_n540_), .A2(new_n560_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n512_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n598_), .A2(G29gat), .A3(new_n500_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n323_), .A2(new_n560_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n544_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT43), .B1(new_n511_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n509_), .A2(new_n510_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n493_), .A2(new_n501_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(new_n372_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT43), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n544_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n600_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT44), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n600_), .A2(new_n608_), .A3(KEYINPUT44), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n443_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n599_), .B1(new_n615_), .B2(G29gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT104), .ZN(G1328gat));
  NOR2_X1   g416(.A1(new_n499_), .A2(G36gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT106), .B1(new_n598_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT106), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n512_), .A2(new_n621_), .A3(new_n597_), .A4(new_n618_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n620_), .A2(KEYINPUT45), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT45), .B1(new_n620_), .B2(new_n622_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n611_), .A2(new_n507_), .A3(new_n612_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n626_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT105), .B1(new_n626_), .B2(G36gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT46), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n625_), .B(KEYINPUT46), .C1(new_n627_), .C2(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1329gat));
  NAND2_X1  g432(.A1(new_n372_), .A2(G43gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n598_), .A2(new_n371_), .ZN(new_n635_));
  OAI22_X1  g434(.A1(new_n613_), .A2(new_n634_), .B1(G43gat), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g436(.A(new_n598_), .ZN(new_n638_));
  AOI21_X1  g437(.A(G50gat), .B1(new_n638_), .B2(new_n494_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n494_), .A2(G50gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n614_), .B2(new_n640_), .ZN(G1331gat));
  INV_X1    g440(.A(new_n322_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n605_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT107), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n287_), .A2(new_n288_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n644_), .A2(new_n562_), .A3(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT108), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT108), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n500_), .A2(G57gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(G57gat), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n322_), .A2(new_n561_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n568_), .A2(new_n645_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(new_n653_), .B2(new_n443_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT109), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT109), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n650_), .A2(new_n658_), .A3(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(G1332gat));
  INV_X1    g459(.A(G64gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n653_), .B2(new_n507_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT48), .Z(new_n663_));
  NOR2_X1   g462(.A1(new_n499_), .A2(G64gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT110), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n646_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT111), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1333gat));
  INV_X1    g468(.A(G71gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n653_), .B2(new_n372_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT49), .Z(new_n672_));
  NAND3_X1  g471(.A1(new_n646_), .A2(new_n670_), .A3(new_n372_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1334gat));
  INV_X1    g473(.A(G78gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n653_), .B2(new_n494_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT50), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n494_), .A2(new_n675_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT112), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n646_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT113), .ZN(G1335gat));
  AND2_X1   g481(.A1(new_n645_), .A2(new_n597_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n644_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n203_), .A3(new_n443_), .ZN(new_n685_));
  AND4_X1   g484(.A1(new_n561_), .A2(new_n608_), .A3(new_n642_), .A4(new_n645_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(new_n443_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(new_n687_), .B2(new_n203_), .ZN(G1336gat));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n204_), .A3(new_n507_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n686_), .A2(new_n507_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(new_n204_), .ZN(G1337gat));
  AOI21_X1  g490(.A(new_n224_), .B1(new_n686_), .B2(new_n372_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n372_), .A2(new_n217_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n684_), .B2(new_n693_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g494(.A1(new_n684_), .A2(new_n218_), .A3(new_n494_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n218_), .B1(new_n686_), .B2(new_n494_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT52), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n698_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT53), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT53), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n703_), .B(new_n696_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1339gat));
  INV_X1    g504(.A(KEYINPUT120), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT118), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n371_), .A2(new_n500_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT115), .B1(new_n509_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n509_), .A2(KEYINPUT115), .A3(new_n708_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n322_), .A2(new_n280_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT55), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n271_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n264_), .A2(new_n267_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT73), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n268_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n720_), .A2(KEYINPUT55), .A3(new_n260_), .A4(new_n263_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n260_), .A2(new_n264_), .A3(new_n263_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n260_), .A2(new_n263_), .A3(KEYINPUT114), .A4(new_n264_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n273_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n716_), .B(new_n721_), .C1(new_n724_), .C2(new_n726_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n727_), .A2(KEYINPUT56), .A3(new_n279_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT56), .B1(new_n727_), .B2(new_n279_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n714_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n313_), .B1(new_n308_), .B2(new_n306_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n303_), .A2(new_n305_), .A3(new_n309_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n315_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n282_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n567_), .B1(new_n730_), .B2(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n280_), .A2(new_n734_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT58), .B(new_n737_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n544_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n724_), .A2(new_n726_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n716_), .A2(new_n721_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n279_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT56), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n727_), .A2(KEYINPUT56), .A3(new_n279_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT58), .B1(new_n746_), .B2(new_n737_), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n736_), .A2(KEYINPUT57), .B1(new_n739_), .B2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n713_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n735_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n540_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT57), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n561_), .B1(new_n748_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n284_), .A2(new_n285_), .A3(new_n652_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n601_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n601_), .B2(new_n756_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n712_), .B1(new_n754_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT59), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT116), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n757_), .A2(new_n758_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n751_), .A2(new_n752_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n736_), .A2(KEYINPUT57), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n765_), .B(new_n766_), .C1(new_n747_), .C2(new_n739_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n764_), .B1(new_n767_), .B2(new_n561_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n763_), .B(KEYINPUT59), .C1(new_n768_), .C2(new_n712_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n762_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n711_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT117), .B1(new_n771_), .B2(new_n709_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n710_), .A2(new_n773_), .A3(new_n711_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n774_), .A3(new_n761_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n768_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n707_), .B1(new_n770_), .B2(new_n777_), .ZN(new_n778_));
  AOI211_X1 g577(.A(KEYINPUT118), .B(new_n776_), .C1(new_n762_), .C2(new_n769_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n322_), .A2(G113gat), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT119), .Z(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n778_), .A2(new_n779_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n760_), .A2(new_n322_), .ZN(new_n784_));
  INV_X1    g583(.A(G113gat), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n706_), .B1(new_n783_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n770_), .A2(new_n777_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT118), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n770_), .A2(new_n707_), .A3(new_n777_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n781_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(KEYINPUT120), .A3(new_n786_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(new_n793_), .ZN(G1340gat));
  OAI21_X1  g593(.A(G120gat), .B1(new_n789_), .B2(new_n289_), .ZN(new_n795_));
  INV_X1    g594(.A(G120gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n289_), .B2(KEYINPUT60), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n760_), .B(new_n797_), .C1(KEYINPUT60), .C2(new_n796_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n795_), .A2(new_n798_), .ZN(G1341gat));
  INV_X1    g598(.A(G127gat), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n760_), .A2(new_n800_), .A3(new_n560_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n778_), .A2(new_n779_), .A3(new_n561_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n800_), .ZN(G1342gat));
  INV_X1    g602(.A(G134gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n760_), .A2(new_n804_), .A3(new_n567_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n778_), .A2(new_n779_), .A3(new_n601_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n804_), .ZN(G1343gat));
  NAND2_X1  g606(.A1(new_n754_), .A2(new_n759_), .ZN(new_n808_));
  NOR4_X1   g607(.A1(new_n426_), .A2(new_n507_), .A3(new_n500_), .A4(new_n372_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n322_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n645_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g614(.A1(new_n810_), .A2(new_n561_), .ZN(new_n816_));
  XOR2_X1   g615(.A(KEYINPUT61), .B(G155gat), .Z(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1346gat));
  OAI21_X1  g617(.A(G162gat), .B1(new_n810_), .B2(new_n601_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n540_), .A2(G162gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n810_), .B2(new_n820_), .ZN(G1347gat));
  AND3_X1   g620(.A1(new_n426_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n808_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n322_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G169gat), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n825_), .A2(KEYINPUT121), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT62), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(KEYINPUT121), .B2(new_n825_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n824_), .A2(new_n450_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1348gat));
  AND3_X1   g631(.A1(new_n823_), .A2(G176gat), .A3(new_n645_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n833_), .A2(KEYINPUT123), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(KEYINPUT123), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n449_), .B1(new_n823_), .B2(new_n645_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n836_), .A2(KEYINPUT122), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(KEYINPUT122), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n834_), .A2(new_n835_), .B1(new_n837_), .B2(new_n838_), .ZN(G1349gat));
  NAND2_X1  g638(.A1(new_n823_), .A2(new_n560_), .ZN(new_n840_));
  MUX2_X1   g639(.A(new_n336_), .B(G183gat), .S(new_n840_), .Z(G1350gat));
  INV_X1    g640(.A(new_n823_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G190gat), .B1(new_n842_), .B2(new_n601_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n823_), .A2(new_n567_), .A3(new_n339_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1351gat));
  NAND3_X1  g644(.A1(new_n494_), .A2(new_n500_), .A3(new_n371_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n507_), .B1(new_n846_), .B2(KEYINPUT124), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(KEYINPUT124), .B2(new_n846_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n808_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n322_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n645_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G204gat), .ZN(new_n853_));
  XOR2_X1   g652(.A(new_n853_), .B(KEYINPUT125), .Z(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(G204gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT126), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1353gat));
  NAND2_X1  g656(.A1(new_n849_), .A2(new_n560_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n859_));
  AND2_X1   g658(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n858_), .B2(new_n859_), .ZN(G1354gat));
  INV_X1    g661(.A(G218gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n849_), .A2(new_n863_), .A3(new_n567_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n849_), .A2(new_n544_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n863_), .ZN(G1355gat));
endmodule


