//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT69), .B(G8gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G1gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n204_), .B2(KEYINPUT14), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT70), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT70), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n205_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n207_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G29gat), .B(G36gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n216_), .B(new_n217_), .Z(new_n218_));
  OR3_X1    g017(.A1(new_n213_), .A2(KEYINPUT72), .A3(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT72), .B1(new_n213_), .B2(new_n218_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n216_), .B(new_n217_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT15), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n213_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT73), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n219_), .A2(new_n220_), .B1(new_n218_), .B2(new_n213_), .ZN(new_n228_));
  OAI22_X1  g027(.A1(new_n223_), .A2(new_n227_), .B1(new_n228_), .B2(new_n222_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G113gat), .B(G141gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G169gat), .B(G197gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n230_), .B(new_n231_), .Z(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT74), .ZN(new_n235_));
  OAI221_X1 g034(.A(new_n232_), .B1(new_n228_), .B2(new_n222_), .C1(new_n223_), .C2(new_n227_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n229_), .A2(KEYINPUT74), .A3(new_n233_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240_));
  INV_X1    g039(.A(G183gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT76), .B1(new_n241_), .B2(KEYINPUT25), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(G183gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n241_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(KEYINPUT75), .A2(G183gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(KEYINPUT25), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT77), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT26), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n252_), .B1(new_n253_), .B2(G190gat), .ZN(new_n254_));
  INV_X1    g053(.A(G190gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT77), .A3(KEYINPUT26), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(G190gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n240_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n260_), .A2(KEYINPUT78), .A3(new_n250_), .A4(new_n246_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G183gat), .A2(G190gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT23), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G176gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n264_), .B(new_n265_), .C1(new_n268_), .C2(KEYINPUT24), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT24), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n270_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n268_), .A2(KEYINPUT79), .A3(KEYINPUT24), .A4(new_n271_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n269_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n259_), .A2(new_n261_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT81), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n264_), .A2(new_n265_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n248_), .A2(new_n249_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(G190gat), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT80), .B1(new_n266_), .B2(KEYINPUT22), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n267_), .B(new_n282_), .C1(new_n283_), .C2(KEYINPUT80), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n284_), .A3(new_n271_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n277_), .A2(new_n278_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n278_), .B1(new_n277_), .B2(new_n285_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT82), .B(G15gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G227gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n286_), .A2(new_n287_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n290_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n277_), .A2(new_n285_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT81), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n277_), .A2(new_n278_), .A3(new_n285_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n292_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT83), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G127gat), .B(G134gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G113gat), .B(G120gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n299_), .A2(new_n300_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n298_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G127gat), .B(G134gat), .Z(new_n304_));
  XOR2_X1   g103(.A(G113gat), .B(G120gat), .Z(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT83), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n297_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G71gat), .B(G99gat), .ZN(new_n311_));
  INV_X1    g110(.A(G43gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT30), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT31), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n297_), .A2(new_n308_), .ZN(new_n317_));
  OR3_X1    g116(.A1(new_n310_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n310_), .B2(new_n317_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT18), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G64gat), .B(G92gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  XOR2_X1   g123(.A(new_n324_), .B(KEYINPUT101), .Z(new_n325_));
  INV_X1    g124(.A(G218gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G211gat), .ZN(new_n327_));
  INV_X1    g126(.A(G211gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G218gat), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n327_), .A2(new_n329_), .A3(KEYINPUT91), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT91), .B1(new_n327_), .B2(new_n329_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G197gat), .ZN(new_n333_));
  INV_X1    g132(.A(G204gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT90), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT90), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G204gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G197gat), .A2(G204gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT92), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT92), .ZN(new_n341_));
  INV_X1    g140(.A(new_n339_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT90), .B(G204gat), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n341_), .B(new_n342_), .C1(new_n343_), .C2(new_n333_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n332_), .A2(new_n340_), .A3(KEYINPUT21), .A4(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(G197gat), .B1(new_n335_), .B2(new_n337_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT89), .B1(new_n333_), .B2(G204gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT89), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(new_n334_), .A3(G197gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT21), .B1(new_n346_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n327_), .A2(new_n329_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT91), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n327_), .A2(new_n329_), .A3(KEYINPUT91), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n351_), .A2(new_n353_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n345_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n294_), .A2(new_n295_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT25), .B(G183gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT96), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT26), .B(G190gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n272_), .A2(new_n273_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n269_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n279_), .B1(G183gat), .B2(G190gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n271_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n283_), .B2(new_n267_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n363_), .B1(new_n375_), .B2(new_n360_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT19), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n362_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n360_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n367_), .A2(new_n369_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n363_), .B1(new_n361_), .B2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n379_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT99), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n380_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AOI211_X1 g185(.A(KEYINPUT99), .B(new_n379_), .C1(new_n381_), .C2(new_n383_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n325_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n286_), .A2(new_n287_), .A3(new_n360_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT20), .B1(new_n361_), .B2(new_n382_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n378_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n381_), .A2(new_n379_), .A3(new_n383_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n324_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(KEYINPUT27), .A3(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G1gat), .B(G29gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G85gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT0), .B(G57gat), .ZN(new_n397_));
  XOR2_X1   g196(.A(new_n396_), .B(new_n397_), .Z(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT1), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(G155gat), .A3(G162gat), .ZN(new_n403_));
  OR2_X1    g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n401_), .A2(new_n403_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n402_), .A2(KEYINPUT84), .A3(G155gat), .A4(G162gat), .ZN(new_n407_));
  INV_X1    g206(.A(G141gat), .ZN(new_n408_));
  INV_X1    g207(.A(G148gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G141gat), .A2(G148gat), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n406_), .A2(new_n407_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT2), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .A4(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n404_), .A2(new_n400_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n413_), .A2(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT98), .B(KEYINPUT4), .Z(new_n424_));
  NAND4_X1  g223(.A1(new_n303_), .A2(new_n423_), .A3(new_n307_), .A4(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n299_), .A2(new_n300_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n306_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT97), .B1(new_n431_), .B2(new_n423_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n303_), .A2(new_n423_), .A3(new_n307_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n407_), .A2(new_n411_), .A3(new_n410_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n434_), .A2(new_n406_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT97), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n430_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n432_), .A2(KEYINPUT4), .A3(new_n433_), .A4(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n428_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n437_), .A3(new_n433_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n427_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n399_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n428_), .A2(new_n438_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(new_n398_), .C1(new_n427_), .C2(new_n440_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT95), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G228gat), .A2(G233gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n423_), .A2(KEYINPUT29), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G78gat), .B(G106gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT93), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n360_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n452_), .B1(new_n360_), .B2(new_n449_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n448_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n360_), .A2(new_n449_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n451_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n448_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n360_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G22gat), .B(G50gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n462_), .B(new_n463_), .Z(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT29), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n413_), .A2(new_n422_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n435_), .A2(KEYINPUT85), .A3(new_n466_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n471_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n465_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n469_), .A2(new_n470_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n471_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n472_), .A3(new_n464_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n447_), .B1(new_n461_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n455_), .A2(new_n460_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n475_), .A2(new_n479_), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n482_), .A2(new_n483_), .A3(KEYINPUT95), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n482_), .A2(KEYINPUT94), .A3(new_n483_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT94), .B1(new_n482_), .B2(new_n483_), .ZN(new_n486_));
  OAI22_X1  g285(.A1(new_n481_), .A2(new_n484_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n324_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n381_), .A2(new_n379_), .A3(new_n383_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n379_), .B1(new_n362_), .B2(new_n376_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n393_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT27), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n394_), .A2(new_n446_), .A3(new_n487_), .A4(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n324_), .A2(KEYINPUT32), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n391_), .A2(new_n496_), .A3(new_n392_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n497_), .A2(new_n445_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n496_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n499_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT33), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n444_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n440_), .A2(new_n426_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(new_n398_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n438_), .A2(new_n426_), .A3(new_n425_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n444_), .A2(new_n502_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n503_), .A2(new_n491_), .A3(new_n507_), .A4(new_n393_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n487_), .B1(new_n501_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT100), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n495_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AOI211_X1 g310(.A(KEYINPUT100), .B(new_n487_), .C1(new_n501_), .C2(new_n508_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n320_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT102), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n394_), .A2(new_n494_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(new_n487_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n320_), .A2(new_n445_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n513_), .A2(new_n514_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT102), .B(new_n320_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n239_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G85gat), .B(G92gat), .Z(new_n522_));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n523_), .B(KEYINPUT6), .Z(new_n524_));
  OR3_X1    g323(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n522_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT8), .ZN(new_n529_));
  INV_X1    g328(.A(G106gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT10), .B(G99gat), .Z(new_n531_));
  AOI21_X1  g330(.A(new_n524_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT64), .B(G92gat), .Z(new_n534_));
  INV_X1    g333(.A(G85gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n532_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  XOR2_X1   g340(.A(G71gat), .B(G78gat), .Z(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n541_), .A2(new_n542_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n529_), .A2(new_n539_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n528_), .A2(KEYINPUT8), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n528_), .A2(KEYINPUT8), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n539_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT12), .B1(new_n553_), .B2(new_n547_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G230gat), .A2(G233gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(KEYINPUT65), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT65), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n529_), .A2(new_n558_), .A3(new_n539_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n557_), .A2(new_n559_), .A3(KEYINPUT12), .A4(new_n547_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n555_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n548_), .B1(new_n529_), .B2(new_n539_), .ZN(new_n562_));
  OAI211_X1 g361(.A(G230gat), .B(G233gat), .C1(new_n550_), .C2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G120gat), .B(G148gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n561_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(KEYINPUT13), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT13), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT36), .Z(new_n580_));
  NOR2_X1   g379(.A1(new_n553_), .A2(new_n218_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT68), .Z(new_n582_));
  NAND3_X1  g381(.A1(new_n225_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n582_), .B(new_n583_), .C1(KEYINPUT35), .C2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT35), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n586_), .A2(new_n589_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n580_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n586_), .A2(new_n589_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n579_), .A2(KEYINPUT36), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n586_), .A2(new_n589_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT37), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n592_), .A2(new_n596_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n213_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(new_n547_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n605_), .A2(KEYINPUT17), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(KEYINPUT17), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n605_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n602_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n521_), .A2(new_n576_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(G1gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(new_n445_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT38), .ZN(new_n621_));
  INV_X1    g420(.A(new_n597_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(KEYINPUT103), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(KEYINPUT103), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n239_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n576_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(new_n615_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n445_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n621_), .B1(new_n632_), .B2(new_n619_), .ZN(G1324gat));
  OR3_X1    g432(.A1(new_n617_), .A2(new_n515_), .A3(new_n203_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n516_), .B(new_n629_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n635_), .A2(new_n636_), .A3(G8gat), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n635_), .B2(G8gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g439(.A(G15gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n320_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n630_), .B2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n618_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n644_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(G1326gat));
  NAND2_X1  g447(.A1(new_n630_), .A2(new_n487_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(G22gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n649_), .B2(G22gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n487_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(G22gat), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT105), .Z(new_n655_));
  OAI22_X1  g454(.A1(new_n651_), .A2(new_n652_), .B1(new_n617_), .B2(new_n655_), .ZN(G1327gat));
  NOR2_X1   g455(.A1(new_n628_), .A2(new_n614_), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT43), .B(new_n601_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n513_), .A2(new_n514_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n517_), .A2(new_n518_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n520_), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n660_), .B1(new_n663_), .B2(new_n602_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n657_), .B1(new_n658_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT44), .B(new_n657_), .C1(new_n658_), .C2(new_n664_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n445_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT107), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n667_), .A2(new_n671_), .A3(new_n445_), .A4(new_n668_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n670_), .A2(G29gat), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n576_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n674_), .A2(new_n597_), .A3(new_n614_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n521_), .A2(new_n675_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n676_), .A2(G29gat), .A3(new_n446_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n673_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT108), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n673_), .A2(new_n680_), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1328gat));
  NOR3_X1   g481(.A1(new_n676_), .A2(G36gat), .A3(new_n515_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT45), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n667_), .A2(new_n516_), .A3(new_n668_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT109), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(KEYINPUT46), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT109), .B(new_n689_), .C1(new_n684_), .C2(new_n686_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1329gat));
  AND2_X1   g490(.A1(new_n667_), .A2(new_n668_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(G43gat), .A3(new_n642_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n312_), .B1(new_n676_), .B2(new_n320_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g495(.A(G50gat), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n653_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n521_), .A2(new_n487_), .A3(new_n675_), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n692_), .A2(new_n698_), .B1(new_n697_), .B2(new_n699_), .ZN(G1331gat));
  NOR3_X1   g499(.A1(new_n627_), .A2(new_n615_), .A3(new_n576_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n626_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n446_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n627_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT110), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n674_), .A3(new_n616_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT111), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n446_), .A2(G57gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n703_), .B1(new_n707_), .B2(new_n708_), .ZN(G1332gat));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710_));
  INV_X1    g509(.A(new_n702_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n516_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n710_), .B1(new_n712_), .B2(G64gat), .ZN(new_n713_));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  AOI211_X1 g513(.A(KEYINPUT48), .B(new_n714_), .C1(new_n711_), .C2(new_n516_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n516_), .A2(new_n714_), .ZN(new_n716_));
  OAI22_X1  g515(.A1(new_n713_), .A2(new_n715_), .B1(new_n707_), .B2(new_n716_), .ZN(G1333gat));
  INV_X1    g516(.A(KEYINPUT49), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n711_), .A2(new_n642_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(G71gat), .ZN(new_n720_));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT49), .B(new_n721_), .C1(new_n711_), .C2(new_n642_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n642_), .A2(new_n721_), .ZN(new_n723_));
  OAI22_X1  g522(.A1(new_n720_), .A2(new_n722_), .B1(new_n707_), .B2(new_n723_), .ZN(G1334gat));
  OAI21_X1  g523(.A(G78gat), .B1(new_n702_), .B2(new_n653_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(KEYINPUT50), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(KEYINPUT50), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n653_), .A2(G78gat), .ZN(new_n728_));
  OAI22_X1  g527(.A1(new_n726_), .A2(new_n727_), .B1(new_n707_), .B2(new_n728_), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n597_), .A2(new_n614_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n705_), .A2(new_n674_), .A3(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G85gat), .B1(new_n732_), .B2(new_n445_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n658_), .A2(new_n664_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n627_), .A2(new_n614_), .A3(new_n576_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT112), .Z(new_n737_));
  NOR2_X1   g536(.A1(new_n446_), .A2(new_n535_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n733_), .B1(new_n737_), .B2(new_n738_), .ZN(G1336gat));
  AOI21_X1  g538(.A(G92gat), .B1(new_n732_), .B2(new_n516_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n515_), .A2(new_n534_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n737_), .B2(new_n741_), .ZN(G1337gat));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(KEYINPUT51), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n642_), .A2(new_n531_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n731_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G99gat), .B1(new_n736_), .B2(new_n320_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n744_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n743_), .A2(KEYINPUT51), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT114), .Z(new_n750_));
  XNOR2_X1  g549(.A(new_n748_), .B(new_n750_), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n732_), .A2(new_n530_), .A3(new_n487_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n487_), .B(new_n735_), .C1(new_n658_), .C2(new_n664_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(G106gat), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n753_), .B2(G106gat), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(KEYINPUT52), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n753_), .A2(G106gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT115), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n759_), .B1(new_n761_), .B2(new_n755_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n752_), .B1(new_n758_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n752_), .C1(new_n758_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  NAND3_X1  g566(.A1(new_n517_), .A2(new_n445_), .A3(new_n642_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n222_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n221_), .A2(new_n769_), .ZN(new_n770_));
  OAI221_X1 g569(.A(new_n233_), .B1(new_n228_), .B2(new_n769_), .C1(new_n770_), .C2(new_n227_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n236_), .A2(new_n771_), .A3(KEYINPUT116), .A4(new_n573_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n236_), .A2(new_n771_), .A3(new_n573_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n237_), .A2(new_n572_), .A3(new_n238_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n556_), .B1(new_n555_), .B2(new_n560_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n561_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n555_), .A2(KEYINPUT55), .A3(new_n556_), .A4(new_n560_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n569_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n772_), .B(new_n775_), .C1(new_n776_), .C2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(KEYINPUT57), .A3(new_n597_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n784_), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n597_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  OR3_X1    g589(.A1(new_n781_), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n781_), .A2(KEYINPUT56), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT117), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT118), .B1(new_n781_), .B2(KEYINPUT56), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n781_), .A2(new_n795_), .A3(KEYINPUT56), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n791_), .A2(new_n793_), .A3(new_n794_), .A4(new_n796_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n236_), .A2(new_n771_), .A3(new_n572_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n797_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n602_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n789_), .B1(new_n790_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n784_), .A2(new_n597_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n802_), .A2(new_n790_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n615_), .B1(new_n803_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n601_), .A2(new_n614_), .A3(new_n576_), .ZN(new_n809_));
  OR3_X1    g608(.A1(new_n809_), .A2(KEYINPUT54), .A3(new_n627_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT54), .B1(new_n809_), .B2(new_n627_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n768_), .B1(new_n808_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  INV_X1    g613(.A(new_n812_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n805_), .A2(new_n804_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n802_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT121), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT121), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n802_), .A2(new_n816_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n789_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n815_), .B1(new_n821_), .B2(new_n615_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n768_), .A2(KEYINPUT59), .ZN(new_n823_));
  OAI22_X1  g622(.A1(new_n813_), .A2(new_n814_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n239_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n813_), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n239_), .A2(G113gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(G1340gat));
  OAI21_X1  g627(.A(G120gat), .B1(new_n824_), .B2(new_n576_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT60), .ZN(new_n830_));
  AOI21_X1  g629(.A(G120gat), .B1(new_n674_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n830_), .B2(G120gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT122), .B1(new_n813_), .B2(new_n832_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n813_), .A2(KEYINPUT122), .A3(new_n832_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n829_), .B1(new_n833_), .B2(new_n834_), .ZN(G1341gat));
  OAI21_X1  g634(.A(G127gat), .B1(new_n824_), .B2(new_n615_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n615_), .A2(G127gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n826_), .B2(new_n837_), .ZN(G1342gat));
  OAI21_X1  g637(.A(G134gat), .B1(new_n824_), .B2(new_n601_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n597_), .A2(G134gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n826_), .B2(new_n840_), .ZN(G1343gat));
  AOI21_X1  g640(.A(new_n642_), .B1(new_n808_), .B2(new_n812_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n516_), .A2(new_n446_), .A3(new_n653_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n627_), .A3(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g644(.A1(new_n842_), .A2(new_n674_), .A3(new_n843_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g646(.A1(new_n842_), .A2(new_n614_), .A3(new_n843_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  NAND2_X1  g649(.A1(new_n842_), .A2(new_n843_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G162gat), .B1(new_n851_), .B2(new_n601_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n597_), .A2(G162gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n851_), .B2(new_n853_), .ZN(G1347gat));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n516_), .A2(new_n653_), .A3(new_n518_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n822_), .A2(new_n239_), .A3(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n855_), .B(new_n856_), .C1(new_n858_), .C2(new_n266_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n283_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n820_), .A2(new_n789_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n819_), .B1(new_n802_), .B2(new_n816_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n615_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n857_), .B1(new_n863_), .B2(new_n812_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n266_), .B1(new_n864_), .B2(new_n627_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT62), .B1(new_n865_), .B2(KEYINPUT123), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n858_), .A2(new_n855_), .A3(new_n266_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n859_), .B(new_n860_), .C1(new_n866_), .C2(new_n867_), .ZN(G1348gat));
  AOI21_X1  g667(.A(G176gat), .B1(new_n864_), .B2(new_n674_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n487_), .B1(new_n808_), .B2(new_n812_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n516_), .A2(new_n518_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n871_), .A2(new_n267_), .A3(new_n576_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n870_), .B2(new_n872_), .ZN(G1349gat));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  INV_X1    g673(.A(new_n365_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n864_), .A2(new_n875_), .A3(new_n614_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n871_), .A2(new_n615_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n870_), .A2(new_n877_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n874_), .B(new_n876_), .C1(new_n878_), .C2(new_n280_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n280_), .B1(new_n870_), .B2(new_n877_), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n822_), .A2(new_n365_), .A3(new_n615_), .A4(new_n857_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT124), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1350gat));
  NAND3_X1  g682(.A1(new_n864_), .A2(new_n622_), .A3(new_n366_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n822_), .A2(new_n601_), .A3(new_n857_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n255_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT125), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n884_), .B(new_n888_), .C1(new_n885_), .C2(new_n255_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1351gat));
  NOR3_X1   g689(.A1(new_n515_), .A2(new_n445_), .A3(new_n653_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n842_), .A2(G197gat), .A3(new_n627_), .A4(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n802_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n895_), .A2(KEYINPUT119), .B1(new_n787_), .B2(new_n788_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n614_), .B1(new_n896_), .B2(new_n806_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n320_), .B(new_n891_), .C1(new_n897_), .C2(new_n815_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n333_), .B1(new_n898_), .B2(new_n239_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n894_), .A2(new_n900_), .ZN(G1352gat));
  NOR2_X1   g700(.A1(new_n898_), .A2(new_n576_), .ZN(new_n902_));
  MUX2_X1   g701(.A(G204gat), .B(new_n343_), .S(new_n902_), .Z(G1353gat));
  NAND3_X1  g702(.A1(new_n842_), .A2(new_n614_), .A3(new_n891_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT63), .B(G211gat), .Z(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n904_), .B2(new_n906_), .ZN(G1354gat));
  OAI21_X1  g706(.A(G218gat), .B1(new_n898_), .B2(new_n601_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n622_), .A2(new_n326_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n898_), .B2(new_n909_), .ZN(G1355gat));
endmodule


