//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n833_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G8gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT75), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT76), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n207_), .B(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G231gat), .A2(G233gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n210_), .B(new_n211_), .Z(new_n212_));
  XNOR2_X1  g011(.A(G71gat), .B(G78gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(G57gat), .B(G64gat), .Z(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT11), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n213_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n213_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(new_n215_), .B2(KEYINPUT11), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n212_), .B(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G127gat), .B(G155gat), .ZN(new_n225_));
  INV_X1    g024(.A(G211gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT16), .B(G183gat), .Z(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT17), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n229_), .A2(KEYINPUT17), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n224_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT78), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n222_), .B(KEYINPUT68), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n212_), .B(new_n234_), .Z(new_n235_));
  XOR2_X1   g034(.A(new_n230_), .B(KEYINPUT77), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G15gat), .B(G43gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT79), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(G190gat), .ZN(new_n244_));
  INV_X1    g043(.A(G190gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(KEYINPUT79), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT26), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT80), .ZN(new_n248_));
  AND2_X1   g047(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT26), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G190gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n247_), .A2(new_n248_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT81), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT24), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n245_), .A2(KEYINPUT79), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n243_), .A2(G190gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n252_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n253_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT80), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n254_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT82), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n256_), .A2(KEYINPUT24), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT23), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT83), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n269_), .ZN(new_n273_));
  NOR3_X1   g072(.A1(new_n268_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT82), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n254_), .A2(new_n260_), .A3(new_n265_), .A4(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n267_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n271_), .B1(new_n273_), .B2(new_n272_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n269_), .A2(KEYINPUT83), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n244_), .A2(new_n246_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n278_), .B(new_n279_), .C1(G183gat), .C2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n257_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n277_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n277_), .B2(new_n286_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n242_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n288_), .A2(new_n289_), .A3(new_n242_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n241_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(G127gat), .A2(G134gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G127gat), .A2(G134gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(G113gat), .A2(G120gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G113gat), .A2(G120gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n295_), .A2(new_n298_), .A3(new_n296_), .A4(new_n299_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(KEYINPUT85), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(KEYINPUT85), .B2(new_n302_), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT31), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT86), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n291_), .A2(new_n241_), .A3(new_n292_), .ZN(new_n307_));
  OR3_X1    g106(.A1(new_n294_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n309_));
  OAI22_X1  g108(.A1(new_n307_), .A2(new_n294_), .B1(new_n309_), .B2(new_n305_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G141gat), .ZN(new_n312_));
  INV_X1    g111(.A(G148gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT3), .B1(new_n314_), .B2(KEYINPUT87), .ZN(new_n315_));
  AND3_X1   g114(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT87), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G155gat), .B(G162gat), .Z(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G155gat), .ZN(new_n325_));
  INV_X1    g124(.A(G162gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT1), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(G155gat), .A3(G162gat), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n327_), .B(new_n329_), .C1(G155gat), .C2(G162gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n314_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n324_), .A2(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(KEYINPUT29), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G22gat), .B(G50gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT28), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n334_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(KEYINPUT29), .ZN(new_n339_));
  OR2_X1    g138(.A1(G211gat), .A2(G218gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G211gat), .A2(G218gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(G197gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(G204gat), .ZN(new_n344_));
  INV_X1    g143(.A(G204gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n345_), .A2(G197gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT21), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT89), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n343_), .B2(G204gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n350_), .B2(new_n344_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n342_), .B(new_n347_), .C1(new_n351_), .C2(KEYINPUT21), .ZN(new_n352_));
  INV_X1    g151(.A(new_n341_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G211gat), .A2(G218gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT90), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT90), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n340_), .A2(new_n356_), .A3(new_n341_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(KEYINPUT21), .A3(new_n351_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n339_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(G228gat), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n352_), .A2(new_n359_), .A3(KEYINPUT91), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT91), .B1(new_n352_), .B2(new_n359_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n339_), .B(new_n365_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n367_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n372_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n338_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n337_), .A3(new_n373_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT24), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n255_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n278_), .A2(new_n279_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT94), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n258_), .B(KEYINPUT93), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT26), .B(G190gat), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n385_), .A2(new_n256_), .B1(new_n251_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT94), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n278_), .A2(new_n388_), .A3(new_n279_), .A4(new_n382_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n384_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n352_), .A2(new_n359_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n273_), .A2(new_n272_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(G183gat), .B2(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n285_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n395_), .A2(KEYINPUT20), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT91), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n360_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n352_), .A2(new_n359_), .A3(KEYINPUT91), .ZN(new_n399_));
  AOI221_X4 g198(.A(KEYINPUT96), .B1(new_n398_), .B2(new_n399_), .C1(new_n277_), .C2(new_n286_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n277_), .A2(new_n286_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n399_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n396_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT95), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n390_), .A2(new_n394_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(new_n360_), .ZN(new_n412_));
  AOI211_X1 g211(.A(KEYINPUT95), .B(new_n391_), .C1(new_n390_), .C2(new_n394_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n408_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n277_), .A2(new_n398_), .A3(new_n399_), .A4(new_n286_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n414_), .A2(KEYINPUT20), .A3(new_n415_), .A4(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n409_), .A2(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G64gat), .B(G92gat), .Z(new_n419_));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT32), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n418_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n301_), .A2(new_n302_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n324_), .A2(new_n428_), .A3(new_n332_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT98), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n304_), .A2(new_n333_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT98), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n324_), .A2(new_n332_), .A3(new_n432_), .A4(new_n428_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT4), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT4), .B1(new_n304_), .B2(new_n333_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(KEYINPUT99), .B(KEYINPUT0), .Z(new_n442_));
  XNOR2_X1  g241(.A(G1gat), .B(G29gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G57gat), .B(G85gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n444_), .B(new_n445_), .Z(new_n446_));
  OR2_X1    g245(.A1(new_n434_), .A2(new_n440_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n441_), .A2(KEYINPUT102), .A3(new_n446_), .A4(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n436_), .B1(new_n434_), .B2(KEYINPUT4), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n449_), .B2(new_n439_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n446_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT102), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n447_), .B(new_n446_), .C1(new_n449_), .C2(new_n439_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n411_), .A2(new_n360_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT95), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n411_), .A2(new_n410_), .A3(new_n360_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n456_), .A2(KEYINPUT20), .A3(new_n416_), .A4(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n408_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n415_), .B(new_n396_), .C1(new_n400_), .C2(new_n404_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n425_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n427_), .A2(new_n448_), .A3(new_n454_), .A4(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n453_), .A2(KEYINPUT100), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT100), .B1(new_n453_), .B2(new_n463_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n438_), .A2(KEYINPUT101), .A3(new_n439_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT101), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n449_), .B2(new_n440_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n434_), .A2(new_n439_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n451_), .A4(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n441_), .A2(KEYINPUT33), .A3(new_n446_), .A4(new_n447_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n459_), .A2(new_n460_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n423_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n459_), .A2(new_n460_), .A3(new_n424_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n466_), .A2(new_n473_), .A3(new_n475_), .A4(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n380_), .B1(new_n462_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n416_), .A2(KEYINPUT20), .ZN(new_n479_));
  NOR4_X1   g278(.A1(new_n479_), .A2(new_n412_), .A3(new_n413_), .A4(new_n408_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n408_), .B2(new_n405_), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT27), .B(new_n476_), .C1(new_n481_), .C2(new_n424_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT27), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n459_), .A2(new_n424_), .A3(new_n460_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n424_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n379_), .B1(new_n448_), .B2(new_n454_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n482_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n311_), .B1(new_n478_), .B2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n454_), .A2(new_n448_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n482_), .A2(new_n486_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n379_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n238_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G29gat), .B(G36gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G29gat), .B(G36gat), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n496_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n499_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n495_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n499_), .A2(new_n501_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n502_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n499_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(KEYINPUT15), .A3(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n505_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G85gat), .B(G92gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT65), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT6), .ZN(new_n517_));
  INV_X1    g316(.A(G99gat), .ZN(new_n518_));
  INV_X1    g317(.A(G106gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(KEYINPUT64), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT7), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT7), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n522_), .A2(new_n518_), .A3(new_n519_), .A4(KEYINPUT64), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n514_), .A2(new_n515_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n515_), .B1(new_n514_), .B2(new_n524_), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT10), .B(G99gat), .Z(new_n528_));
  AND2_X1   g327(.A1(new_n528_), .A2(new_n519_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT9), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(G85gat), .A3(G92gat), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n517_), .B(new_n531_), .C1(new_n530_), .C2(new_n512_), .ZN(new_n532_));
  OAI22_X1  g331(.A1(new_n526_), .A2(new_n527_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT73), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n511_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n505_), .A2(new_n510_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n532_), .A2(new_n529_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n514_), .A2(new_n524_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT8), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n539_), .B2(new_n525_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT73), .B1(new_n536_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n508_), .A2(new_n509_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n544_), .A2(KEYINPUT74), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT74), .B1(new_n544_), .B2(new_n549_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554_));
  XOR2_X1   g353(.A(G190gat), .B(G218gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n511_), .A2(new_n533_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n549_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n547_), .A2(new_n548_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n543_), .A4(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n553_), .A2(new_n554_), .A3(new_n557_), .A4(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n544_), .A2(new_n549_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT74), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(new_n550_), .A3(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n557_), .A2(new_n554_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n557_), .A2(new_n554_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n562_), .A2(new_n569_), .A3(KEYINPUT37), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT37), .B1(new_n562_), .B2(new_n569_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n494_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n533_), .A2(new_n223_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT67), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n540_), .A2(new_n222_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT66), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n575_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n234_), .A2(KEYINPUT12), .A3(new_n533_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n576_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT69), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n578_), .B2(new_n574_), .ZN(new_n586_));
  AOI211_X1 g385(.A(KEYINPUT69), .B(new_n575_), .C1(new_n540_), .C2(new_n222_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n582_), .B(new_n584_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(KEYINPUT70), .B(KEYINPUT5), .Z(new_n589_));
  XNOR2_X1  g388(.A(G120gat), .B(G148gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G176gat), .B(G204gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n581_), .A2(new_n588_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n581_), .B2(new_n588_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n597_), .A2(KEYINPUT13), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(KEYINPUT13), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n210_), .B(new_n542_), .Z(new_n601_));
  NAND2_X1  g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n511_), .A2(new_n210_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n210_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n542_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(new_n607_), .A3(new_n602_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n604_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G113gat), .B(G141gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G169gat), .B(G197gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n604_), .A2(new_n608_), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n600_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n573_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(new_n202_), .A3(new_n490_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT38), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n562_), .A2(new_n569_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT103), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT104), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n494_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n490_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n618_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n621_), .B1(new_n202_), .B2(new_n627_), .ZN(G1324gat));
  NOR2_X1   g427(.A1(new_n625_), .A2(new_n618_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n492_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n203_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT39), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n619_), .A2(new_n203_), .A3(new_n630_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n311_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n629_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT41), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n619_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1326gat));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n629_), .B2(new_n380_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT42), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n380_), .A2(new_n643_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT105), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n619_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(G1327gat));
  NAND2_X1  g448(.A1(new_n489_), .A2(new_n493_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(new_n623_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n600_), .A2(new_n617_), .A3(new_n238_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(G29gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n490_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  INV_X1    g456(.A(new_n572_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n650_), .B2(new_n658_), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT43), .B(new_n572_), .C1(new_n489_), .C2(new_n493_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n653_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT106), .B(new_n653_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n650_), .A2(new_n658_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT43), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n650_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n652_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT107), .B1(new_n670_), .B2(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n666_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n663_), .A2(KEYINPUT107), .A3(new_n664_), .A4(new_n665_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n626_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n656_), .B1(new_n674_), .B2(new_n655_), .ZN(G1328gat));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n672_), .A2(new_n673_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT108), .B1(new_n677_), .B2(new_n630_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n679_), .B(new_n492_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n680_));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n678_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n654_), .A2(new_n681_), .A3(new_n630_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT45), .Z(new_n684_));
  OAI21_X1  g483(.A(new_n676_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n677_), .A2(new_n630_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n679_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n677_), .A2(KEYINPUT108), .A3(new_n630_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(G36gat), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n684_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(KEYINPUT46), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n685_), .A2(new_n691_), .ZN(G1329gat));
  XOR2_X1   g491(.A(KEYINPUT109), .B(G43gat), .Z(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n654_), .B2(new_n638_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n311_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G43gat), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g496(.A(G50gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n654_), .A2(new_n698_), .A3(new_n380_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n379_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n698_), .ZN(G1331gat));
  INV_X1    g500(.A(new_n600_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n616_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n573_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n490_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n625_), .A2(new_n703_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n490_), .A2(G57gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n706_), .B2(new_n707_), .ZN(G1332gat));
  INV_X1    g507(.A(G64gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n706_), .B2(new_n630_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT48), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n704_), .A2(new_n709_), .A3(new_n630_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1333gat));
  INV_X1    g512(.A(G71gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n706_), .B2(new_n638_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT49), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n704_), .A2(new_n714_), .A3(new_n638_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1334gat));
  INV_X1    g517(.A(G78gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n706_), .B2(new_n380_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT50), .Z(new_n721_));
  NAND2_X1  g520(.A1(new_n380_), .A2(new_n719_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT110), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n704_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1335gat));
  INV_X1    g524(.A(new_n238_), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n726_), .B(new_n703_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(G85gat), .A3(new_n490_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n703_), .A2(new_n726_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n651_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(new_n626_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(G85gat), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT111), .ZN(G1336gat));
  INV_X1    g532(.A(new_n730_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G92gat), .B1(new_n734_), .B2(new_n630_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT112), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n630_), .A2(G92gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n727_), .B2(new_n737_), .ZN(G1337gat));
  AOI21_X1  g537(.A(new_n518_), .B1(new_n727_), .B2(new_n638_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n638_), .A2(new_n528_), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT113), .B(new_n739_), .C1(new_n734_), .C2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g541(.A(new_n519_), .B1(new_n727_), .B2(new_n380_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT52), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n734_), .A2(new_n519_), .A3(new_n380_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(G1339gat));
  NOR4_X1   g547(.A1(new_n702_), .A2(new_n658_), .A3(new_n617_), .A4(new_n238_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT54), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n582_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n752_));
  AOI22_X1  g551(.A1(new_n588_), .A2(new_n751_), .B1(new_n752_), .B2(new_n575_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n582_), .A2(new_n584_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n586_), .A2(new_n587_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(KEYINPUT115), .A4(KEYINPUT55), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n588_), .B2(new_n751_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n753_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n593_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT56), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(KEYINPUT56), .A3(new_n760_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(KEYINPUT116), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n759_), .A2(new_n765_), .A3(KEYINPUT56), .A4(new_n760_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n764_), .A2(new_n617_), .A3(new_n594_), .A4(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n601_), .A2(new_n602_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n605_), .A2(new_n607_), .A3(new_n603_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n612_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n768_), .A2(KEYINPUT117), .A3(new_n612_), .A4(new_n769_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(new_n615_), .A3(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n767_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n623_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n595_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT58), .A3(new_n774_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n763_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n594_), .B(new_n774_), .C1(new_n785_), .C2(new_n761_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(new_n658_), .A3(new_n788_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n780_), .A2(new_n781_), .B1(new_n782_), .B2(new_n789_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n789_), .A2(new_n782_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n623_), .B1(new_n767_), .B2(new_n777_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n792_), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT120), .B1(new_n792_), .B2(KEYINPUT57), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n790_), .B(new_n791_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n750_), .B1(new_n795_), .B2(new_n238_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NOR4_X1   g596(.A1(new_n630_), .A2(new_n311_), .A3(new_n626_), .A4(new_n380_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(G113gat), .B1(new_n800_), .B2(new_n617_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n780_), .A2(new_n781_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n789_), .B(new_n803_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n750_), .B1(new_n804_), .B2(new_n238_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n798_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT121), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n806_), .A2(KEYINPUT121), .A3(new_n807_), .A4(new_n798_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G113gat), .B1(new_n616_), .B2(KEYINPUT122), .ZN(new_n812_));
  AND4_X1   g611(.A1(new_n802_), .A2(new_n810_), .A3(new_n811_), .A4(new_n812_), .ZN(new_n813_));
  OR2_X1    g612(.A1(KEYINPUT122), .A2(G113gat), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n801_), .B1(new_n813_), .B2(new_n814_), .ZN(G1340gat));
  INV_X1    g614(.A(G120gat), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n600_), .B2(KEYINPUT60), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT123), .Z(new_n818_));
  OAI211_X1 g617(.A(new_n800_), .B(new_n818_), .C1(KEYINPUT60), .C2(new_n816_), .ZN(new_n819_));
  AND4_X1   g618(.A1(new_n702_), .A2(new_n810_), .A3(new_n802_), .A4(new_n811_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n816_), .ZN(G1341gat));
  AOI21_X1  g620(.A(G127gat), .B1(new_n800_), .B2(new_n726_), .ZN(new_n822_));
  AND4_X1   g621(.A1(G127gat), .A2(new_n810_), .A3(new_n802_), .A4(new_n811_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n726_), .ZN(G1342gat));
  INV_X1    g623(.A(new_n624_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G134gat), .B1(new_n800_), .B2(new_n825_), .ZN(new_n826_));
  AND4_X1   g625(.A1(new_n658_), .A2(new_n810_), .A3(new_n802_), .A4(new_n811_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g627(.A1(new_n796_), .A2(new_n379_), .A3(new_n638_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n630_), .A2(new_n626_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n617_), .A3(new_n830_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n702_), .A3(new_n830_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g633(.A1(new_n829_), .A2(new_n726_), .A3(new_n830_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT61), .B(G155gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1346gat));
  AND4_X1   g636(.A1(G162gat), .A2(new_n829_), .A3(new_n658_), .A4(new_n830_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n829_), .A2(new_n825_), .A3(new_n830_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n326_), .B2(new_n839_), .ZN(G1347gat));
  NAND3_X1  g639(.A1(new_n630_), .A2(new_n379_), .A3(new_n491_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n805_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n842_), .A2(new_n843_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n617_), .B(new_n283_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n842_), .A2(new_n617_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n848_), .A2(new_n849_), .A3(G169gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n848_), .B2(G169gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n847_), .B1(new_n850_), .B2(new_n851_), .ZN(G1348gat));
  NOR4_X1   g651(.A1(new_n796_), .A2(new_n284_), .A3(new_n600_), .A4(new_n841_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n702_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n284_), .ZN(G1349gat));
  NOR2_X1   g654(.A1(new_n796_), .A2(new_n841_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G183gat), .B1(new_n856_), .B2(new_n726_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n846_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n238_), .B1(new_n858_), .B2(new_n844_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n251_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n859_), .B2(new_n860_), .ZN(G1350gat));
  NAND2_X1  g660(.A1(new_n825_), .A2(new_n386_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT125), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n572_), .B1(new_n858_), .B2(new_n844_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n245_), .ZN(G1351gat));
  INV_X1    g665(.A(new_n487_), .ZN(new_n867_));
  NOR4_X1   g666(.A1(new_n796_), .A2(new_n867_), .A3(new_n492_), .A4(new_n638_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n617_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n702_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT126), .B(G204gat), .Z(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1353gat));
  NAND2_X1  g672(.A1(new_n795_), .A2(new_n238_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n750_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n638_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  AND4_X1   g675(.A1(new_n487_), .A2(new_n876_), .A3(new_n630_), .A4(new_n726_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT127), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT63), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n226_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n877_), .A2(new_n878_), .A3(new_n880_), .A4(new_n881_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n868_), .A2(new_n726_), .A3(new_n880_), .A4(new_n881_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT127), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n868_), .A2(new_n726_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n879_), .A3(new_n226_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n882_), .A2(new_n884_), .A3(new_n886_), .ZN(G1354gat));
  AOI21_X1  g686(.A(G218gat), .B1(new_n868_), .B2(new_n825_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n868_), .A2(new_n658_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(G218gat), .B2(new_n889_), .ZN(G1355gat));
endmodule


