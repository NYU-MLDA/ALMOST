//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n599_, new_n600_,
    new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n203_));
  NAND2_X1  g002(.A1(G232gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n205_), .A2(KEYINPUT35), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT7), .ZN(new_n207_));
  INV_X1    g006(.A(G99gat), .ZN(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(KEYINPUT65), .A3(new_n207_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(new_n213_), .B2(new_n207_), .ZN(new_n216_));
  OAI211_X1 g015(.A(KEYINPUT64), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n212_), .A2(new_n214_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  XOR2_X1   g024(.A(G85gat), .B(G92gat), .Z(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n220_), .A2(new_n222_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n232_), .B1(new_n218_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n212_), .A2(new_n214_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n216_), .A2(new_n217_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n235_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n228_), .B(new_n226_), .C1(new_n234_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT8), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n236_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT67), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n218_), .A2(new_n233_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n232_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n228_), .B1(new_n243_), .B2(new_n226_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n227_), .B1(new_n239_), .B2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT10), .B(G99gat), .Z(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n209_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n226_), .A2(KEYINPUT9), .ZN(new_n248_));
  INV_X1    g047(.A(G85gat), .ZN(new_n249_));
  INV_X1    g048(.A(G92gat), .ZN(new_n250_));
  OR3_X1    g049(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT9), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n247_), .A2(new_n248_), .A3(new_n223_), .A4(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n245_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G29gat), .B(G36gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G43gat), .B(G50gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT15), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT71), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n253_), .A2(new_n260_), .A3(new_n257_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n252_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n226_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT68), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT8), .A3(new_n238_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n263_), .B1(new_n266_), .B2(new_n227_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT72), .B1(new_n267_), .B2(new_n256_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n245_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n206_), .B1(new_n262_), .B2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G190gat), .B(G218gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(G134gat), .B(G162gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT36), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT73), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT74), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n269_), .B(new_n270_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT75), .B1(new_n205_), .B2(KEYINPUT35), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n206_), .B(new_n282_), .Z(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT76), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  OAI211_X1 g084(.A(KEYINPUT76), .B(new_n284_), .C1(new_n268_), .C2(new_n271_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n273_), .B(new_n280_), .C1(new_n285_), .C2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n276_), .B(KEYINPUT36), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n284_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n286_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n291_), .B1(new_n295_), .B2(new_n273_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n289_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT37), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n202_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n281_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n294_), .A2(new_n286_), .B1(new_n300_), .B2(new_n206_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n288_), .B1(new_n301_), .B2(new_n291_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(KEYINPUT77), .A3(KEYINPUT37), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n302_), .B2(KEYINPUT37), .ZN(new_n305_));
  INV_X1    g104(.A(new_n296_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n306_), .A2(KEYINPUT78), .A3(new_n298_), .A4(new_n288_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n299_), .A2(new_n303_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G15gat), .B(G22gat), .ZN(new_n309_));
  INV_X1    g108(.A(G1gat), .ZN(new_n310_));
  INV_X1    g109(.A(G8gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT14), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G8gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G231gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G57gat), .B(G64gat), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n318_), .A2(KEYINPUT11), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(KEYINPUT11), .ZN(new_n320_));
  XOR2_X1   g119(.A(G71gat), .B(G78gat), .Z(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n320_), .A2(new_n321_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n317_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G127gat), .B(G155gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT16), .ZN(new_n328_));
  XOR2_X1   g127(.A(G183gat), .B(G211gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OR3_X1    g130(.A1(new_n326_), .A2(KEYINPUT17), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(KEYINPUT79), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(KEYINPUT17), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n333_), .A2(new_n334_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n332_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT80), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT81), .B1(new_n308_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n305_), .A2(new_n307_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT77), .B1(new_n302_), .B2(KEYINPUT37), .ZN(new_n342_));
  INV_X1    g141(.A(new_n303_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n338_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT82), .ZN(new_n347_));
  AND2_X1   g146(.A1(G230gat), .A2(G233gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n267_), .A2(new_n324_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n267_), .A2(new_n324_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n348_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(new_n267_), .B2(new_n324_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n348_), .B1(new_n267_), .B2(new_n324_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n253_), .A2(KEYINPUT12), .A3(new_n325_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G120gat), .B(G148gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT5), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G176gat), .B(G204gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n352_), .A2(new_n357_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT13), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n363_), .A2(KEYINPUT13), .A3(new_n365_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n340_), .A2(new_n346_), .A3(new_n347_), .A4(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G78gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(G197gat), .B(G204gat), .Z(new_n374_));
  OR2_X1    g173(.A1(new_n374_), .A2(KEYINPUT21), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(KEYINPUT21), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n376_), .A2(new_n377_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G228gat), .A2(G233gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(KEYINPUT1), .ZN(new_n383_));
  OR2_X1    g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(KEYINPUT1), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n386_), .B2(new_n385_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT90), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n383_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n389_), .B2(new_n388_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G141gat), .A2(G148gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(KEYINPUT88), .Z(new_n393_));
  NOR2_X1   g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n394_), .B(KEYINPUT3), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(new_n393_), .B2(KEYINPUT2), .ZN(new_n398_));
  NAND3_X1  g197(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT91), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n382_), .B(new_n384_), .C1(new_n398_), .C2(new_n400_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n380_), .B(new_n381_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n396_), .B2(new_n401_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n380_), .B(KEYINPUT93), .ZN(new_n406_));
  OAI211_X1 g205(.A(G228gat), .B(G233gat), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n373_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n404_), .A2(new_n407_), .A3(new_n373_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(G106gat), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n410_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n209_), .B1(new_n412_), .B2(new_n408_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(KEYINPUT92), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT94), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT94), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n411_), .A2(new_n413_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n402_), .A2(new_n403_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT28), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G22gat), .B(G50gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n415_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n414_), .A3(KEYINPUT94), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G8gat), .B(G36gat), .Z(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G64gat), .B(G92gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT25), .B(G183gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT26), .B(G190gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n433_), .A2(KEYINPUT84), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G183gat), .A2(G190gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT85), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT23), .ZN(new_n437_));
  MUX2_X1   g236(.A(new_n435_), .B(new_n436_), .S(new_n437_), .Z(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(G169gat), .B2(G176gat), .ZN(new_n440_));
  NOR3_X1   g239(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(KEYINPUT84), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n434_), .A2(new_n438_), .A3(new_n442_), .A4(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n445_), .B1(new_n436_), .B2(KEYINPUT23), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(G183gat), .B2(G190gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(G169gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n444_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT20), .B1(new_n451_), .B2(new_n380_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n432_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n431_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(new_n446_), .A3(new_n442_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT96), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n438_), .B1(G183gat), .B2(G190gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n449_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n452_), .B1(new_n461_), .B2(new_n380_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n463_), .B(KEYINPUT19), .Z(new_n464_));
  AND2_X1   g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n406_), .A2(new_n460_), .A3(new_n456_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n451_), .B2(new_n380_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n464_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(KEYINPUT32), .B(new_n430_), .C1(new_n465_), .C2(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n470_), .A2(KEYINPUT101), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n462_), .A2(new_n464_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n458_), .A2(new_n378_), .A3(new_n379_), .A4(new_n460_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n430_), .A2(KEYINPUT32), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n470_), .A2(KEYINPUT101), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G127gat), .B(G134gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G113gat), .B(G120gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  AND3_X1   g280(.A1(new_n402_), .A2(KEYINPUT99), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n402_), .B2(KEYINPUT99), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT4), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G225gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT100), .ZN(new_n486_));
  INV_X1    g285(.A(new_n481_), .ZN(new_n487_));
  OR3_X1    g286(.A1(new_n402_), .A2(KEYINPUT4), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n484_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n482_), .A2(new_n483_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n485_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G1gat), .B(G29gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G85gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT0), .B(G57gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  NAND3_X1  g294(.A1(new_n489_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n495_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n471_), .B(new_n478_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT33), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n430_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n502_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT98), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n474_), .B(new_n430_), .C1(new_n462_), .C2(new_n464_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(KEYINPUT98), .B(new_n502_), .C1(new_n472_), .C2(new_n475_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n495_), .B1(new_n490_), .B2(new_n486_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n484_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n489_), .A2(new_n491_), .A3(KEYINPUT33), .A4(new_n495_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n501_), .A2(new_n508_), .A3(new_n511_), .A4(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n499_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n425_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT27), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n506_), .A2(new_n516_), .A3(new_n507_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n502_), .B1(new_n465_), .B2(new_n469_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(KEYINPUT27), .A3(new_n505_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n497_), .A2(new_n498_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n422_), .A2(new_n520_), .A3(new_n521_), .A4(new_n424_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G227gat), .A2(G233gat), .ZN(new_n524_));
  INV_X1    g323(.A(G71gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G99gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n451_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n481_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G15gat), .B(G43gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT86), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT30), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT31), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n529_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT87), .ZN(new_n535_));
  INV_X1    g334(.A(new_n520_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n536_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n521_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n534_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n523_), .A2(new_n535_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n257_), .A2(new_n315_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n315_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n256_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n315_), .B(new_n256_), .Z(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(G229gat), .A3(G233gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G113gat), .B(G141gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT83), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G169gat), .B(G197gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n548_), .A2(new_n550_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n541_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n372_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n340_), .A2(new_n346_), .A3(new_n371_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT82), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n562_), .A2(new_n310_), .A3(new_n564_), .A4(new_n538_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT38), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n522_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n422_), .A2(new_n424_), .B1(new_n499_), .B2(new_n513_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n535_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n537_), .A2(new_n540_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n370_), .A2(new_n560_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n297_), .A2(new_n339_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(G1gat), .B1(new_n575_), .B2(new_n521_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n565_), .A2(new_n566_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n567_), .A2(new_n576_), .A3(new_n577_), .ZN(G1324gat));
  OAI21_X1  g377(.A(G8gat), .B1(new_n575_), .B2(new_n520_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT39), .B1(new_n579_), .B2(KEYINPUT103), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT103), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n520_), .A2(G8gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n562_), .A2(new_n564_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT102), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT102), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n562_), .A2(new_n586_), .A3(new_n564_), .A4(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT40), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n582_), .A2(KEYINPUT40), .A3(new_n588_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(G1325gat));
  OAI21_X1  g392(.A(G15gat), .B1(new_n575_), .B2(new_n535_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT41), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n562_), .A2(new_n564_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n535_), .A2(G15gat), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(G1326gat));
  OAI21_X1  g397(.A(G22gat), .B1(new_n575_), .B2(new_n425_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT42), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n425_), .A2(G22gat), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n600_), .B1(new_n596_), .B2(new_n601_), .ZN(G1327gat));
  NAND2_X1  g401(.A1(new_n572_), .A2(new_n308_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT43), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n338_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n572_), .A2(KEYINPUT43), .A3(new_n308_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n573_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n605_), .A2(KEYINPUT44), .A3(new_n573_), .A4(new_n606_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(G29gat), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n521_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n297_), .A2(new_n339_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(new_n370_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n561_), .A2(new_n538_), .A3(new_n615_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n611_), .A2(new_n613_), .B1(new_n612_), .B2(new_n616_), .ZN(G1328gat));
  NAND3_X1  g416(.A1(new_n609_), .A2(new_n536_), .A3(new_n610_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(G36gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n561_), .A2(new_n615_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n520_), .A2(G36gat), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT105), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT105), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n561_), .A2(new_n624_), .A3(new_n615_), .A4(new_n621_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n623_), .A2(KEYINPUT45), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT45), .B1(new_n623_), .B2(new_n625_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n619_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT46), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n619_), .A2(new_n628_), .A3(KEYINPUT46), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1329gat));
  NAND4_X1  g432(.A1(new_n609_), .A2(G43gat), .A3(new_n534_), .A4(new_n610_), .ZN(new_n634_));
  INV_X1    g433(.A(G43gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n620_), .B2(new_n535_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n634_), .A2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g439(.A(new_n425_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n609_), .A2(G50gat), .A3(new_n641_), .A4(new_n610_), .ZN(new_n642_));
  INV_X1    g441(.A(G50gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(new_n620_), .B2(new_n425_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT107), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(G1331gat));
  NAND2_X1  g446(.A1(new_n370_), .A2(new_n560_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n541_), .A2(new_n648_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n649_), .A2(new_n340_), .A3(new_n346_), .ZN(new_n650_));
  INV_X1    g449(.A(G57gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n538_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n649_), .A2(new_n574_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G57gat), .B1(new_n653_), .B2(new_n521_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(G1332gat));
  OAI21_X1  g454(.A(G64gat), .B1(new_n653_), .B2(new_n520_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT108), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n658_), .B(G64gat), .C1(new_n653_), .C2(new_n520_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT48), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(G64gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n650_), .A2(new_n663_), .A3(new_n536_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n657_), .A2(KEYINPUT48), .A3(new_n659_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n662_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT109), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n662_), .A2(new_n668_), .A3(new_n664_), .A4(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1333gat));
  OAI21_X1  g469(.A(G71gat), .B1(new_n653_), .B2(new_n535_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT49), .ZN(new_n672_));
  INV_X1    g471(.A(new_n535_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n650_), .A2(new_n525_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1334gat));
  OAI21_X1  g474(.A(G78gat), .B1(new_n653_), .B2(new_n425_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT50), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n641_), .A2(new_n373_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT110), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n650_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n680_), .ZN(G1335gat));
  INV_X1    g480(.A(new_n614_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n649_), .A2(new_n682_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n683_), .A2(G85gat), .A3(new_n521_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n648_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n605_), .A2(new_n606_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n605_), .A2(KEYINPUT111), .A3(new_n606_), .A4(new_n686_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n521_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n685_), .B1(new_n691_), .B2(new_n249_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT112), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT112), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n694_), .B(new_n685_), .C1(new_n691_), .C2(new_n249_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1336gat));
  INV_X1    g495(.A(new_n683_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(new_n250_), .A3(new_n536_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n520_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n250_), .ZN(G1337gat));
  NAND3_X1  g499(.A1(new_n697_), .A2(new_n246_), .A3(new_n534_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n535_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(new_n208_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT51), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT51), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n705_), .B(new_n701_), .C1(new_n702_), .C2(new_n208_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1338gat));
  NAND3_X1  g506(.A1(new_n697_), .A2(new_n209_), .A3(new_n641_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n605_), .A2(new_n641_), .A3(new_n606_), .A4(new_n686_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(G106gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G106gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n713_), .B(new_n715_), .ZN(G1339gat));
  NAND4_X1  g515(.A1(new_n368_), .A2(new_n369_), .A3(new_n338_), .A4(new_n560_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT114), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n344_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT54), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT54), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n344_), .A2(new_n719_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n546_), .A2(KEYINPUT115), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n546_), .A2(KEYINPUT115), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n547_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n557_), .B1(new_n549_), .B2(new_n547_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n558_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(new_n365_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n357_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n354_), .A2(new_n349_), .A3(new_n356_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n348_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n354_), .A2(new_n355_), .A3(KEYINPUT55), .A4(new_n356_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(KEYINPUT56), .A3(new_n362_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT56), .B1(new_n738_), .B2(new_n362_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(KEYINPUT118), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT118), .ZN(new_n742_));
  AOI211_X1 g541(.A(new_n742_), .B(KEYINPUT56), .C1(new_n738_), .C2(new_n362_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n732_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT119), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT58), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT58), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(KEYINPUT119), .A3(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n308_), .A3(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n365_), .A2(new_n559_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n738_), .A2(KEYINPUT56), .A3(new_n362_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n740_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n730_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n297_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n758_), .B(new_n297_), .C1(new_n752_), .C2(new_n754_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n749_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n724_), .B1(new_n761_), .B2(new_n338_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT59), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n521_), .A2(new_n539_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n537_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n763_), .A3(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT117), .B1(new_n755_), .B2(new_n756_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  INV_X1    g568(.A(new_n756_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n738_), .A2(new_n362_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n739_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n753_), .B1(new_n774_), .B2(new_n750_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n769_), .B(new_n770_), .C1(new_n775_), .C2(new_n297_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n759_), .B1(new_n768_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n749_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT120), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n749_), .A3(KEYINPUT120), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n339_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n765_), .B1(new_n782_), .B2(new_n724_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n767_), .B1(new_n783_), .B2(new_n763_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G113gat), .B1(new_n784_), .B2(new_n560_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n781_), .A2(new_n339_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT120), .B1(new_n777_), .B2(new_n749_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n724_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n766_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n560_), .A2(G113gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n785_), .B1(new_n789_), .B2(new_n790_), .ZN(G1340gat));
  NOR2_X1   g590(.A1(new_n371_), .A2(KEYINPUT60), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT121), .B(G120gat), .Z(new_n793_));
  MUX2_X1   g592(.A(KEYINPUT60), .B(new_n792_), .S(new_n793_), .Z(new_n794_));
  NAND2_X1  g593(.A1(new_n783_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n723_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n722_), .B1(new_n344_), .B2(new_n719_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n338_), .B1(new_n749_), .B2(new_n760_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n766_), .A2(new_n763_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n370_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n789_), .B2(KEYINPUT59), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n795_), .B1(new_n803_), .B2(new_n793_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT122), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT122), .B(new_n795_), .C1(new_n803_), .C2(new_n793_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1341gat));
  INV_X1    g607(.A(G127gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n789_), .B2(new_n339_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n339_), .A2(new_n809_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n784_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT123), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n810_), .C1(new_n784_), .C2(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1342gat));
  OAI21_X1  g616(.A(G134gat), .B1(new_n784_), .B2(new_n344_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n302_), .A2(G134gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n789_), .B2(new_n819_), .ZN(G1343gat));
  NOR4_X1   g619(.A1(new_n425_), .A2(new_n536_), .A3(new_n521_), .A4(new_n673_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n788_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n559_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n370_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g626(.A1(new_n822_), .A2(new_n339_), .ZN(new_n828_));
  XOR2_X1   g627(.A(KEYINPUT61), .B(G155gat), .Z(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1346gat));
  OAI21_X1  g629(.A(G162gat), .B1(new_n822_), .B2(new_n344_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n302_), .A2(G162gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n822_), .B2(new_n832_), .ZN(G1347gat));
  INV_X1    g632(.A(G169gat), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n520_), .A2(new_n538_), .A3(new_n535_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n762_), .A2(new_n425_), .A3(new_n559_), .A4(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT62), .B(new_n834_), .C1(new_n836_), .C2(KEYINPUT22), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT62), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n425_), .B(new_n835_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n560_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT22), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n838_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G169gat), .B1(new_n836_), .B2(KEYINPUT62), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n837_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT124), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(new_n837_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1348gat));
  INV_X1    g647(.A(G176gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n839_), .B2(new_n371_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT125), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n641_), .B1(new_n782_), .B2(new_n724_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n835_), .A2(G176gat), .A3(new_n370_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1349gat));
  AND2_X1   g653(.A1(new_n835_), .A2(new_n338_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G183gat), .B1(new_n852_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n431_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n762_), .A2(new_n857_), .A3(new_n425_), .A4(new_n855_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n856_), .A2(new_n859_), .ZN(G1350gat));
  OAI21_X1  g659(.A(G190gat), .B1(new_n839_), .B2(new_n344_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n297_), .A2(new_n454_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n839_), .B2(new_n862_), .ZN(G1351gat));
  NOR4_X1   g662(.A1(new_n425_), .A2(new_n538_), .A3(new_n673_), .A4(new_n520_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n788_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n560_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT126), .B(G197gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1352gat));
  AND2_X1   g667(.A1(new_n788_), .A2(new_n864_), .ZN(new_n869_));
  INV_X1    g668(.A(G204gat), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n869_), .B(new_n370_), .C1(KEYINPUT127), .C2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(KEYINPUT127), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1353gat));
  NOR2_X1   g672(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n874_));
  AND2_X1   g673(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n875_));
  NOR4_X1   g674(.A1(new_n865_), .A2(new_n339_), .A3(new_n874_), .A4(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n869_), .A2(new_n338_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n874_), .ZN(G1354gat));
  OR3_X1    g677(.A1(new_n865_), .A2(G218gat), .A3(new_n302_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G218gat), .B1(new_n865_), .B2(new_n344_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1355gat));
endmodule


