//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT10), .B(G99gat), .Z(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT64), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(new_n215_), .B2(new_n214_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n210_), .B(new_n213_), .C1(new_n217_), .C2(new_n221_), .ZN(new_n222_));
  OR3_X1    g021(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n210_), .A2(new_n223_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT8), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n220_), .A2(new_n214_), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n222_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n205_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G232gat), .A2(G233gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT34), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT35), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n204_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n234_), .B(new_n239_), .C1(new_n233_), .C2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n237_), .A2(new_n238_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n241_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT36), .ZN(new_n245_));
  XOR2_X1   g044(.A(G134gat), .B(G162gat), .Z(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT73), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G190gat), .B(G218gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n244_), .A2(new_n245_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n245_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n244_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n254_), .B2(KEYINPUT74), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n241_), .B(new_n242_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n251_), .B(KEYINPUT36), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n256_), .A2(KEYINPUT74), .A3(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT37), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n257_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n252_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G15gat), .B(G22gat), .ZN(new_n265_));
  INV_X1    g064(.A(G1gat), .ZN(new_n266_));
  INV_X1    g065(.A(G8gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT14), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n265_), .B1(new_n268_), .B2(KEYINPUT76), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(KEYINPUT76), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G1gat), .B(G8gat), .ZN(new_n271_));
  OR3_X1    g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G57gat), .B(G64gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT11), .ZN(new_n276_));
  XOR2_X1   g075(.A(G71gat), .B(G78gat), .Z(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n276_), .A2(new_n277_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n275_), .A2(KEYINPUT11), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n274_), .B(new_n281_), .Z(new_n282_));
  NAND2_X1  g081(.A1(G231gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G127gat), .B(G155gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G183gat), .B(G211gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT17), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n289_), .A2(new_n290_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n284_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(new_n291_), .B2(new_n284_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT78), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n264_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT79), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n233_), .A2(KEYINPUT12), .A3(new_n281_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n233_), .A2(KEYINPUT67), .A3(KEYINPUT12), .A4(new_n281_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G230gat), .A2(G233gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT12), .B1(new_n233_), .B2(new_n281_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n233_), .A2(new_n281_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n303_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n304_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n306_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(new_n281_), .B2(new_n233_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n306_), .A2(new_n310_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n308_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G176gat), .B(G204gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G120gat), .B(G148gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n315_), .B(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n323_), .A2(KEYINPUT13), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(KEYINPUT13), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n298_), .A2(KEYINPUT80), .A3(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G8gat), .B(G36gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT101), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT19), .ZN(new_n335_));
  INV_X1    g134(.A(G197gat), .ZN(new_n336_));
  INV_X1    g135(.A(G204gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT21), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(KEYINPUT90), .B(G197gat), .Z(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n337_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT91), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT92), .B1(new_n336_), .B2(G204gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT90), .B(G197gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(new_n337_), .ZN(new_n345_));
  MUX2_X1   g144(.A(new_n343_), .B(KEYINPUT92), .S(new_n345_), .Z(new_n346_));
  OAI211_X1 g145(.A(new_n341_), .B(new_n342_), .C1(new_n346_), .C2(KEYINPUT21), .ZN(new_n347_));
  INV_X1    g146(.A(new_n342_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(KEYINPUT21), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT25), .B(G183gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G190gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT24), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(G169gat), .B2(G176gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(G169gat), .B2(G176gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n357_), .A2(KEYINPUT83), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(KEYINPUT83), .ZN(new_n359_));
  NOR3_X1   g158(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT23), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G183gat), .A3(G190gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n360_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n358_), .A2(new_n359_), .A3(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT84), .B(G176gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G169gat), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n367_), .A2(new_n368_), .B1(G169gat), .B2(G176gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(KEYINPUT85), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(new_n362_), .Z(new_n371_));
  NOR2_X1   g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n369_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n366_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n350_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n372_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n369_), .A2(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n357_), .A2(new_n360_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(new_n371_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n350_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n335_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n347_), .A2(new_n349_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n374_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n350_), .B2(new_n382_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n335_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n333_), .B1(new_n384_), .B2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n391_), .A2(new_n333_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n332_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n382_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT20), .B1(new_n385_), .B2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n350_), .A2(new_n374_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n335_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n385_), .A2(new_n395_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n335_), .A2(new_n388_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n375_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n331_), .A3(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n402_), .A2(KEYINPUT27), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n394_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n401_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n390_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n332_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n402_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT27), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT102), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT102), .ZN(new_n411_));
  AOI211_X1 g210(.A(new_n411_), .B(KEYINPUT27), .C1(new_n407_), .C2(new_n402_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n404_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G155gat), .B(G162gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT88), .ZN(new_n415_));
  OR2_X1    g214(.A1(G141gat), .A2(G148gat), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n416_), .A2(KEYINPUT3), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G141gat), .A2(G148gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT2), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n416_), .A2(KEYINPUT3), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n417_), .A2(new_n420_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n415_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G155gat), .ZN(new_n425_));
  INV_X1    g224(.A(G162gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT1), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(G155gat), .B2(G162gat), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT1), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n418_), .B(new_n416_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n430_), .ZN(new_n431_));
  OR3_X1    g230(.A1(new_n431_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT28), .B1(new_n431_), .B2(KEYINPUT29), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G22gat), .B(G50gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT94), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(KEYINPUT94), .A3(new_n438_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G228gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT89), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n431_), .A2(KEYINPUT29), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n444_), .B1(new_n385_), .B2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n447_));
  AOI21_X1  g246(.A(new_n444_), .B1(new_n431_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n350_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G78gat), .B(G106gat), .Z(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n446_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n441_), .B(new_n442_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n454_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n456_), .A2(new_n440_), .A3(new_n439_), .A4(new_n452_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G225gat), .A2(G233gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G127gat), .B(G134gat), .Z(new_n462_));
  XOR2_X1   g261(.A(G113gat), .B(G120gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT4), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT96), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n465_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT95), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n424_), .A2(new_n464_), .A3(new_n430_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n464_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n431_), .A2(KEYINPUT95), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n466_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n461_), .B1(new_n469_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n460_), .A3(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G1gat), .B(G29gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G57gat), .B(G85gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n479_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n477_), .A2(new_n484_), .A3(new_n478_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G71gat), .B(G99gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT86), .B(G43gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n374_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G227gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(G15gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT30), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n493_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n464_), .B(KEYINPUT31), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(KEYINPUT87), .A3(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n498_), .A2(KEYINPUT87), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(KEYINPUT87), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n499_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n489_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n413_), .A2(new_n459_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT98), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n398_), .A2(new_n401_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT99), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n398_), .A2(KEYINPUT99), .A3(new_n401_), .A4(new_n508_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n507_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n513_), .A2(new_n488_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n473_), .A2(new_n475_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n485_), .B1(new_n517_), .B2(new_n461_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n469_), .A2(new_n476_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n461_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(new_n407_), .A3(new_n402_), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT33), .B1(new_n479_), .B2(new_n485_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT33), .ZN(new_n523_));
  AOI211_X1 g322(.A(new_n523_), .B(new_n484_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n458_), .B1(new_n516_), .B2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n458_), .A2(new_n488_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n527_), .B(new_n404_), .C1(new_n410_), .C2(new_n412_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n504_), .A2(new_n501_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n506_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n205_), .A2(new_n274_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n274_), .A2(new_n240_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT81), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n204_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n538_));
  OAI211_X1 g337(.A(G229gat), .B(G233gat), .C1(new_n533_), .C2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G169gat), .B(G197gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n539_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT82), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n537_), .A2(new_n539_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n544_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n531_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n327_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT80), .B1(new_n298_), .B2(new_n326_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(new_n266_), .A3(new_n488_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT38), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n261_), .B(KEYINPUT103), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n531_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n326_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n296_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n549_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(G1gat), .B1(new_n562_), .B2(new_n489_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n554_), .A2(new_n555_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n556_), .A2(new_n563_), .A3(new_n564_), .ZN(G1324gat));
  NAND3_X1  g364(.A1(new_n553_), .A2(new_n267_), .A3(new_n413_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n558_), .A2(new_n413_), .A3(new_n561_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n267_), .B1(KEYINPUT104), .B2(KEYINPUT39), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n568_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n566_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g373(.A(G15gat), .B1(new_n562_), .B2(new_n530_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT41), .Z(new_n576_));
  INV_X1    g375(.A(new_n530_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n553_), .A2(new_n495_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(G1326gat));
  OAI21_X1  g378(.A(G22gat), .B1(new_n562_), .B2(new_n458_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT42), .ZN(new_n581_));
  INV_X1    g380(.A(G22gat), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n553_), .A2(new_n582_), .A3(new_n459_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(G1327gat));
  INV_X1    g383(.A(new_n261_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n296_), .A2(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n326_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n550_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(G29gat), .B1(new_n589_), .B2(new_n488_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n326_), .A2(new_n560_), .A3(new_n548_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT43), .B1(new_n264_), .B2(KEYINPUT105), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n531_), .B2(new_n264_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n264_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n577_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n595_), .B(new_n592_), .C1(new_n596_), .C2(new_n506_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n591_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(KEYINPUT44), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT44), .ZN(new_n600_));
  AOI211_X1 g399(.A(new_n600_), .B(new_n591_), .C1(new_n594_), .C2(new_n597_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n488_), .A2(G29gat), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n590_), .B1(new_n602_), .B2(new_n603_), .ZN(G1328gat));
  XOR2_X1   g403(.A(new_n413_), .B(KEYINPUT106), .Z(new_n605_));
  INV_X1    g404(.A(G36gat), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n588_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT45), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n407_), .A2(new_n402_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n411_), .B1(new_n611_), .B2(KEYINPUT27), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n408_), .A2(KEYINPUT102), .A3(new_n409_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n612_), .A2(new_n613_), .B1(new_n394_), .B2(new_n403_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n599_), .A2(new_n601_), .A3(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n610_), .B1(new_n615_), .B2(new_n606_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI221_X1 g417(.A(new_n610_), .B1(KEYINPUT107), .B2(KEYINPUT46), .C1(new_n615_), .C2(new_n606_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1329gat));
  AOI21_X1  g419(.A(G43gat), .B1(new_n589_), .B2(new_n577_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n577_), .A2(G43gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n602_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT47), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(G1330gat));
  AOI21_X1  g424(.A(G50gat), .B1(new_n589_), .B2(new_n459_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n459_), .A2(G50gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n602_), .B2(new_n627_), .ZN(G1331gat));
  NOR3_X1   g427(.A1(new_n531_), .A2(new_n326_), .A3(new_n548_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n298_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(G57gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(new_n488_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n505_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n614_), .A2(new_n634_), .A3(new_n458_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n522_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n479_), .A2(KEYINPUT33), .A3(new_n485_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n636_), .A2(new_n611_), .A3(new_n520_), .A4(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n513_), .A2(new_n488_), .A3(new_n515_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AOI22_X1  g439(.A1(new_n614_), .A2(new_n527_), .B1(new_n640_), .B2(new_n458_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n635_), .B1(new_n641_), .B2(new_n577_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n557_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n326_), .A2(new_n560_), .A3(new_n548_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT108), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT108), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n558_), .A2(new_n647_), .A3(new_n644_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(new_n488_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n633_), .B1(new_n650_), .B2(new_n632_), .ZN(G1332gat));
  INV_X1    g450(.A(G64gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n631_), .A2(new_n652_), .A3(new_n605_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n605_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G64gat), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n655_), .A2(KEYINPUT48), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(KEYINPUT48), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(G1333gat));
  NOR2_X1   g457(.A1(new_n530_), .A2(G71gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT109), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n631_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n646_), .A2(new_n648_), .A3(new_n577_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT49), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n662_), .A2(new_n663_), .A3(G71gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n662_), .B2(G71gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT110), .B(new_n661_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1334gat));
  OR3_X1    g469(.A1(new_n630_), .A2(G78gat), .A3(new_n458_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n649_), .A2(new_n459_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G78gat), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n673_), .A2(KEYINPUT50), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(KEYINPUT50), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(G1335gat));
  NAND2_X1  g475(.A1(new_n629_), .A2(new_n586_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n218_), .B1(new_n677_), .B2(new_n489_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT111), .Z(new_n679_));
  NOR3_X1   g478(.A1(new_n326_), .A2(new_n296_), .A3(new_n548_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n489_), .A2(new_n218_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n679_), .B1(new_n682_), .B2(new_n683_), .ZN(G1336gat));
  INV_X1    g483(.A(new_n677_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n219_), .A3(new_n413_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n682_), .A2(new_n605_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n687_), .B2(new_n219_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT112), .ZN(G1337gat));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n211_), .A3(new_n577_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n682_), .A2(new_n577_), .ZN(new_n691_));
  INV_X1    g490(.A(G99gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g493(.A(new_n592_), .B1(new_n642_), .B2(new_n595_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n597_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n459_), .B(new_n680_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT113), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(G106gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n697_), .B2(G106gat), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT52), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n699_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n458_), .B(new_n681_), .C1(new_n594_), .C2(new_n597_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT113), .B(new_n701_), .C1(new_n703_), .C2(new_n212_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n685_), .A2(new_n212_), .A3(new_n459_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT53), .B1(new_n702_), .B2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT113), .B1(new_n703_), .B2(new_n212_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n697_), .A2(new_n698_), .A3(G106gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(KEYINPUT52), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT53), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n704_), .A4(new_n705_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n707_), .A2(new_n712_), .ZN(G1339gat));
  NOR4_X1   g512(.A1(new_n413_), .A2(new_n530_), .A3(new_n489_), .A4(new_n459_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n315_), .A2(new_n322_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n548_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT56), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n322_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AND4_X1   g519(.A1(KEYINPUT55), .A2(new_n303_), .A3(new_n304_), .A4(new_n307_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n722_));
  AOI22_X1  g521(.A1(new_n301_), .A2(new_n302_), .B1(new_n306_), .B2(new_n305_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n304_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n721_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n303_), .A2(new_n307_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(KEYINPUT115), .A3(new_n309_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT115), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n728_), .B1(new_n723_), .B2(new_n304_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n720_), .B1(new_n725_), .B2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n322_), .B1(new_n725_), .B2(new_n730_), .ZN(new_n732_));
  OAI22_X1  g531(.A1(KEYINPUT116), .A2(new_n731_), .B1(new_n732_), .B2(KEYINPUT56), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT115), .B1(new_n726_), .B2(new_n309_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n723_), .A2(new_n728_), .A3(new_n304_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n723_), .A2(KEYINPUT55), .A3(new_n304_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n308_), .B2(new_n722_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n719_), .B1(new_n736_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT116), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n717_), .B1(new_n733_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT117), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n322_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n745_), .B1(new_n736_), .B2(new_n738_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n718_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n739_), .A2(new_n740_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n731_), .A2(KEYINPUT116), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(KEYINPUT117), .A3(new_n717_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n536_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n532_), .A2(new_n534_), .A3(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n536_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n546_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n543_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n323_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n744_), .A2(new_n751_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n261_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n716_), .A2(new_n756_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n732_), .A2(KEYINPUT56), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n731_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT58), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(KEYINPUT58), .B(new_n762_), .C1(new_n763_), .C2(new_n731_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n595_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n761_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT57), .B1(new_n758_), .B2(new_n585_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n560_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n326_), .A2(new_n296_), .A3(new_n264_), .A4(new_n549_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n715_), .B1(new_n772_), .B2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(G113gat), .B1(new_n777_), .B2(new_n548_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n750_), .A2(KEYINPUT117), .A3(new_n717_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT117), .B1(new_n750_), .B2(new_n717_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n757_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n759_), .B1(new_n783_), .B2(new_n261_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n768_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n296_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n779_), .B(new_n714_), .C1(new_n786_), .C2(new_n775_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n772_), .A2(new_n776_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n790_), .A2(new_n779_), .A3(KEYINPUT59), .A4(new_n714_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n549_), .A2(KEYINPUT119), .ZN(new_n793_));
  MUX2_X1   g592(.A(KEYINPUT119), .B(new_n793_), .S(G113gat), .Z(new_n794_));
  AOI21_X1  g593(.A(new_n778_), .B1(new_n792_), .B2(new_n794_), .ZN(G1340gat));
  NAND2_X1  g594(.A1(new_n790_), .A2(new_n714_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT120), .B(G120gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT60), .B1(new_n559_), .B2(new_n797_), .ZN(new_n798_));
  OR3_X1    g597(.A1(new_n796_), .A2(KEYINPUT60), .A3(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n559_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n801_), .B2(new_n797_), .ZN(G1341gat));
  INV_X1    g601(.A(G127gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n777_), .A2(new_n803_), .A3(new_n296_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n560_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n803_), .ZN(G1342gat));
  INV_X1    g605(.A(G134gat), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n264_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT59), .B1(new_n777_), .B2(new_n779_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n782_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n261_), .B1(new_n810_), .B2(new_n751_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n761_), .B(new_n769_), .C1(new_n811_), .C2(KEYINPUT57), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n775_), .B1(new_n812_), .B2(new_n560_), .ZN(new_n813_));
  NOR4_X1   g612(.A1(new_n813_), .A2(KEYINPUT118), .A3(new_n788_), .A4(new_n715_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n808_), .B1(new_n809_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  AOI21_X1  g615(.A(G134gat), .B1(new_n777_), .B2(new_n557_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n808_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT121), .B1(new_n821_), .B2(new_n817_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n822_), .ZN(G1343gat));
  NOR3_X1   g622(.A1(new_n605_), .A2(new_n489_), .A3(new_n458_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n790_), .A2(new_n530_), .A3(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n549_), .ZN(new_n826_));
  XOR2_X1   g625(.A(KEYINPUT122), .B(G141gat), .Z(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1344gat));
  NOR2_X1   g627(.A1(new_n825_), .A2(new_n326_), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(G148gat), .Z(G1345gat));
  OAI21_X1  g629(.A(KEYINPUT123), .B1(new_n825_), .B2(new_n560_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n813_), .A2(new_n577_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n296_), .A4(new_n824_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT61), .B(G155gat), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n831_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1346gat));
  OAI21_X1  g639(.A(G162gat), .B1(new_n825_), .B2(new_n264_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n557_), .A2(new_n426_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n825_), .B2(new_n842_), .ZN(G1347gat));
  AND3_X1   g642(.A1(new_n605_), .A2(new_n458_), .A3(new_n634_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n790_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G169gat), .B1(new_n845_), .B2(new_n549_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n845_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(new_n368_), .A3(new_n548_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n847_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(new_n850_), .A3(new_n851_), .ZN(G1348gat));
  NOR2_X1   g651(.A1(new_n845_), .A2(new_n326_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(G176gat), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(G176gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT124), .ZN(new_n857_));
  INV_X1    g656(.A(new_n367_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n853_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n857_), .B2(new_n859_), .ZN(G1349gat));
  NOR2_X1   g659(.A1(new_n845_), .A2(new_n560_), .ZN(new_n861_));
  MUX2_X1   g660(.A(G183gat), .B(new_n351_), .S(new_n861_), .Z(G1350gat));
  OAI21_X1  g661(.A(G190gat), .B1(new_n845_), .B2(new_n264_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n557_), .A2(new_n352_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n845_), .B2(new_n864_), .ZN(G1351gat));
  XNOR2_X1  g664(.A(KEYINPUT126), .B(G197gat), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n605_), .A2(new_n527_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n530_), .B(new_n867_), .C1(new_n786_), .C2(new_n775_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT125), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n790_), .A2(new_n870_), .A3(new_n530_), .A4(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n866_), .B1(new_n872_), .B2(new_n548_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n336_), .A2(KEYINPUT126), .ZN(new_n874_));
  AOI211_X1 g673(.A(new_n549_), .B(new_n874_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1352gat));
  AOI21_X1  g675(.A(new_n326_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT127), .B(G204gat), .Z(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n877_), .B2(new_n880_), .ZN(G1353gat));
  NOR2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  AND2_X1   g681(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n872_), .B(new_n296_), .C1(new_n882_), .C2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n560_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n882_), .ZN(G1354gat));
  INV_X1    g685(.A(G218gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n872_), .A2(new_n887_), .A3(new_n557_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n264_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n887_), .ZN(G1355gat));
endmodule


