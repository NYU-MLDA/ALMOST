//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT35), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n207_));
  AND3_X1   g006(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  OR3_X1    g010(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n210_), .A2(KEYINPUT66), .A3(new_n211_), .A4(new_n212_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n215_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n213_), .A2(new_n219_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT68), .B1(new_n223_), .B2(KEYINPUT8), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  AOI211_X1 g025(.A(new_n225_), .B(new_n226_), .C1(new_n213_), .C2(new_n219_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n222_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT10), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(G99gat), .ZN(new_n232_));
  INV_X1    g031(.A(G99gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(KEYINPUT10), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n230_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(KEYINPUT10), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(G99gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(KEYINPUT64), .ZN(new_n238_));
  AOI21_X1  g037(.A(G106gat), .B1(new_n235_), .B2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(G85gat), .A2(G92gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(KEYINPUT9), .A3(new_n216_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT9), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(G85gat), .A3(G92gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n210_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n229_), .B1(new_n239_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G106gat), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n236_), .A2(new_n237_), .A3(KEYINPUT64), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT64), .B1(new_n236_), .B2(new_n237_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n217_), .A2(new_n218_), .A3(new_n242_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT6), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n243_), .A3(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n249_), .A2(KEYINPUT65), .A3(new_n256_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n245_), .A2(KEYINPUT69), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT69), .B1(new_n245_), .B2(new_n257_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n228_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(KEYINPUT70), .B(new_n228_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G29gat), .B(G36gat), .ZN(new_n265_));
  INV_X1    g064(.A(G43gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G50gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n265_), .B(G43gat), .ZN(new_n269_));
  INV_X1    g068(.A(G50gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT15), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n207_), .B1(new_n264_), .B2(new_n274_), .ZN(new_n275_));
  AOI211_X1 g074(.A(KEYINPUT73), .B(new_n273_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n228_), .A2(new_n257_), .A3(new_n245_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(new_n272_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n206_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n263_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n239_), .A2(new_n229_), .A3(new_n244_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT65), .B1(new_n249_), .B2(new_n256_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n245_), .A2(KEYINPUT69), .A3(new_n257_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT70), .B1(new_n287_), .B2(new_n228_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n274_), .B1(new_n281_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT73), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n264_), .A2(new_n207_), .A3(new_n274_), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n206_), .B(KEYINPUT74), .Z(new_n292_));
  NAND4_X1  g091(.A1(new_n290_), .A2(new_n279_), .A3(new_n291_), .A4(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n204_), .A2(new_n205_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n280_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G190gat), .B(G218gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(G134gat), .ZN(new_n298_));
  INV_X1    g097(.A(G162gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(KEYINPUT36), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(KEYINPUT36), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  OAI211_X1 g104(.A(KEYINPUT75), .B(new_n302_), .C1(new_n280_), .C2(new_n295_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n290_), .A2(new_n279_), .A3(new_n291_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n206_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(new_n294_), .A3(new_n293_), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT75), .B1(new_n311_), .B2(new_n302_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n305_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT37), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(KEYINPUT37), .B(new_n305_), .C1(new_n307_), .C2(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G15gat), .B(G22gat), .ZN(new_n318_));
  INV_X1    g117(.A(G1gat), .ZN(new_n319_));
  INV_X1    g118(.A(G8gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT14), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G8gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT76), .B(KEYINPUT77), .Z(new_n325_));
  NAND2_X1  g124(.A1(G231gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n324_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G57gat), .B(G64gat), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n329_), .A2(KEYINPUT11), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(KEYINPUT11), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G71gat), .B(G78gat), .ZN(new_n332_));
  OR3_X1    g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n329_), .A2(new_n332_), .A3(KEYINPUT11), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n328_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT16), .B(G183gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G211gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G127gat), .B(G155gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n337_), .B1(KEYINPUT71), .B2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n341_), .B(KEYINPUT17), .Z(new_n345_));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n336_), .B(new_n345_), .C1(new_n346_), .C2(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n317_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT94), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT91), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G155gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(new_n299_), .ZN(new_n359_));
  INV_X1    g158(.A(G141gat), .ZN(new_n360_));
  INV_X1    g159(.A(G148gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT2), .B1(new_n362_), .B2(KEYINPUT93), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT93), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n364_), .B(new_n365_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n363_), .A2(new_n366_), .A3(new_n367_), .A4(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n354_), .B1(new_n359_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n359_), .A2(new_n354_), .A3(new_n371_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT92), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT1), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n357_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n358_), .A2(new_n299_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n357_), .A2(new_n377_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n362_), .A2(new_n368_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n376_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n380_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n376_), .B(new_n383_), .C1(new_n385_), .C2(new_n378_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n375_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT90), .B(G113gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G120gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(G127gat), .B(G134gat), .Z(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(KEYINPUT102), .A3(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n383_), .B1(new_n385_), .B2(new_n378_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT92), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n395_), .A2(new_n386_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n392_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n353_), .B1(new_n393_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n396_), .A2(new_n397_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT4), .B1(new_n400_), .B2(KEYINPUT102), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n352_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n396_), .B(new_n392_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n351_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G57gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G85gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(G1gat), .B(G29gat), .Z(new_n408_));
  XOR2_X1   g207(.A(new_n407_), .B(new_n408_), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT106), .ZN(new_n411_));
  INV_X1    g210(.A(new_n409_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n402_), .A2(KEYINPUT105), .A3(new_n404_), .A4(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n402_), .A2(new_n404_), .A3(new_n412_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT105), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT106), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n405_), .A2(new_n417_), .A3(new_n409_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n411_), .A2(new_n413_), .A3(new_n416_), .A4(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT18), .B(G64gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G92gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  AND2_X1   g222(.A1(new_n423_), .A2(KEYINPUT32), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT19), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G197gat), .B(G204gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT21), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G211gat), .B(G218gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n429_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT95), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n430_), .A2(new_n431_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT22), .B(G169gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n438_), .B(KEYINPUT101), .Z(new_n439_));
  INV_X1    g238(.A(G176gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G183gat), .ZN(new_n442_));
  INV_X1    g241(.A(G190gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT23), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT86), .ZN(new_n445_));
  OR3_X1    g244(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT23), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n443_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n447_), .A2(new_n448_), .B1(G169gat), .B2(G176gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT25), .B(G183gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT26), .B(G190gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G169gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n440_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G169gat), .A2(G176gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT24), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT100), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n446_), .A2(new_n444_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n454_), .A2(KEYINPUT24), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n441_), .A2(new_n449_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n427_), .B1(new_n437_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n447_), .A2(new_n464_), .A3(new_n460_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n464_), .B1(new_n447_), .B2(new_n460_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n452_), .B(KEYINPUT84), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n456_), .B(KEYINPUT85), .Z(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n466_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n459_), .A2(new_n448_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n438_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n455_), .B1(new_n473_), .B2(G176gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n436_), .B1(new_n471_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n426_), .B1(new_n463_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n475_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n467_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n480_), .A2(new_n469_), .A3(new_n468_), .A4(new_n465_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n437_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n449_), .A2(new_n441_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n458_), .A2(new_n461_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n436_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n482_), .A2(new_n485_), .A3(KEYINPUT20), .A4(new_n426_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n424_), .B1(new_n478_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n463_), .A2(new_n476_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n426_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n485_), .A3(KEYINPUT20), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n489_), .B1(new_n426_), .B2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n487_), .B1(new_n491_), .B2(new_n424_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n419_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n486_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n423_), .B1(new_n494_), .B2(new_n477_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n423_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n478_), .A2(new_n496_), .A3(new_n486_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n351_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n403_), .A2(new_n352_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n409_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT104), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n499_), .A2(KEYINPUT104), .A3(new_n500_), .A4(new_n409_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n498_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT33), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n414_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n414_), .A2(new_n506_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT103), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n414_), .A2(KEYINPUT103), .A3(new_n506_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n505_), .A2(new_n507_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n493_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G43gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G227gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G71gat), .B(G99gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT30), .B1(new_n471_), .B2(new_n475_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n481_), .A2(new_n520_), .A3(new_n479_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT89), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n521_), .A3(new_n518_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT88), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n392_), .B(KEYINPUT31), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n523_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT98), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n388_), .A2(KEYINPUT29), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G228gat), .A2(G233gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n436_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT96), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT96), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n531_), .A2(new_n535_), .A3(new_n436_), .A4(new_n532_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT29), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n538_), .B1(new_n396_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n388_), .A2(KEYINPUT97), .A3(KEYINPUT29), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(new_n541_), .A3(new_n436_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(G228gat), .A3(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G78gat), .B(G106gat), .Z(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n530_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n396_), .A2(new_n539_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G22gat), .B(G50gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT28), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n548_), .B(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n551_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n537_), .A2(new_n543_), .A3(KEYINPUT98), .A4(new_n545_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT99), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n544_), .B1(new_n555_), .B2(new_n545_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n537_), .A2(KEYINPUT99), .A3(new_n543_), .A4(new_n546_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n551_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n513_), .A2(new_n529_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT27), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n478_), .A2(new_n486_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(new_n423_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n491_), .A2(new_n496_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n563_), .A2(new_n564_), .A3(KEYINPUT107), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT107), .B1(new_n563_), .B2(new_n564_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT27), .B1(new_n495_), .B2(new_n497_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n419_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n529_), .A2(new_n554_), .A3(new_n558_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n527_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n528_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n554_), .A2(new_n558_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n568_), .B(new_n569_), .C1(new_n570_), .C2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n560_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n350_), .A2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n273_), .A2(new_n324_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n268_), .A2(new_n271_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n324_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT79), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n580_), .B1(new_n324_), .B2(new_n578_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT80), .ZN(new_n586_));
  INV_X1    g385(.A(new_n582_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n584_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT80), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n585_), .B(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n583_), .B(new_n593_), .C1(new_n596_), .C2(new_n582_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT83), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(KEYINPUT83), .A3(new_n593_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n594_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n335_), .B(KEYINPUT71), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n264_), .A2(KEYINPUT12), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604_));
  INV_X1    g403(.A(new_n335_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n278_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n278_), .A2(new_n605_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .A4(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n607_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(G230gat), .A3(G233gat), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(G120gat), .B(G148gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n610_), .A2(new_n612_), .A3(new_n618_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT13), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n620_), .A2(KEYINPUT13), .A3(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n601_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n576_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n319_), .A3(new_n419_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT38), .ZN(new_n631_));
  INV_X1    g430(.A(new_n313_), .ZN(new_n632_));
  AOI211_X1 g431(.A(new_n349_), .B(new_n632_), .C1(new_n574_), .C2(new_n560_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n627_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n634_), .B2(new_n569_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n631_), .A2(new_n635_), .ZN(G1324gat));
  OAI21_X1  g435(.A(G8gat), .B1(new_n634_), .B2(new_n568_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT39), .ZN(new_n638_));
  INV_X1    g437(.A(new_n568_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n629_), .A2(new_n320_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g441(.A(G15gat), .B1(new_n634_), .B2(new_n529_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT41), .Z(new_n644_));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n529_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n629_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(G1326gat));
  INV_X1    g447(.A(G22gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n559_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n629_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G22gat), .B1(new_n634_), .B2(new_n559_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(KEYINPUT108), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(KEYINPUT108), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(KEYINPUT42), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT42), .B1(new_n653_), .B2(new_n654_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n651_), .B1(new_n655_), .B2(new_n656_), .ZN(G1327gat));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n575_), .A2(new_n658_), .A3(new_n317_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT109), .ZN(new_n660_));
  INV_X1    g459(.A(new_n316_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n302_), .B1(new_n280_), .B2(new_n295_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT75), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n306_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT37), .B1(new_n665_), .B2(new_n305_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n660_), .B1(new_n661_), .B2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n315_), .A2(KEYINPUT109), .A3(new_n316_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n667_), .A2(new_n668_), .B1(new_n574_), .B2(new_n560_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n659_), .B1(new_n669_), .B2(new_n658_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n628_), .A2(new_n348_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT110), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n672_), .B(new_n674_), .Z(new_n675_));
  OAI21_X1  g474(.A(G29gat), .B1(new_n675_), .B2(new_n569_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n313_), .B1(new_n560_), .B2(new_n574_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n671_), .ZN(new_n678_));
  OR3_X1    g477(.A1(new_n678_), .A2(G29gat), .A3(new_n569_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT111), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT111), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n676_), .A2(new_n682_), .A3(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1328gat));
  OAI21_X1  g483(.A(G36gat), .B1(new_n675_), .B2(new_n568_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n678_), .A2(G36gat), .A3(new_n568_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n685_), .B(new_n688_), .C1(KEYINPUT113), .C2(KEYINPUT46), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  OAI21_X1  g492(.A(G43gat), .B1(new_n675_), .B2(new_n529_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n678_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n266_), .A3(new_n646_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n694_), .A2(KEYINPUT47), .A3(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1330gat));
  OAI21_X1  g500(.A(G50gat), .B1(new_n675_), .B2(new_n559_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n695_), .A2(new_n270_), .A3(new_n650_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1331gat));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n419_), .B2(KEYINPUT114), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n633_), .A2(new_n601_), .A3(new_n626_), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n706_), .B(new_n707_), .C1(KEYINPUT114), .C2(new_n705_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n601_), .A2(new_n626_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n576_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n419_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n708_), .A2(new_n711_), .ZN(G1332gat));
  OAI21_X1  g511(.A(G64gat), .B1(new_n707_), .B2(new_n568_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT48), .ZN(new_n714_));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n710_), .A2(new_n715_), .A3(new_n639_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n707_), .B2(new_n529_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT49), .ZN(new_n719_));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n710_), .A2(new_n720_), .A3(new_n646_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1334gat));
  OAI21_X1  g521(.A(G78gat), .B1(new_n707_), .B2(new_n559_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT50), .ZN(new_n724_));
  INV_X1    g523(.A(G78gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n710_), .A2(new_n725_), .A3(new_n650_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1335gat));
  INV_X1    g526(.A(KEYINPUT116), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n709_), .A2(new_n348_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n670_), .A2(KEYINPUT115), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT115), .B1(new_n670_), .B2(new_n729_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n575_), .A2(new_n658_), .A3(new_n317_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n667_), .A2(new_n668_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n575_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n737_), .B2(KEYINPUT43), .ZN(new_n738_));
  INV_X1    g537(.A(new_n729_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n734_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(KEYINPUT116), .A3(new_n730_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n733_), .A2(new_n419_), .A3(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G85gat), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n677_), .A2(new_n729_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n569_), .A2(G85gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(G1336gat));
  NAND3_X1  g545(.A1(new_n733_), .A2(new_n639_), .A3(new_n741_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G92gat), .ZN(new_n748_));
  OR3_X1    g547(.A1(new_n744_), .A2(G92gat), .A3(new_n568_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT117), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT117), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n752_), .A3(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1337gat));
  INV_X1    g553(.A(new_n744_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n646_), .C1(new_n248_), .C2(new_n247_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n731_), .A2(new_n529_), .A3(new_n732_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n233_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g558(.A(new_n658_), .B1(new_n736_), .B2(new_n575_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n650_), .B(new_n729_), .C1(new_n760_), .C2(new_n735_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT118), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n670_), .A2(KEYINPUT118), .A3(new_n650_), .A4(new_n729_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(G106gat), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT119), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT119), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n763_), .A2(new_n764_), .A3(new_n767_), .A4(G106gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(KEYINPUT52), .A3(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n755_), .A2(new_n246_), .A3(new_n650_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n765_), .A2(KEYINPUT119), .A3(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT53), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n769_), .A2(new_n775_), .A3(new_n770_), .A4(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1339gat));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n610_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT120), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n610_), .A2(new_n779_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n603_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(G230gat), .A3(G233gat), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n610_), .A2(new_n785_), .A3(new_n779_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n781_), .A2(new_n782_), .A3(new_n784_), .A4(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n619_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT121), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n601_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n621_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n586_), .A2(new_n582_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n593_), .B1(new_n581_), .B2(new_n587_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n600_), .A2(new_n599_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n791_), .A2(new_n793_), .B1(new_n622_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n778_), .B1(new_n797_), .B2(new_n632_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n622_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n601_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n788_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n790_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n803_), .B2(new_n792_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(KEYINPUT57), .A3(new_n313_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(KEYINPUT122), .A2(KEYINPUT56), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n787_), .A2(new_n619_), .A3(new_n806_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(new_n621_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(KEYINPUT122), .A2(KEYINPUT56), .ZN(new_n809_));
  INV_X1    g608(.A(new_n806_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n788_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n796_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n808_), .A2(KEYINPUT58), .A3(new_n796_), .A4(new_n811_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n317_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n798_), .A2(new_n805_), .A3(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n800_), .A2(new_n626_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n350_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT54), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n350_), .A2(new_n821_), .A3(new_n818_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n817_), .A2(new_n349_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n573_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n639_), .A2(new_n569_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828_), .B2(new_n800_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(KEYINPUT59), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n601_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n829_), .B1(new_n833_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g633(.A(G120gat), .ZN(new_n835_));
  INV_X1    g634(.A(new_n626_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(KEYINPUT60), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n828_), .B(new_n837_), .C1(KEYINPUT60), .C2(new_n835_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n835_), .ZN(G1341gat));
  AOI21_X1  g639(.A(G127gat), .B1(new_n828_), .B2(new_n348_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n349_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g642(.A(G134gat), .B1(new_n828_), .B2(new_n632_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n830_), .A2(new_n832_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n317_), .A2(G134gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT123), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n844_), .B1(new_n845_), .B2(new_n847_), .ZN(G1343gat));
  NOR3_X1   g647(.A1(new_n823_), .A2(new_n646_), .A3(new_n559_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n849_), .A2(new_n826_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n800_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n626_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT124), .B(G148gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1345gat));
  NAND2_X1  g654(.A1(new_n850_), .A2(new_n348_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT125), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n856_), .B(new_n858_), .ZN(G1346gat));
  AOI21_X1  g658(.A(G162gat), .B1(new_n850_), .B2(new_n632_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n299_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n850_), .B2(new_n861_), .ZN(G1347gat));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n568_), .A2(new_n419_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR4_X1   g664(.A1(new_n823_), .A2(new_n601_), .A3(new_n824_), .A4(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT126), .B(new_n863_), .C1(new_n866_), .C2(new_n453_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n823_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n868_), .A2(new_n800_), .A3(new_n573_), .A4(new_n864_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n863_), .A2(KEYINPUT126), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n863_), .A2(KEYINPUT126), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n869_), .A2(G169gat), .A3(new_n870_), .A4(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n866_), .A2(new_n439_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n867_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT127), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n867_), .A2(new_n872_), .A3(KEYINPUT127), .A4(new_n873_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1348gat));
  NAND2_X1  g677(.A1(new_n825_), .A2(new_n864_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n836_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n440_), .ZN(G1349gat));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n349_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n450_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n882_), .B2(new_n442_), .ZN(G1350gat));
  INV_X1    g683(.A(new_n317_), .ZN(new_n885_));
  OAI21_X1  g684(.A(G190gat), .B1(new_n879_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n632_), .A2(new_n451_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n879_), .B2(new_n887_), .ZN(G1351gat));
  AND2_X1   g687(.A1(new_n849_), .A2(new_n864_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n800_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n626_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g692(.A(KEYINPUT63), .B(G211gat), .Z(new_n894_));
  AND3_X1   g693(.A1(new_n889_), .A2(new_n348_), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n889_), .A2(new_n348_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1354gat));
  AOI21_X1  g697(.A(G218gat), .B1(new_n889_), .B2(new_n632_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n889_), .A2(new_n317_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(G218gat), .B2(new_n900_), .ZN(G1355gat));
endmodule


