//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT8), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(G99gat), .ZN(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n205_), .A2(new_n207_), .B1(new_n210_), .B2(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n215_));
  NAND2_X1  g014(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n211_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G85gat), .B(G92gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n203_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G29gat), .B(G36gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(G43gat), .B(G50gat), .Z(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n219_), .B1(new_n211_), .B2(new_n217_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT8), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT10), .B(G99gat), .Z(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n209_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G85gat), .B(G92gat), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT9), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n205_), .A2(new_n207_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT9), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G85gat), .A3(G92gat), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .A4(new_n236_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n220_), .A2(new_n227_), .A3(new_n229_), .A4(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT34), .Z(new_n240_));
  INV_X1    g039(.A(KEYINPUT35), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT70), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n224_), .A2(KEYINPUT15), .A3(new_n226_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT15), .B1(new_n224_), .B2(new_n226_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n237_), .B1(new_n228_), .B2(KEYINPUT8), .ZN(new_n248_));
  INV_X1    g047(.A(new_n229_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n240_), .A2(new_n241_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n244_), .B(new_n250_), .C1(KEYINPUT69), .C2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n250_), .A2(new_n238_), .A3(new_n243_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n238_), .A2(KEYINPUT69), .A3(new_n243_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(new_n251_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G190gat), .B(G218gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(G134gat), .B(G162gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT36), .Z(new_n263_));
  NAND2_X1  g062(.A1(new_n257_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n262_), .A2(KEYINPUT36), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n253_), .A2(new_n256_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n202_), .B1(new_n267_), .B2(KEYINPUT37), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT37), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n264_), .A2(KEYINPUT74), .A3(new_n269_), .A4(new_n266_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n266_), .B1(new_n264_), .B2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT73), .B1(new_n257_), .B2(new_n263_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT37), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n271_), .A2(KEYINPUT75), .A3(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT76), .B(G8gat), .Z(new_n281_));
  INV_X1    g080(.A(G1gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT14), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G15gat), .B(G22gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G1gat), .B(G8gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n283_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G57gat), .B(G64gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(KEYINPUT11), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n292_), .A2(KEYINPUT11), .ZN(new_n295_));
  XOR2_X1   g094(.A(G71gat), .B(G78gat), .Z(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n291_), .A3(KEYINPUT11), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(KEYINPUT11), .B2(new_n292_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n297_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n299_), .B1(new_n300_), .B2(new_n293_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n290_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G231gat), .A2(G233gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n307_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT17), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G127gat), .B(G155gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT16), .ZN(new_n313_));
  XOR2_X1   g112(.A(G183gat), .B(G211gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n310_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n311_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n308_), .A2(new_n317_), .A3(new_n309_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n280_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT27), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT23), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT23), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(G183gat), .A3(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(G183gat), .ZN(new_n327_));
  INV_X1    g126(.A(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G169gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT24), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n335_), .A2(G169gat), .A3(G176gat), .ZN(new_n336_));
  INV_X1    g135(.A(G169gat), .ZN(new_n337_));
  INV_X1    g136(.A(G176gat), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT82), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n334_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n334_), .B1(G169gat), .B2(G176gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n338_), .A3(KEYINPUT82), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n335_), .B1(G169gat), .B2(G176gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n327_), .A2(KEYINPUT25), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT25), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G183gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n328_), .A2(KEYINPUT26), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT26), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G190gat), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n340_), .A2(new_n344_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n323_), .A2(new_n325_), .A3(KEYINPUT83), .ZN(new_n353_));
  OR3_X1    g152(.A1(new_n322_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n333_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G218gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G211gat), .ZN(new_n358_));
  INV_X1    g157(.A(G211gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G218gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT88), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(KEYINPUT21), .A3(new_n365_), .ZN(new_n366_));
  OR2_X1    g165(.A1(G197gat), .A2(G204gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G197gat), .A2(G204gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(KEYINPUT21), .A3(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n361_), .A3(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n358_), .B(new_n360_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT89), .B(KEYINPUT21), .Z(new_n374_));
  AOI22_X1  g173(.A1(new_n366_), .A2(new_n371_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT90), .B1(new_n356_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n353_), .A2(new_n354_), .A3(new_n329_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n332_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n340_), .A2(new_n326_), .A3(new_n344_), .A4(new_n351_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n377_), .B1(new_n381_), .B2(new_n375_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n371_), .A2(new_n366_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n373_), .A2(new_n374_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n353_), .A2(new_n354_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n386_), .A2(new_n344_), .A3(new_n340_), .A4(new_n351_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT90), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n385_), .A2(new_n387_), .A3(new_n388_), .A4(new_n333_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n376_), .A2(new_n382_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT19), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G8gat), .B(G36gat), .Z(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT18), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G64gat), .B(G92gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n356_), .A2(new_n375_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n385_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT20), .A4(new_n392_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n394_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n399_), .B1(new_n394_), .B2(new_n402_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n321_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n404_), .ZN(new_n406_));
  AND4_X1   g205(.A1(KEYINPUT20), .A2(new_n400_), .A3(new_n401_), .A4(new_n393_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n385_), .A2(new_n387_), .A3(new_n333_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n393_), .B1(new_n382_), .B2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT94), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT20), .A4(new_n393_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT94), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n398_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT95), .ZN(new_n415_));
  OAI211_X1 g214(.A(KEYINPUT27), .B(new_n406_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n416_));
  AOI211_X1 g215(.A(KEYINPUT95), .B(new_n398_), .C1(new_n410_), .C2(new_n413_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n405_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G1gat), .B(G29gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(G85gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT0), .B(G57gat), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(new_n421_), .Z(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(G155gat), .A2(G162gat), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n426_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n430_));
  INV_X1    g229(.A(G155gat), .ZN(new_n431_));
  INV_X1    g230(.A(G162gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI221_X1 g234(.A(new_n427_), .B1(new_n429_), .B2(new_n430_), .C1(KEYINPUT1), .C2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT86), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G155gat), .A2(G162gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n426_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n433_), .A2(KEYINPUT86), .A3(new_n434_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G141gat), .ZN(new_n442_));
  INV_X1    g241(.A(G148gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT3), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT3), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(G141gat), .B2(G148gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  AND3_X1   g246(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n447_), .A2(new_n450_), .A3(KEYINPUT85), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n441_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT85), .B1(new_n447_), .B2(new_n450_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n436_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G127gat), .B(G134gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G113gat), .B(G120gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n425_), .B1(new_n459_), .B2(KEYINPUT4), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n457_), .B(new_n436_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(KEYINPUT4), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT91), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT91), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n459_), .A2(new_n464_), .A3(KEYINPUT4), .A4(new_n461_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n460_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n459_), .A2(new_n461_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(new_n425_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n423_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n460_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n461_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n444_), .A2(new_n446_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n449_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n472_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(new_n451_), .A3(new_n441_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n457_), .B1(new_n478_), .B2(new_n436_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n471_), .A2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n464_), .B1(new_n480_), .B2(KEYINPUT4), .ZN(new_n481_));
  INV_X1    g280(.A(new_n465_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n470_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n422_), .B1(new_n467_), .B2(new_n425_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n469_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G71gat), .B(G99gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(G43gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n381_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(new_n458_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G227gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(G15gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT30), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT31), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n491_), .B(new_n496_), .Z(new_n497_));
  NAND2_X1  g296(.A1(new_n487_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G233gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n500_), .A2(G228gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(G228gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n499_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(G78gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(new_n209_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G22gat), .B(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OR3_X1    g307(.A1(new_n454_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT28), .B1(new_n454_), .B2(KEYINPUT29), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n454_), .A2(KEYINPUT29), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(new_n385_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n509_), .B(new_n510_), .C1(new_n385_), .C2(new_n512_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n508_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n507_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n418_), .A2(new_n498_), .A3(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n414_), .A2(new_n415_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n414_), .A2(new_n415_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n521_), .A2(KEYINPUT27), .A3(new_n406_), .A4(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n523_), .A2(new_n487_), .A3(new_n519_), .A4(new_n405_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT32), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n399_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n381_), .A2(new_n375_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n408_), .A2(new_n527_), .A3(KEYINPUT20), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n392_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n412_), .B1(new_n529_), .B2(new_n411_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n413_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n526_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n394_), .A2(new_n402_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n525_), .B2(new_n399_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(new_n486_), .B2(new_n469_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT33), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n486_), .B2(KEYINPUT92), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n403_), .A2(new_n404_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(KEYINPUT33), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n541_), .B1(new_n466_), .B2(new_n484_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n463_), .A2(new_n465_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT4), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n425_), .B1(new_n479_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT93), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n545_), .A2(new_n550_), .A3(new_n547_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n422_), .B1(new_n480_), .B2(new_n425_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n536_), .B1(new_n544_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n524_), .B1(new_n554_), .B2(new_n519_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n497_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n520_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT79), .ZN(new_n558_));
  INV_X1    g357(.A(new_n289_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n286_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n559_), .A2(new_n227_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n227_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n558_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n227_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n288_), .A2(new_n562_), .A3(new_n289_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(KEYINPUT79), .A3(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n247_), .A2(new_n289_), .A3(new_n288_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT80), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT80), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n571_), .A2(new_n574_), .A3(new_n565_), .A4(new_n567_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n570_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G113gat), .B(G141gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT81), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G169gat), .B(G197gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n570_), .A2(new_n573_), .A3(new_n575_), .A4(new_n580_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT64), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n248_), .A2(new_n249_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(new_n302_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n298_), .A2(new_n301_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n589_), .A2(new_n249_), .A3(new_n248_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n586_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT12), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n587_), .B2(new_n302_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n586_), .B1(new_n587_), .B2(new_n302_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n589_), .B(KEYINPUT12), .C1(new_n249_), .C2(new_n248_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G120gat), .B(G148gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT5), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n598_), .B(new_n599_), .Z(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n591_), .A2(new_n596_), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n591_), .B2(new_n596_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT13), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n591_), .A2(new_n596_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n600_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n591_), .A2(new_n596_), .A3(new_n601_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT13), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n605_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT68), .ZN(new_n613_));
  NOR4_X1   g412(.A1(new_n320_), .A2(new_n557_), .A3(new_n584_), .A4(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n469_), .A2(new_n486_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n282_), .A3(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n267_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n557_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n612_), .A2(new_n584_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n319_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT97), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT98), .ZN(new_n625_));
  OAI21_X1  g424(.A(G1gat), .B1(new_n625_), .B2(new_n487_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n618_), .A2(new_n626_), .ZN(G1324gat));
  NAND3_X1  g426(.A1(new_n614_), .A2(new_n418_), .A3(new_n281_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT99), .ZN(new_n629_));
  INV_X1    g428(.A(new_n418_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G8gat), .B1(new_n624_), .B2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT39), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1325gat));
  OAI21_X1  g434(.A(G15gat), .B1(new_n625_), .B2(new_n556_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT41), .Z(new_n637_));
  NAND3_X1  g436(.A1(new_n614_), .A2(new_n493_), .A3(new_n497_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1326gat));
  INV_X1    g438(.A(new_n519_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G22gat), .B1(new_n625_), .B2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT42), .ZN(new_n642_));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n614_), .A2(new_n643_), .A3(new_n519_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1327gat));
  NOR2_X1   g444(.A1(new_n557_), .A2(new_n584_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n319_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n619_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n612_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G29gat), .B1(new_n651_), .B2(new_n615_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n647_), .A2(new_n621_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT43), .B1(new_n557_), .B2(new_n280_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n484_), .B1(new_n545_), .B2(new_n470_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT33), .B1(new_n656_), .B2(new_n540_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n553_), .A2(new_n657_), .A3(new_n539_), .A4(new_n542_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n615_), .A2(new_n534_), .A3(new_n532_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n519_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n487_), .A2(new_n519_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n418_), .A2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n556_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n520_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n271_), .A2(KEYINPUT75), .A3(new_n275_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT75), .B1(new_n271_), .B2(new_n275_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n654_), .B1(new_n655_), .B2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n653_), .B1(new_n671_), .B2(KEYINPUT44), .ZN(new_n672_));
  INV_X1    g471(.A(new_n654_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n665_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n669_), .B1(new_n665_), .B2(new_n668_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(KEYINPUT100), .A3(new_n677_), .ZN(new_n678_));
  AOI22_X1  g477(.A1(new_n672_), .A2(new_n678_), .B1(KEYINPUT44), .B2(new_n671_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n615_), .A2(G29gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n652_), .B1(new_n679_), .B2(new_n680_), .ZN(G1328gat));
  INV_X1    g480(.A(G36gat), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n646_), .A2(new_n682_), .A3(new_n418_), .A4(new_n649_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT45), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT44), .B(new_n673_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n418_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n672_), .B2(new_n678_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(new_n687_), .B2(new_n682_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(KEYINPUT101), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n688_), .B2(KEYINPUT101), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1329gat));
  NAND3_X1  g491(.A1(new_n679_), .A2(G43gat), .A3(new_n497_), .ZN(new_n693_));
  INV_X1    g492(.A(G43gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(new_n650_), .B2(new_n556_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n693_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1330gat));
  OR3_X1    g498(.A1(new_n650_), .A2(G50gat), .A3(new_n640_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n679_), .A2(new_n519_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(G50gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n701_), .B2(G50gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(G1331gat));
  INV_X1    g504(.A(new_n613_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n319_), .A2(new_n584_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT105), .B(G57gat), .Z(new_n709_));
  NAND4_X1  g508(.A1(new_n620_), .A2(new_n615_), .A3(new_n708_), .A4(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT106), .ZN(new_n711_));
  INV_X1    g510(.A(new_n612_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n320_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n584_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n557_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n615_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n711_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT107), .ZN(G1332gat));
  NAND2_X1  g519(.A1(new_n620_), .A2(new_n708_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G64gat), .B1(new_n721_), .B2(new_n630_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT48), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n630_), .A2(G64gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n716_), .B2(new_n724_), .ZN(G1333gat));
  OR3_X1    g524(.A1(new_n716_), .A2(G71gat), .A3(new_n556_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G71gat), .B1(new_n721_), .B2(new_n556_), .ZN(new_n727_));
  XOR2_X1   g526(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n727_), .A2(new_n729_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n726_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT109), .Z(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n721_), .B2(new_n640_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n640_), .A2(G78gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n716_), .B2(new_n736_), .ZN(G1335gat));
  NAND2_X1  g536(.A1(new_n655_), .A2(new_n670_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n319_), .A2(new_n714_), .A3(new_n712_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n487_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n706_), .A2(new_n648_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n715_), .A2(new_n742_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n487_), .A2(G85gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n741_), .B1(new_n743_), .B2(new_n744_), .ZN(G1336gat));
  OAI21_X1  g544(.A(G92gat), .B1(new_n740_), .B2(new_n630_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n630_), .A2(G92gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n743_), .B2(new_n747_), .ZN(G1337gat));
  NAND3_X1  g547(.A1(new_n738_), .A2(new_n497_), .A3(new_n739_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G99gat), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT110), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT110), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n497_), .A2(new_n230_), .ZN(new_n753_));
  OAI22_X1  g552(.A1(new_n751_), .A2(new_n752_), .B1(new_n743_), .B2(new_n753_), .ZN(new_n754_));
  AND2_X1   g553(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(G1338gat));
  XNOR2_X1  g555(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n738_), .A2(new_n519_), .A3(new_n739_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G106gat), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n715_), .A2(new_n209_), .A3(new_n519_), .A4(new_n742_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n757_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n763_), .B(new_n757_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  NOR4_X1   g566(.A1(new_n418_), .A2(new_n556_), .A3(new_n487_), .A4(new_n519_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n564_), .A2(new_n565_), .A3(new_n569_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n571_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n581_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n583_), .A2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(new_n602_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n596_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n587_), .A2(new_n302_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n593_), .A2(new_n777_), .A3(new_n595_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n586_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n593_), .A2(new_n594_), .A3(KEYINPUT55), .A4(new_n595_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n776_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n600_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n600_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n774_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT58), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(KEYINPUT116), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n786_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n278_), .A2(new_n279_), .A3(new_n787_), .A4(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT115), .B1(new_n604_), .B2(new_n773_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n773_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n609_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n602_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(KEYINPUT114), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n798_), .B(new_n795_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n619_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n789_), .B1(new_n800_), .B2(KEYINPUT57), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n796_), .A2(KEYINPUT114), .ZN(new_n802_));
  INV_X1    g601(.A(new_n794_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n799_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n267_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n647_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n707_), .A2(new_n612_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n280_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n810_), .B(new_n280_), .C1(KEYINPUT113), .C2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n769_), .B1(new_n809_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(G113gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n714_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT117), .B(new_n647_), .C1(new_n801_), .C2(new_n808_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n806_), .A2(new_n807_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n800_), .A2(KEYINPUT57), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n789_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT117), .B1(new_n824_), .B2(new_n647_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n816_), .B1(new_n821_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n768_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n817_), .A2(new_n827_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n714_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n819_), .B1(new_n831_), .B2(new_n818_), .ZN(G1340gat));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n828_), .A2(new_n833_), .A3(new_n613_), .A4(new_n829_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n816_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n809_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n837_), .B2(new_n820_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n768_), .A2(new_n827_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n613_), .B1(new_n817_), .B2(new_n827_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT118), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n834_), .A2(new_n842_), .A3(G120gat), .ZN(new_n843_));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n712_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n817_), .B(new_n845_), .C1(KEYINPUT60), .C2(new_n844_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(G1341gat));
  INV_X1    g646(.A(G127gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n817_), .A2(new_n848_), .A3(new_n319_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n828_), .A2(new_n319_), .A3(new_n829_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n849_), .B1(new_n851_), .B2(new_n848_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n817_), .A2(new_n853_), .A3(new_n619_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n828_), .A2(new_n668_), .A3(new_n829_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n856_), .B2(new_n853_), .ZN(G1343gat));
  NAND2_X1  g656(.A1(new_n809_), .A2(new_n816_), .ZN(new_n858_));
  NOR4_X1   g657(.A1(new_n418_), .A2(new_n640_), .A3(new_n487_), .A4(new_n497_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT119), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n584_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n442_), .ZN(G1344gat));
  NOR2_X1   g662(.A1(new_n861_), .A2(new_n706_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT120), .B(G148gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1345gat));
  NOR2_X1   g665(.A1(new_n861_), .A2(new_n647_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT61), .B(G155gat), .Z(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n861_), .B2(new_n280_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n619_), .A2(new_n432_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n861_), .B2(new_n871_), .ZN(G1347gat));
  INV_X1    g671(.A(KEYINPUT22), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n630_), .A2(new_n498_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n519_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n826_), .A2(new_n873_), .A3(new_n714_), .A4(new_n876_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n877_), .A2(KEYINPUT62), .A3(new_n337_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(KEYINPUT62), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n826_), .A2(new_n880_), .A3(new_n714_), .A4(new_n876_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(G169gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n878_), .B1(new_n879_), .B2(new_n882_), .ZN(G1348gat));
  NAND2_X1  g682(.A1(new_n826_), .A2(new_n876_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n338_), .B1(new_n884_), .B2(new_n712_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(KEYINPUT121), .B(new_n338_), .C1(new_n884_), .C2(new_n712_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n519_), .B1(new_n809_), .B2(new_n816_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n706_), .A2(new_n338_), .A3(new_n875_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n887_), .A2(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(G1349gat));
  NOR2_X1   g690(.A1(new_n875_), .A2(new_n647_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G183gat), .B1(new_n889_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n884_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n647_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1350gat));
  NAND4_X1  g695(.A1(new_n894_), .A2(new_n619_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n826_), .A2(new_n668_), .A3(new_n876_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(G190gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(G190gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n897_), .B1(new_n900_), .B2(new_n901_), .ZN(G1351gat));
  NOR3_X1   g701(.A1(new_n630_), .A2(new_n661_), .A3(new_n497_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n858_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n714_), .ZN(new_n905_));
  INV_X1    g704(.A(G197gat), .ZN(new_n906_));
  OR3_X1    g705(.A1(new_n905_), .A2(KEYINPUT123), .A3(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT123), .B1(new_n905_), .B2(new_n906_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n906_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(G1352gat));
  INV_X1    g709(.A(new_n904_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n706_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT124), .B(G204gat), .Z(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n912_), .B2(new_n915_), .ZN(G1353gat));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n319_), .B1(new_n917_), .B2(new_n359_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT125), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n904_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n917_), .A2(new_n359_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1354gat));
  XOR2_X1   g721(.A(KEYINPUT127), .B(G218gat), .Z(new_n923_));
  NOR3_X1   g722(.A1(new_n911_), .A2(new_n280_), .A3(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n904_), .A2(new_n619_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT126), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n926_), .B2(new_n923_), .ZN(G1355gat));
endmodule


