//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  INV_X1    g006(.A(G1gat), .ZN(new_n208_));
  INV_X1    g007(.A(G8gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n212_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G29gat), .B(G36gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G43gat), .B(G50gat), .Z(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n216_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT15), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT15), .B1(new_n219_), .B2(new_n221_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n215_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT78), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n219_), .A2(new_n221_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(new_n214_), .A3(new_n213_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT78), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n215_), .B(new_n230_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n225_), .A2(new_n226_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n215_), .A2(new_n227_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n233_), .A3(KEYINPUT76), .ZN(new_n234_));
  INV_X1    g033(.A(new_n226_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n215_), .A2(new_n236_), .A3(new_n227_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n206_), .B1(new_n232_), .B2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n206_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n205_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(KEYINPUT79), .B(new_n204_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G113gat), .B(G120gat), .Z(new_n247_));
  NOR2_X1   g046(.A1(G127gat), .A2(G134gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT82), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G127gat), .A2(G134gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT82), .B1(new_n253_), .B2(new_n248_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n247_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT83), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n252_), .A2(new_n254_), .A3(new_n247_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT84), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n252_), .A2(new_n254_), .A3(new_n247_), .A4(KEYINPUT84), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT83), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n255_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n257_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G227gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G15gat), .B(G43gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT31), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n271_), .B(new_n272_), .Z(new_n273_));
  INV_X1    g072(.A(KEYINPUT80), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT25), .B(G183gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT23), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(G183gat), .A3(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT24), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n279_), .A2(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(KEYINPUT24), .A3(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n277_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n290_));
  OR2_X1    g089(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(G176gat), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n286_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n290_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n274_), .B1(new_n288_), .B2(new_n295_), .ZN(new_n296_));
  OR3_X1    g095(.A1(new_n290_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n277_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(KEYINPUT80), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n273_), .B(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n269_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(KEYINPUT86), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n303_), .A2(G155gat), .A3(G162gat), .ZN(new_n304_));
  INV_X1    g103(.A(G155gat), .ZN(new_n305_));
  INV_X1    g104(.A(G162gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT86), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n305_), .A2(new_n306_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n309_));
  OAI22_X1  g108(.A1(new_n304_), .A2(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT87), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n309_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT87), .ZN(new_n313_));
  OAI221_X1 g112(.A(new_n313_), .B1(new_n308_), .B2(new_n309_), .C1(new_n307_), .C2(new_n304_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT85), .Z(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(KEYINPUT88), .A2(KEYINPUT3), .ZN(new_n323_));
  OAI22_X1  g122(.A1(new_n322_), .A2(new_n323_), .B1(G141gat), .B2(G148gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n316_), .B(KEYINPUT2), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n317_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT89), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n304_), .A2(new_n307_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n324_), .A2(new_n325_), .A3(new_n330_), .A4(new_n326_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n308_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n319_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT29), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G228gat), .A2(G233gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(KEYINPUT29), .ZN(new_n337_));
  OR2_X1    g136(.A1(G211gat), .A2(G218gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G211gat), .A2(G218gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT90), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n338_), .A2(KEYINPUT90), .A3(new_n339_), .ZN(new_n343_));
  INV_X1    g142(.A(G204gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G197gat), .ZN(new_n345_));
  INV_X1    g144(.A(G197gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G204gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n342_), .A2(new_n343_), .B1(new_n348_), .B2(KEYINPUT21), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(KEYINPUT21), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n343_), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT90), .B1(new_n338_), .B2(new_n339_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n349_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n336_), .B1(new_n337_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(new_n319_), .B2(new_n333_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n348_), .A2(KEYINPUT21), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n351_), .A2(new_n352_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n342_), .B(new_n343_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n350_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n336_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n361_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n335_), .B1(new_n359_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n337_), .A2(new_n358_), .A3(new_n336_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n335_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n367_), .B1(new_n361_), .B2(new_n366_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G78gat), .B(G106gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT91), .B(G50gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT28), .B(G22gat), .Z(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n369_), .A2(new_n373_), .A3(new_n379_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n257_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n334_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n256_), .A2(new_n258_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n319_), .A2(new_n333_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n265_), .B1(new_n333_), .B2(new_n319_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(KEYINPUT4), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n385_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n388_), .A2(new_n384_), .A3(new_n390_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT96), .ZN(new_n397_));
  XOR2_X1   g196(.A(G57gat), .B(G85gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n394_), .A2(new_n395_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT97), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT33), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n384_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n388_), .A2(new_n385_), .A3(new_n390_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n401_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n403_), .A2(new_n404_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n297_), .A2(new_n298_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT93), .B1(new_n358_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n358_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT93), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n366_), .A2(new_n415_), .A3(new_n297_), .A4(new_n298_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n413_), .A2(new_n414_), .A3(new_n416_), .A4(KEYINPUT20), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G226gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n300_), .A2(new_n366_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n420_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n358_), .A2(new_n412_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n422_), .A2(KEYINPUT20), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n426_));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G8gat), .B(G36gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n421_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(new_n421_), .B2(new_n425_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n406_), .A2(new_n409_), .A3(new_n411_), .A4(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n390_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT4), .B1(new_n392_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n388_), .A2(new_n386_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n384_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n395_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n401_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n403_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n421_), .A2(new_n425_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT32), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n444_), .B1(new_n445_), .B2(new_n431_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n414_), .B(KEYINPUT20), .C1(new_n412_), .C2(new_n358_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n423_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n422_), .A2(KEYINPUT20), .A3(new_n420_), .A4(new_n424_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(KEYINPUT32), .A3(new_n430_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(new_n446_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n383_), .B1(new_n436_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT98), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n369_), .A2(new_n373_), .A3(new_n379_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n379_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n442_), .B(new_n403_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n430_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n444_), .A2(new_n430_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT27), .A3(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n435_), .B2(KEYINPUT27), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n454_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT27), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n434_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT27), .B1(new_n460_), .B2(new_n432_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n442_), .A2(new_n403_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(KEYINPUT98), .A4(new_n383_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n463_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n302_), .B1(new_n453_), .B2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n302_), .A2(new_n443_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n383_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n467_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n246_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G232gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT34), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT68), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT6), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT7), .ZN(new_n484_));
  INV_X1    g283(.A(G99gat), .ZN(new_n485_));
  INV_X1    g284(.A(G106gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n478_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n481_), .A2(new_n483_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G85gat), .A2(G92gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G85gat), .A2(G92gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT8), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT69), .ZN(new_n497_));
  XOR2_X1   g296(.A(KEYINPUT66), .B(KEYINPUT8), .Z(new_n498_));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n482_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n487_), .A2(new_n478_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n494_), .B(new_n498_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT67), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT69), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n495_), .A2(new_n505_), .A3(KEYINPUT8), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n497_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT9), .ZN(new_n508_));
  INV_X1    g307(.A(G85gat), .ZN(new_n509_));
  INV_X1    g308(.A(G92gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n508_), .B1(new_n511_), .B2(new_n491_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n491_), .A2(new_n508_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT65), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n516_), .B(new_n513_), .C1(new_n494_), .C2(new_n508_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT10), .B(G99gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT64), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n486_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT64), .B1(new_n519_), .B2(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n518_), .A2(new_n524_), .A3(new_n483_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n507_), .A2(new_n525_), .A3(new_n228_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n222_), .A2(new_n223_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n500_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(KEYINPUT70), .A3(new_n524_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n527_), .B1(new_n507_), .B2(new_n532_), .ZN(new_n533_));
  OAI211_X1 g332(.A(KEYINPUT35), .B(new_n477_), .C1(new_n526_), .C2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n502_), .B(KEYINPUT67), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n505_), .B1(new_n495_), .B2(KEYINPUT8), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT8), .ZN(new_n537_));
  AOI211_X1 g336(.A(KEYINPUT69), .B(new_n537_), .C1(new_n490_), .C2(new_n494_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n535_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n530_), .A2(KEYINPUT70), .A3(new_n524_), .ZN(new_n540_));
  AOI21_X1  g339(.A(KEYINPUT70), .B1(new_n530_), .B2(new_n524_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI22_X1  g341(.A1(new_n539_), .A2(new_n542_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n477_), .A2(KEYINPUT35), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n477_), .A2(KEYINPUT35), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n507_), .A2(new_n525_), .A3(new_n228_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n534_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT36), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n534_), .A2(new_n547_), .A3(KEYINPUT73), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n550_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n534_), .A2(new_n547_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G71gat), .B(G78gat), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n566_), .A3(KEYINPUT11), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(new_n215_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(G211gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(KEYINPUT16), .B(G183gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n572_), .A2(new_n573_), .A3(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(KEYINPUT17), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n572_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n507_), .A2(new_n525_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n569_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT12), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(G230gat), .ZN(new_n587_));
  INV_X1    g386(.A(G233gat), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n507_), .A2(new_n525_), .A3(new_n569_), .ZN(new_n591_));
  OAI211_X1 g390(.A(KEYINPUT12), .B(new_n583_), .C1(new_n539_), .C2(new_n542_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n586_), .A2(new_n590_), .A3(new_n591_), .A4(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n584_), .A2(new_n591_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n589_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G204gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT5), .B(G176gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n593_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT13), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT71), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(KEYINPUT71), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n601_), .A2(new_n602_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n593_), .A2(new_n595_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n599_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n593_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n604_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n581_), .B1(new_n606_), .B2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n475_), .A2(new_n562_), .A3(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n468_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n556_), .A2(new_n615_), .A3(new_n561_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT74), .ZN(new_n617_));
  INV_X1    g416(.A(new_n554_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n534_), .B2(new_n547_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT37), .B1(new_n560_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT72), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT72), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n622_), .B(KEYINPUT37), .C1(new_n560_), .C2(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT74), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n556_), .A2(new_n625_), .A3(new_n615_), .A4(new_n561_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n617_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n581_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT75), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n606_), .A2(new_n611_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n475_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n208_), .A3(new_n443_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT99), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(KEYINPUT99), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n614_), .B1(new_n638_), .B2(new_n639_), .ZN(G1324gat));
  XNOR2_X1  g439(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n613_), .A2(new_n467_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(G8gat), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(KEYINPUT39), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(KEYINPUT39), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n633_), .A2(new_n209_), .A3(new_n462_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n641_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n647_), .B(new_n641_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n648_), .A2(new_n650_), .ZN(G1325gat));
  OAI21_X1  g450(.A(G15gat), .B1(new_n613_), .B2(new_n302_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT41), .Z(new_n653_));
  INV_X1    g452(.A(new_n633_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n302_), .A2(G15gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n653_), .B1(new_n654_), .B2(new_n655_), .ZN(G1326gat));
  OAI21_X1  g455(.A(G22gat), .B1(new_n613_), .B2(new_n473_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT42), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n473_), .A2(G22gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n654_), .B2(new_n659_), .ZN(G1327gat));
  AOI211_X1 g459(.A(new_n246_), .B(new_n628_), .C1(new_n606_), .C2(new_n611_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n627_), .A2(KEYINPUT102), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n617_), .A2(new_n624_), .A3(new_n664_), .A4(new_n626_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n471_), .A2(new_n474_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n662_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  AOI211_X1 g467(.A(KEYINPUT43), .B(new_n627_), .C1(new_n471_), .C2(new_n474_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n661_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n673_), .B(new_n661_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(new_n443_), .A3(new_n674_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(KEYINPUT104), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(KEYINPUT104), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(G29gat), .A3(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n562_), .A2(new_n628_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n632_), .A2(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n468_), .A2(G29gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(G1328gat));
  NOR3_X1   g481(.A1(new_n680_), .A2(G36gat), .A3(new_n467_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n672_), .A2(new_n462_), .A3(new_n674_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n686_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT105), .B1(new_n686_), .B2(G36gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n685_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n685_), .B(KEYINPUT46), .C1(new_n687_), .C2(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  NOR3_X1   g492(.A1(new_n680_), .A2(G43gat), .A3(new_n302_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n302_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n672_), .A2(new_n695_), .A3(new_n674_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n696_), .B2(G43gat), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g497(.A1(new_n672_), .A2(new_n383_), .A3(new_n674_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(new_n700_), .A3(G50gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(G50gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n473_), .A2(G50gat), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT107), .Z(new_n704_));
  OAI22_X1  g503(.A1(new_n701_), .A2(new_n702_), .B1(new_n680_), .B2(new_n704_), .ZN(G1331gat));
  AOI21_X1  g504(.A(new_n245_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n631_), .A2(new_n581_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n562_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(G57gat), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n468_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT109), .Z(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n706_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n706_), .A2(new_n712_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n631_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n443_), .A3(new_n630_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n711_), .B1(new_n716_), .B2(new_n709_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n708_), .B2(new_n467_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT48), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(new_n630_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n467_), .A2(G64gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n720_), .B2(new_n721_), .ZN(G1333gat));
  OAI21_X1  g521(.A(G71gat), .B1(new_n708_), .B2(new_n302_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT49), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n302_), .A2(G71gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n720_), .B2(new_n725_), .ZN(G1334gat));
  OAI21_X1  g525(.A(G78gat), .B1(new_n708_), .B2(new_n473_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT50), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n473_), .A2(G78gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n720_), .B2(new_n729_), .ZN(G1335gat));
  OR2_X1    g529(.A1(new_n668_), .A2(new_n669_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n631_), .A2(new_n628_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n246_), .A3(new_n732_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n733_), .A2(new_n509_), .A3(new_n468_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n679_), .ZN(new_n735_));
  NOR4_X1   g534(.A1(new_n713_), .A2(new_n714_), .A3(new_n631_), .A4(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n443_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n734_), .A2(new_n737_), .ZN(G1336gat));
  NOR3_X1   g537(.A1(new_n733_), .A2(new_n510_), .A3(new_n467_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G92gat), .B1(new_n736_), .B2(new_n462_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n733_), .B2(new_n302_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n736_), .A2(new_n520_), .A3(new_n695_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g544(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n736_), .A2(new_n486_), .A3(new_n383_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n736_), .A2(KEYINPUT110), .A3(new_n486_), .A4(new_n383_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n731_), .A2(new_n246_), .A3(new_n383_), .A4(new_n732_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G106gat), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n747_), .B1(new_n752_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n750_), .A2(new_n751_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n760_), .A2(new_n746_), .A3(new_n757_), .A4(new_n756_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  AND2_X1   g561(.A1(new_n234_), .A2(new_n237_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n205_), .B1(new_n763_), .B2(new_n226_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n764_), .B(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n225_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n768_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n235_), .A3(new_n770_), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n766_), .A2(new_n771_), .B1(new_n241_), .B2(new_n205_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(new_n609_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n590_), .A2(KEYINPUT114), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n586_), .A2(new_n591_), .A3(new_n592_), .A4(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n569_), .B1(new_n507_), .B2(new_n525_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n592_), .B(new_n591_), .C1(KEYINPUT12), .C2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n775_), .B1(new_n779_), .B2(new_n774_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n589_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n782_), .A2(KEYINPUT56), .A3(new_n599_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n782_), .B2(new_n599_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT58), .B(new_n773_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT117), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n773_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  INV_X1    g589(.A(new_n777_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n591_), .B1(new_n778_), .B2(KEYINPUT12), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n585_), .B(new_n569_), .C1(new_n507_), .C2(new_n532_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n774_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT55), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n795_), .B2(new_n593_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n790_), .B1(new_n796_), .B2(new_n600_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n782_), .A2(KEYINPUT56), .A3(new_n599_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n799_), .A2(new_n800_), .A3(KEYINPUT58), .A4(new_n773_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n617_), .A2(new_n626_), .A3(new_n624_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n786_), .A2(new_n789_), .A3(new_n801_), .A4(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n245_), .A2(KEYINPUT113), .A3(new_n609_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT113), .B1(new_n245_), .B2(new_n609_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n608_), .A2(new_n609_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n799_), .A2(new_n807_), .B1(new_n808_), .B2(new_n772_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n562_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n804_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n806_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n245_), .A2(KEYINPUT113), .A3(new_n609_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n812_), .B(new_n813_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n808_), .A2(new_n772_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(KEYINPUT57), .A3(new_n562_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n803_), .A2(new_n811_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n581_), .ZN(new_n819_));
  AND4_X1   g618(.A1(KEYINPUT112), .A2(new_n631_), .A3(new_n246_), .A4(new_n628_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT112), .B1(new_n612_), .B2(new_n246_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n627_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT54), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n824_), .B(new_n627_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n819_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT118), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n818_), .A2(new_n581_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n462_), .A2(new_n468_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n695_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n828_), .A2(new_n473_), .A3(new_n831_), .A4(new_n834_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n835_), .A2(new_n246_), .ZN(new_n836_));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  NOR4_X1   g636(.A1(new_n829_), .A2(KEYINPUT59), .A3(new_n383_), .A4(new_n833_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n835_), .B2(KEYINPUT59), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n246_), .A2(new_n837_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n836_), .A2(new_n837_), .B1(new_n839_), .B2(new_n840_), .ZN(G1340gat));
  AOI211_X1 g640(.A(new_n631_), .B(new_n838_), .C1(new_n835_), .C2(KEYINPUT59), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT119), .B(G120gat), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n828_), .A2(new_n473_), .A3(new_n831_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n844_), .B1(new_n631_), .B2(KEYINPUT60), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n834_), .A3(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n844_), .A2(KEYINPUT60), .ZN(new_n849_));
  OAI22_X1  g648(.A1(new_n842_), .A2(new_n844_), .B1(new_n848_), .B2(new_n849_), .ZN(G1341gat));
  OR2_X1    g649(.A1(new_n835_), .A2(new_n581_), .ZN(new_n851_));
  INV_X1    g650(.A(G127gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n581_), .A2(new_n852_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n851_), .A2(new_n852_), .B1(new_n839_), .B2(new_n853_), .ZN(G1342gat));
  OR2_X1    g653(.A1(new_n835_), .A2(new_n562_), .ZN(new_n855_));
  INV_X1    g654(.A(G134gat), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n627_), .A2(new_n856_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n855_), .A2(new_n856_), .B1(new_n839_), .B2(new_n857_), .ZN(G1343gat));
  NOR2_X1   g657(.A1(new_n695_), .A2(new_n473_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n828_), .A2(new_n831_), .A3(new_n832_), .A4(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n245_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g662(.A1(new_n860_), .A2(new_n631_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT120), .B(G148gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1345gat));
  NOR2_X1   g665(.A1(new_n860_), .A2(new_n581_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT61), .B(G155gat), .Z(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  AOI21_X1  g668(.A(G162gat), .B1(new_n861_), .B2(new_n810_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n306_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n861_), .B2(new_n871_), .ZN(G1347gat));
  AOI21_X1  g671(.A(new_n246_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n472_), .A2(new_n462_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n819_), .B2(new_n826_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT121), .B1(new_n875_), .B2(new_n473_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  NOR4_X1   g676(.A1(new_n829_), .A2(new_n877_), .A3(new_n383_), .A4(new_n874_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n873_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n874_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n827_), .A2(new_n245_), .A3(new_n473_), .A4(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n881_), .A2(new_n882_), .A3(G169gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(G169gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n879_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT122), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n879_), .B(new_n887_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1348gat));
  NAND2_X1  g688(.A1(new_n845_), .A2(KEYINPUT123), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n828_), .A2(new_n891_), .A3(new_n831_), .A4(new_n473_), .ZN(new_n892_));
  INV_X1    g691(.A(G176gat), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n631_), .A2(new_n893_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n890_), .A2(new_n880_), .A3(new_n892_), .A4(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n876_), .A2(new_n878_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n893_), .B1(new_n896_), .B2(new_n631_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1349gat));
  NOR3_X1   g697(.A1(new_n896_), .A2(new_n275_), .A3(new_n581_), .ZN(new_n899_));
  INV_X1    g698(.A(G183gat), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n890_), .A2(new_n628_), .A3(new_n880_), .A4(new_n892_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1350gat));
  OAI21_X1  g701(.A(G190gat), .B1(new_n896_), .B2(new_n627_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n810_), .A2(new_n276_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n896_), .B2(new_n904_), .ZN(G1351gat));
  NAND3_X1  g704(.A1(new_n302_), .A2(new_n468_), .A3(new_n383_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n467_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n828_), .A2(new_n831_), .A3(new_n908_), .A4(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n346_), .B1(new_n910_), .B2(new_n246_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n910_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n914_), .A2(G197gat), .A3(new_n245_), .ZN(new_n915_));
  OAI211_X1 g714(.A(KEYINPUT125), .B(new_n346_), .C1(new_n910_), .C2(new_n246_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n913_), .A2(new_n915_), .A3(new_n916_), .ZN(G1352gat));
  NOR2_X1   g716(.A1(new_n910_), .A2(new_n631_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT126), .B(G204gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1353gat));
  AOI211_X1 g719(.A(KEYINPUT63), .B(G211gat), .C1(new_n914_), .C2(new_n628_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT63), .B(G211gat), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n910_), .A2(new_n581_), .A3(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1354gat));
  XOR2_X1   g723(.A(KEYINPUT127), .B(G218gat), .Z(new_n925_));
  NOR3_X1   g724(.A1(new_n910_), .A2(new_n627_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n914_), .A2(new_n810_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n925_), .ZN(G1355gat));
endmodule


