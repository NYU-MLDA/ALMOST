//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT65), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n202_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(KEYINPUT65), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n203_), .A2(KEYINPUT6), .ZN(new_n209_));
  AND2_X1   g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT66), .ZN(new_n212_));
  OAI22_X1  g011(.A1(new_n212_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT7), .ZN(new_n214_));
  INV_X1    g013(.A(G99gat), .ZN(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .A4(KEYINPUT66), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n207_), .A2(new_n211_), .A3(new_n213_), .A4(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT68), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  INV_X1    g022(.A(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n219_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n218_), .A2(KEYINPUT67), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(new_n230_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n218_), .A2(new_n228_), .A3(KEYINPUT67), .A4(new_n233_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n217_), .A2(new_n213_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n210_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n222_), .A2(new_n227_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n232_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n225_), .A2(KEYINPUT9), .A3(new_n219_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n243_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n244_));
  OR2_X1    g043(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n245_), .A2(KEYINPUT64), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT64), .B1(new_n245_), .B2(new_n246_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n216_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n231_), .A2(new_n234_), .A3(new_n240_), .A4(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G57gat), .B(G64gat), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(KEYINPUT11), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(KEYINPUT11), .ZN(new_n256_));
  XOR2_X1   g055(.A(G71gat), .B(G78gat), .Z(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n256_), .A2(new_n257_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n218_), .A2(new_n228_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n262_), .A2(new_n232_), .B1(new_n244_), .B2(new_n249_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n263_), .A2(KEYINPUT72), .A3(new_n231_), .A4(new_n234_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n253_), .A2(KEYINPUT12), .A3(new_n261_), .A4(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n263_), .A2(new_n260_), .A3(new_n231_), .A4(new_n234_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G230gat), .A2(G233gat), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n240_), .A2(new_n234_), .A3(new_n250_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n229_), .A2(new_n230_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n261_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT73), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n274_));
  AOI211_X1 g073(.A(new_n274_), .B(KEYINPUT12), .C1(new_n251_), .C2(new_n261_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n265_), .B(new_n268_), .C1(new_n273_), .C2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G120gat), .B(G148gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT5), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G176gat), .B(G204gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n269_), .A2(new_n270_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n260_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n266_), .A2(KEYINPUT70), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n282_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n271_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n266_), .B(new_n284_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n282_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n276_), .B(new_n281_), .C1(new_n292_), .C2(new_n267_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n267_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n276_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n280_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT13), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(KEYINPUT74), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n298_), .A2(KEYINPUT74), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n297_), .B1(new_n301_), .B2(new_n299_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT79), .ZN(new_n304_));
  XOR2_X1   g103(.A(G29gat), .B(G36gat), .Z(new_n305_));
  XOR2_X1   g104(.A(G43gat), .B(G50gat), .Z(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  XNOR2_X1  g106(.A(G15gat), .B(G22gat), .ZN(new_n308_));
  INV_X1    g107(.A(G1gat), .ZN(new_n309_));
  INV_X1    g108(.A(G8gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT14), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G1gat), .B(G8gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n307_), .B(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n307_), .A2(KEYINPUT15), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n305_), .B(new_n306_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT15), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n314_), .A3(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n307_), .A2(new_n314_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n316_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G113gat), .B(G141gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G169gat), .B(G197gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n304_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n318_), .A2(new_n325_), .A3(KEYINPUT79), .A4(new_n329_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n330_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT80), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(KEYINPUT80), .A3(new_n334_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n303_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n343_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G155gat), .B(G162gat), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n342_), .B(new_n344_), .C1(KEYINPUT1), .C2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n340_), .B(KEYINPUT3), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT2), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT90), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n345_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n353_), .B2(new_n352_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n348_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G127gat), .B(G134gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT86), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G113gat), .B(G120gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n357_), .A2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n356_), .A2(new_n361_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G1gat), .B(G29gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G57gat), .B(G85gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT102), .B1(new_n366_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n356_), .B(new_n362_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n365_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT102), .ZN(new_n376_));
  INV_X1    g175(.A(new_n371_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n373_), .A2(KEYINPUT4), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n356_), .A2(new_n380_), .A3(new_n361_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n381_), .A2(KEYINPUT100), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(KEYINPUT100), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n379_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n372_), .B(new_n378_), .C1(new_n384_), .C2(new_n374_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G197gat), .B(G204gat), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT21), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G211gat), .B(G218gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G197gat), .B(G204gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT21), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n393_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT91), .ZN(new_n399_));
  INV_X1    g198(.A(new_n394_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n393_), .B1(KEYINPUT92), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(KEYINPUT92), .B2(new_n400_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(KEYINPUT93), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(KEYINPUT93), .ZN(new_n406_));
  INV_X1    g205(.A(G169gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT22), .B1(new_n407_), .B2(KEYINPUT81), .ZN(new_n408_));
  INV_X1    g207(.A(G176gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT22), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G169gat), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n408_), .B(new_n409_), .C1(KEYINPUT81), .C2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G169gat), .A2(G176gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G183gat), .A2(G190gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT23), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(G183gat), .B2(G190gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n407_), .A2(new_n409_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n420_), .A2(KEYINPUT24), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT25), .B(G183gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT26), .B(G190gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n420_), .A2(KEYINPUT24), .A3(new_n415_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n419_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n405_), .A2(new_n406_), .A3(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G226gat), .A2(G233gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT20), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT22), .B(G169gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n409_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n418_), .A2(new_n415_), .A3(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT98), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n425_), .A2(new_n426_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT97), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n422_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n399_), .A2(new_n402_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n433_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n429_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n406_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n427_), .B(new_n419_), .C1(new_n446_), .C2(new_n404_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n441_), .B2(new_n403_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n391_), .B(new_n445_), .C1(new_n450_), .C2(new_n432_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n445_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n432_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n390_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n385_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n379_), .B(new_n374_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n373_), .A2(new_n365_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n371_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n458_), .A2(new_n459_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n455_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n391_), .A2(KEYINPUT32), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n447_), .A2(new_n432_), .A3(new_n449_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n440_), .A2(new_n436_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n448_), .B1(new_n465_), .B2(new_n443_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n432_), .B1(new_n429_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n463_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n445_), .B1(new_n450_), .B2(new_n432_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(new_n463_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n456_), .A2(new_n457_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n377_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n470_), .B1(new_n458_), .B2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G22gat), .B(G50gat), .ZN(new_n474_));
  AND2_X1   g273(.A1(G228gat), .A2(G233gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n356_), .A2(KEYINPUT29), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n403_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n476_), .A2(new_n477_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n475_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n482_));
  INV_X1    g281(.A(new_n475_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n405_), .A2(new_n406_), .A3(new_n483_), .A4(new_n476_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n482_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n474_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n481_), .A2(new_n484_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT95), .ZN(new_n490_));
  INV_X1    g289(.A(new_n474_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n485_), .A3(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n356_), .A2(KEYINPUT29), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT28), .Z(new_n494_));
  XOR2_X1   g293(.A(G78gat), .B(G106gat), .Z(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n488_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n498_));
  OAI22_X1  g297(.A1(new_n462_), .A2(new_n473_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n488_), .A2(new_n492_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n390_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT27), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n452_), .A2(new_n453_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n505_), .B2(new_n391_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n451_), .A2(new_n454_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n503_), .A2(new_n506_), .B1(new_n507_), .B2(new_n504_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n472_), .A2(new_n458_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n488_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n502_), .A2(new_n508_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n499_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n428_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G71gat), .B(G99gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(G43gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G227gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT83), .B(G15gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  OR3_X1    g321(.A1(new_n515_), .A2(new_n516_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n515_), .A2(new_n522_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT84), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n516_), .B1(new_n515_), .B2(new_n522_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n515_), .A2(KEYINPUT84), .A3(new_n522_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n523_), .A2(new_n526_), .A3(new_n527_), .A4(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT87), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT31), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT31), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(KEYINPUT87), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n362_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n531_), .A2(new_n361_), .A3(new_n533_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n513_), .A2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n508_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n510_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n339_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT34), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n545_), .A2(KEYINPUT35), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(KEYINPUT35), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n546_), .B1(new_n547_), .B2(KEYINPUT77), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n283_), .A2(KEYINPUT75), .A3(new_n320_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT75), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(new_n251_), .B2(new_n307_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n548_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(KEYINPUT77), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n253_), .A2(new_n319_), .A3(new_n322_), .A4(new_n264_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT76), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n557_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n555_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(KEYINPUT76), .A3(new_n562_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT78), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(KEYINPUT37), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n570_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(KEYINPUT78), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n260_), .B(new_n314_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583_));
  XOR2_X1   g382(.A(G127gat), .B(G155gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT16), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n582_), .A2(new_n583_), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(KEYINPUT17), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n582_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n578_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n543_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n309_), .A3(new_n509_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT38), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n572_), .B1(new_n538_), .B2(new_n542_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n339_), .A2(new_n591_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G1gat), .B1(new_n600_), .B2(new_n510_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n596_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n601_), .A3(new_n602_), .ZN(G1324gat));
  INV_X1    g402(.A(new_n508_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n594_), .A2(new_n310_), .A3(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n598_), .A2(new_n604_), .A3(new_n599_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n606_), .A2(G8gat), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n606_), .B2(G8gat), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g410(.A(G15gat), .B1(new_n600_), .B2(new_n537_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n593_), .A2(G15gat), .A3(new_n537_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT105), .Z(G1326gat));
  NAND2_X1  g417(.A1(new_n502_), .A2(new_n511_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G22gat), .B1(new_n600_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT42), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n619_), .A2(G22gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n593_), .B2(new_n622_), .ZN(G1327gat));
  INV_X1    g422(.A(new_n591_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n576_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n543_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n509_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n537_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n499_), .B2(new_n512_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n578_), .B1(new_n630_), .B2(new_n541_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT43), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n633_), .B(new_n578_), .C1(new_n630_), .C2(new_n541_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n339_), .A2(new_n624_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT44), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638_));
  INV_X1    g437(.A(new_n636_), .ZN(new_n639_));
  AOI211_X1 g438(.A(new_n638_), .B(new_n639_), .C1(new_n632_), .C2(new_n634_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n509_), .A2(G29gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n628_), .B1(new_n641_), .B2(new_n642_), .ZN(G1328gat));
  INV_X1    g442(.A(KEYINPUT46), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT107), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT107), .ZN(new_n646_));
  INV_X1    g445(.A(G36gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n641_), .B2(new_n604_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n508_), .A2(G36gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT106), .B1(new_n626_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n543_), .A2(new_n652_), .A3(new_n625_), .A4(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT45), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n651_), .A2(KEYINPUT45), .A3(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n645_), .B(new_n646_), .C1(new_n648_), .C2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n637_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n640_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n604_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G36gat), .ZN(new_n663_));
  INV_X1    g462(.A(new_n657_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT45), .B1(new_n651_), .B2(new_n653_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n663_), .A2(new_n666_), .A3(KEYINPUT107), .A4(new_n644_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n659_), .A2(new_n667_), .ZN(G1329gat));
  AOI21_X1  g467(.A(G43gat), .B1(new_n627_), .B2(new_n629_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n629_), .A2(G43gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n641_), .B2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g471(.A(new_n619_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G50gat), .B1(new_n627_), .B2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(G50gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n641_), .B2(new_n675_), .ZN(G1331gat));
  NOR2_X1   g475(.A1(new_n303_), .A2(new_n338_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n598_), .A2(new_n624_), .A3(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G57gat), .B1(new_n678_), .B2(new_n510_), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n338_), .B(new_n303_), .C1(new_n538_), .C2(new_n542_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n592_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n510_), .A2(G57gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(G1332gat));
  OAI21_X1  g482(.A(G64gat), .B1(new_n678_), .B2(new_n508_), .ZN(new_n684_));
  XOR2_X1   g483(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n508_), .A2(G64gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n681_), .B2(new_n687_), .ZN(G1333gat));
  OAI21_X1  g487(.A(G71gat), .B1(new_n678_), .B2(new_n537_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT49), .ZN(new_n690_));
  OR3_X1    g489(.A1(new_n681_), .A2(G71gat), .A3(new_n537_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT109), .ZN(G1334gat));
  OAI21_X1  g492(.A(G78gat), .B1(new_n678_), .B2(new_n619_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT50), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n619_), .A2(G78gat), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT110), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n695_), .B1(new_n681_), .B2(new_n697_), .ZN(G1335gat));
  AND3_X1   g497(.A1(new_n635_), .A2(new_n591_), .A3(new_n677_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G85gat), .B1(new_n700_), .B2(new_n510_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n680_), .A2(new_n625_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(new_n223_), .A3(new_n509_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1336gat));
  OAI21_X1  g504(.A(G92gat), .B1(new_n700_), .B2(new_n508_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n703_), .A2(new_n224_), .A3(new_n604_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1337gat));
  OAI211_X1 g507(.A(new_n703_), .B(new_n629_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n700_), .A2(new_n537_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(new_n215_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT51), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n713_), .B(new_n709_), .C1(new_n710_), .C2(new_n215_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1338gat));
  NAND3_X1  g514(.A1(new_n703_), .A2(new_n216_), .A3(new_n673_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n635_), .A2(new_n591_), .A3(new_n673_), .A4(new_n677_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(new_n718_), .A3(G106gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n717_), .B2(G106gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g521(.A(new_n338_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n723_), .A2(new_n624_), .A3(new_n577_), .A4(new_n574_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT54), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT113), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n290_), .B(new_n265_), .C1(new_n273_), .C2(new_n275_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n267_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT55), .ZN(new_n730_));
  AOI22_X1  g529(.A1(new_n728_), .A2(new_n729_), .B1(new_n276_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n271_), .A2(new_n272_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n274_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n271_), .A2(KEYINPUT73), .A3(new_n272_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n735_), .A2(KEYINPUT55), .A3(new_n265_), .A4(new_n268_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n281_), .B1(new_n731_), .B2(new_n736_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT112), .B(KEYINPUT56), .Z(new_n738_));
  OAI21_X1  g537(.A(new_n727_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n265_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n290_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n729_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n276_), .A2(new_n730_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n736_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n280_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n738_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(KEYINPUT113), .A3(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n280_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT114), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n744_), .A2(new_n750_), .A3(KEYINPUT56), .A4(new_n280_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n739_), .A2(new_n747_), .A3(new_n749_), .A4(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n337_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(new_n335_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n294_), .A2(new_n295_), .A3(new_n280_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT111), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n338_), .A2(new_n293_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n752_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT115), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n752_), .A2(new_n759_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n315_), .A2(new_n316_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n323_), .A2(new_n324_), .A3(new_n317_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n330_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n333_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n297_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT117), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n297_), .A2(new_n772_), .A3(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n761_), .A2(new_n763_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n572_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n769_), .A2(new_n293_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n737_), .A2(KEYINPUT56), .ZN(new_n780_));
  INV_X1    g579(.A(new_n748_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(new_n578_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n782_), .A2(new_n783_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n760_), .A2(KEYINPUT115), .B1(new_n771_), .B2(new_n773_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n572_), .B1(new_n788_), .B2(new_n763_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n778_), .B(new_n787_), .C1(new_n789_), .C2(KEYINPUT57), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n726_), .B1(new_n790_), .B2(new_n591_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n539_), .A2(new_n537_), .A3(new_n510_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G113gat), .B1(new_n794_), .B2(new_n338_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n795_), .A2(KEYINPUT118), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(KEYINPUT118), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n775_), .A2(new_n576_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n776_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n775_), .A2(new_n777_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n624_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT59), .B(new_n792_), .C1(new_n803_), .C2(new_n726_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n799_), .A2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT119), .B(G113gat), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n754_), .A2(new_n806_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n796_), .A2(new_n797_), .B1(new_n805_), .B2(new_n807_), .ZN(G1340gat));
  OR2_X1    g607(.A1(new_n303_), .A2(KEYINPUT60), .ZN(new_n809_));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n794_), .B(new_n811_), .C1(KEYINPUT60), .C2(new_n810_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n303_), .B1(new_n799_), .B2(new_n804_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT120), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n812_), .C1(new_n813_), .C2(new_n810_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1341gat));
  INV_X1    g617(.A(G127gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n794_), .A2(new_n819_), .A3(new_n624_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n591_), .B1(new_n799_), .B2(new_n804_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n819_), .ZN(G1342gat));
  AOI21_X1  g621(.A(G134gat), .B1(new_n794_), .B2(new_n572_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n578_), .ZN(new_n824_));
  XOR2_X1   g623(.A(KEYINPUT121), .B(G134gat), .Z(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n823_), .B1(new_n805_), .B2(new_n826_), .ZN(G1343gat));
  INV_X1    g626(.A(new_n791_), .ZN(new_n828_));
  NOR4_X1   g627(.A1(new_n629_), .A2(new_n619_), .A3(new_n604_), .A4(new_n510_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(new_n754_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT122), .B(G141gat), .Z(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1344gat));
  NOR2_X1   g632(.A1(new_n830_), .A2(new_n303_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(G148gat), .Z(G1345gat));
  OAI21_X1  g634(.A(KEYINPUT123), .B1(new_n830_), .B2(new_n591_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n828_), .A2(new_n837_), .A3(new_n624_), .A4(new_n829_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT61), .B(G155gat), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n836_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1346gat));
  INV_X1    g641(.A(G162gat), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n830_), .A2(new_n843_), .A3(new_n824_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n830_), .B2(new_n576_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT124), .B(new_n843_), .C1(new_n830_), .C2(new_n576_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n844_), .B1(new_n847_), .B2(new_n848_), .ZN(G1347gat));
  INV_X1    g648(.A(KEYINPUT126), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n673_), .A2(new_n508_), .A3(new_n540_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n828_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n850_), .B1(new_n828_), .B2(new_n851_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n434_), .B(new_n338_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n828_), .A2(new_n851_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G169gat), .B1(new_n856_), .B2(new_n754_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n858_), .A2(KEYINPUT125), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(KEYINPUT125), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n857_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n855_), .B(new_n861_), .C1(new_n857_), .C2(new_n859_), .ZN(G1348gat));
  INV_X1    g661(.A(new_n854_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n852_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n303_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n409_), .A3(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(G176gat), .B1(new_n856_), .B2(new_n303_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1349gat));
  NOR2_X1   g667(.A1(new_n856_), .A2(new_n591_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(G183gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n591_), .A2(new_n423_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n864_), .B2(new_n871_), .ZN(G1350gat));
  OAI211_X1 g671(.A(new_n572_), .B(new_n424_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n824_), .B1(new_n863_), .B2(new_n852_), .ZN(new_n874_));
  INV_X1    g673(.A(G190gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1351gat));
  NOR4_X1   g675(.A1(new_n629_), .A2(new_n619_), .A3(new_n509_), .A4(new_n508_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n828_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n338_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n865_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g682(.A1(new_n828_), .A2(new_n624_), .A3(new_n877_), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT63), .B(G211gat), .Z(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT127), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n884_), .A2(KEYINPUT127), .A3(new_n886_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1354gat));
  OAI21_X1  g691(.A(G218gat), .B1(new_n878_), .B2(new_n824_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n576_), .A2(G218gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n878_), .B2(new_n894_), .ZN(G1355gat));
endmodule


