//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT89), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT90), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n202_), .A2(new_n203_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n205_), .B(KEYINPUT90), .ZN(new_n210_));
  INV_X1    g009(.A(new_n208_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G141gat), .ZN(new_n214_));
  INV_X1    g013(.A(G148gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT94), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT93), .A2(KEYINPUT2), .ZN(new_n219_));
  AND2_X1   g018(.A1(KEYINPUT93), .A2(KEYINPUT2), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n217_), .B(new_n218_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n214_), .A2(new_n215_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT92), .A2(KEYINPUT3), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n220_), .A2(new_n219_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT94), .B1(new_n225_), .B2(new_n216_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n216_), .A2(KEYINPUT2), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n221_), .A2(new_n224_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT91), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n230_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n231_), .B(KEYINPUT1), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n222_), .B(new_n217_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(KEYINPUT95), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT95), .B1(new_n232_), .B2(new_n235_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n213_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n232_), .A2(new_n235_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n211_), .B2(new_n204_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(KEYINPUT102), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT102), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n213_), .B(new_n245_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n243_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n241_), .B1(new_n247_), .B2(new_n240_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  AOI211_X1 g050(.A(new_n250_), .B(new_n243_), .C1(new_n244_), .C2(new_n246_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G57gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G85gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(G1gat), .B(G29gat), .Z(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT33), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n262_));
  OR3_X1    g061(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n263_));
  INV_X1    g062(.A(G190gat), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n264_), .A2(KEYINPUT26), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(KEYINPUT26), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT25), .B(G183gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G183gat), .ZN(new_n270_));
  OR3_X1    g069(.A1(new_n270_), .A2(new_n264_), .A3(KEYINPUT23), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT23), .B1(new_n270_), .B2(new_n264_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AND4_X1   g076(.A1(new_n263_), .A2(new_n269_), .A3(new_n273_), .A4(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n276_), .B(KEYINPUT84), .Z(new_n279_));
  OR2_X1    g078(.A1(new_n272_), .A2(KEYINPUT85), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n272_), .A2(KEYINPUT85), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n271_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n270_), .A2(new_n264_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n279_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT86), .B(G176gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT22), .B(G169gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n278_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT97), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G211gat), .A2(G218gat), .ZN(new_n290_));
  AND2_X1   g089(.A1(G211gat), .A2(G218gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(G197gat), .B(G204gat), .Z(new_n292_));
  OAI221_X1 g091(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .C1(new_n292_), .C2(KEYINPUT21), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(KEYINPUT21), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n262_), .B1(new_n288_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n295_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT87), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n287_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT81), .B(G183gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n264_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n279_), .B1(new_n273_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n279_), .A2(new_n274_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G183gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT82), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n265_), .B1(KEYINPUT83), .B2(new_n266_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n300_), .A2(KEYINPUT25), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n266_), .A2(KEYINPUT83), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .A4(new_n310_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n304_), .A2(new_n311_), .A3(new_n263_), .A4(new_n282_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n303_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n297_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n296_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT19), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n288_), .A2(new_n295_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n295_), .A2(new_n312_), .A3(new_n303_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n320_), .A2(KEYINPUT20), .A3(new_n317_), .A4(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G8gat), .B(G36gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G64gat), .B(G92gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n323_), .A2(new_n328_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI211_X1 g131(.A(new_n249_), .B(new_n243_), .C1(new_n244_), .C2(new_n246_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n334_), .B2(new_n257_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n251_), .A2(KEYINPUT33), .A3(new_n253_), .A4(new_n258_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n261_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT32), .ZN(new_n338_));
  INV_X1    g137(.A(new_n328_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n323_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AND4_X1   g139(.A1(KEYINPUT20), .A2(new_n320_), .A3(new_n318_), .A4(new_n321_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n318_), .B1(new_n296_), .B2(new_n314_), .ZN(new_n342_));
  OAI211_X1 g141(.A(KEYINPUT32), .B(new_n328_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n258_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n344_));
  AOI211_X1 g143(.A(new_n257_), .B(new_n252_), .C1(new_n248_), .C2(new_n250_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n340_), .B(new_n343_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n337_), .A2(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n209_), .A2(new_n212_), .A3(KEYINPUT31), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT31), .B1(new_n209_), .B2(new_n212_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT88), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n303_), .A2(new_n353_), .A3(new_n312_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n353_), .B1(new_n303_), .B2(new_n312_), .ZN(new_n356_));
  OAI21_X1  g155(.A(G43gat), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G227gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(G15gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n313_), .A2(KEYINPUT30), .ZN(new_n361_));
  INV_X1    g160(.A(G43gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(new_n354_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n357_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n360_), .B1(new_n357_), .B2(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n352_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n351_), .A3(new_n364_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n237_), .A2(new_n238_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT28), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n238_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(new_n378_), .A3(new_n236_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n380_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n385_), .A3(KEYINPUT99), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n381_), .A2(new_n385_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(KEYINPUT96), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(KEYINPUT96), .A2(G233gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(G228gat), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n378_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n396_), .B2(new_n295_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT98), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n297_), .B(new_n394_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT100), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n388_), .B(new_n390_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n388_), .A2(new_n390_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n403_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n401_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n376_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n330_), .A2(KEYINPUT27), .A3(new_n331_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n339_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n412_), .A2(KEYINPUT103), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(KEYINPUT103), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n329_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n411_), .B1(new_n415_), .B2(KEYINPUT27), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n375_), .A2(new_n408_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n373_), .A2(new_n404_), .A3(new_n407_), .A4(new_n374_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n344_), .A2(new_n345_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n347_), .A2(new_n410_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT16), .B(G183gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(G211gat), .ZN(new_n423_));
  XOR2_X1   g222(.A(G127gat), .B(G155gat), .Z(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n426_));
  OR2_X1    g225(.A1(G57gat), .A2(G64gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G57gat), .A2(G64gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT11), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G71gat), .B(G78gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT11), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n427_), .A2(new_n433_), .A3(new_n428_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n426_), .B(new_n432_), .C1(new_n435_), .C2(new_n431_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n426_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n431_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n431_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(KEYINPUT11), .B2(new_n429_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n437_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G1gat), .B(G8gat), .ZN(new_n443_));
  AND2_X1   g242(.A1(G15gat), .A2(G22gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G15gat), .A2(G22gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT14), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(G1gat), .B2(G8gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n443_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(G1gat), .A2(G8gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G1gat), .A2(G8gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G15gat), .B(G22gat), .ZN(new_n453_));
  INV_X1    g252(.A(G1gat), .ZN(new_n454_));
  INV_X1    g253(.A(G8gat), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT14), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n449_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n442_), .B(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G231gat), .A2(G233gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT75), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n425_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT17), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n464_), .B1(new_n461_), .B2(new_n425_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n465_), .B1(new_n467_), .B2(new_n463_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n421_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT15), .ZN(new_n470_));
  INV_X1    g269(.A(G50gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G43gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n362_), .A2(G50gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(G29gat), .A2(G36gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G29gat), .A2(G36gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n472_), .B(new_n473_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n470_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n479_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G43gat), .B(G50gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G29gat), .B(G36gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n480_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n484_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT15), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n483_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G85gat), .B(G92gat), .Z(new_n493_));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n494_));
  INV_X1    g293(.A(G99gat), .ZN(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n493_), .B1(new_n499_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT10), .B(G99gat), .ZN(new_n508_));
  OR3_X1    g307(.A1(new_n508_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n493_), .A2(KEYINPUT9), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G85gat), .A2(G92gat), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n511_), .A2(KEYINPUT9), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n504_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT64), .B1(new_n508_), .B2(G106gat), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n505_), .A2(new_n506_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n507_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n492_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT71), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G232gat), .A2(G233gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT34), .Z(new_n521_));
  INV_X1    g320(.A(KEYINPUT35), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(KEYINPUT66), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n507_), .A2(new_n525_), .A3(new_n516_), .A4(new_n515_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(new_n490_), .A3(new_n489_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n519_), .A2(new_n523_), .A3(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n521_), .A2(new_n522_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT72), .B(G134gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(G162gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(KEYINPUT36), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n529_), .A2(new_n530_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n531_), .A2(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(KEYINPUT36), .ZN(new_n542_));
  INV_X1    g341(.A(new_n536_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n538_), .A2(new_n539_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n540_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT37), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT74), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n541_), .A2(KEYINPUT74), .A3(new_n542_), .A4(new_n543_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .A4(new_n538_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n469_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n442_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n527_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n524_), .A2(new_n442_), .A3(new_n526_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(G230gat), .A3(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n442_), .A2(KEYINPUT12), .A3(new_n517_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n561_), .A2(new_n556_), .A3(new_n562_), .A4(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G120gat), .B(G148gat), .ZN(new_n565_));
  INV_X1    g364(.A(G204gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT5), .ZN(new_n568_));
  INV_X1    g367(.A(G176gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n559_), .A2(new_n564_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n559_), .B2(new_n564_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT13), .Z(new_n575_));
  INV_X1    g374(.A(KEYINPUT78), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT76), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n449_), .A2(new_n457_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n490_), .B2(new_n489_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n481_), .A2(new_n482_), .A3(new_n458_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n578_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n489_), .A2(new_n579_), .A3(new_n490_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n458_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n584_), .A3(KEYINPUT76), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n577_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n481_), .A2(new_n482_), .A3(new_n470_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT15), .B1(new_n489_), .B2(new_n490_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT77), .B(new_n458_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n579_), .B1(new_n483_), .B2(new_n491_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT77), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n581_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n589_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n586_), .B1(new_n577_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595_));
  INV_X1    g394(.A(G169gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(G197gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n576_), .B1(new_n594_), .B2(new_n599_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n492_), .A2(new_n458_), .B1(KEYINPUT77), .B2(new_n583_), .ZN(new_n601_));
  AOI211_X1 g400(.A(new_n591_), .B(new_n579_), .C1(new_n483_), .C2(new_n491_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n577_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n577_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n585_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT76), .B1(new_n583_), .B2(new_n584_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n604_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n599_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(KEYINPUT78), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n600_), .A2(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n603_), .A2(new_n607_), .A3(new_n599_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT79), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT79), .ZN(new_n615_));
  AOI211_X1 g414(.A(new_n615_), .B(new_n612_), .C1(new_n600_), .C2(new_n610_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(KEYINPUT80), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n614_), .A2(new_n616_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT80), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n554_), .A2(new_n575_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n420_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n454_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT38), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n575_), .A2(new_n619_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n469_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n549_), .A2(new_n551_), .A3(new_n538_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n420_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n627_), .A2(new_n634_), .ZN(G1324gat));
  INV_X1    g434(.A(new_n416_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n629_), .A2(new_n631_), .A3(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n455_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT104), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(KEYINPUT104), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n624_), .A2(new_n455_), .A3(new_n416_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT104), .B(new_n639_), .C1(new_n637_), .C2(new_n455_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT105), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n642_), .A2(new_n647_), .A3(new_n643_), .A4(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n646_), .A2(KEYINPUT40), .A3(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1325gat));
  AOI21_X1  g452(.A(new_n359_), .B1(new_n632_), .B2(new_n375_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT106), .Z(new_n655_));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n656_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n624_), .A2(new_n359_), .A3(new_n375_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(G1326gat));
  INV_X1    g459(.A(G22gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n408_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n632_), .B2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT42), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n624_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  INV_X1    g466(.A(new_n628_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n347_), .A2(new_n410_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n418_), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n374_), .A2(new_n373_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n420_), .B(new_n636_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n553_), .B1(new_n669_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT107), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n553_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n672_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n409_), .B1(new_n337_), .B2(new_n346_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(KEYINPUT43), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n675_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT108), .B1(new_n679_), .B2(KEYINPUT43), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n669_), .A2(new_n672_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n674_), .A4(new_n676_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n668_), .B1(new_n682_), .B2(new_n687_), .ZN(new_n688_));
  AOI211_X1 g487(.A(KEYINPUT109), .B(new_n667_), .C1(new_n688_), .C2(new_n468_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n681_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n680_), .B1(new_n679_), .B2(KEYINPUT43), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n692_));
  NOR4_X1   g491(.A1(new_n421_), .A2(KEYINPUT108), .A3(KEYINPUT43), .A4(new_n553_), .ZN(new_n693_));
  OAI22_X1  g492(.A1(new_n690_), .A2(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n667_), .A2(KEYINPUT109), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n694_), .A2(new_n628_), .A3(new_n468_), .A4(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n667_), .A2(KEYINPUT109), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n625_), .B1(new_n689_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n696_), .A2(new_n697_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n697_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n688_), .A2(new_n468_), .A3(new_n703_), .A4(new_n695_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(KEYINPUT110), .A3(new_n625_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n701_), .A2(G29gat), .A3(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n421_), .A2(new_n630_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n468_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n623_), .A2(new_n575_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n711_), .A2(G29gat), .A3(new_n420_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n707_), .A2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(new_n711_), .ZN(new_n714_));
  INV_X1    g513(.A(G36gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n416_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT45), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n636_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(new_n715_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT46), .B(new_n717_), .C1(new_n718_), .C2(new_n715_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  AOI211_X1 g522(.A(new_n362_), .B(new_n376_), .C1(new_n702_), .C2(new_n704_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n362_), .B1(new_n711_), .B2(new_n376_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT111), .Z(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT47), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n705_), .A2(G43gat), .A3(new_n375_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729_));
  INV_X1    g528(.A(new_n726_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n728_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n731_), .ZN(G1330gat));
  AOI21_X1  g531(.A(G50gat), .B1(new_n714_), .B2(new_n662_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n471_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n662_), .ZN(G1331gat));
  INV_X1    g534(.A(new_n554_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n575_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n737_), .A2(new_n617_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n625_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n469_), .A2(new_n630_), .A3(new_n575_), .A4(new_n623_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(new_n420_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(G57gat), .B2(new_n743_), .ZN(G1332gat));
  OAI21_X1  g543(.A(G64gat), .B1(new_n742_), .B2(new_n636_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT48), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n636_), .A2(G64gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n739_), .B2(new_n747_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT112), .Z(G1333gat));
  OAI21_X1  g548(.A(G71gat), .B1(new_n742_), .B2(new_n376_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT49), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n376_), .A2(G71gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n739_), .B2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n742_), .B2(new_n408_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n408_), .A2(G78gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n739_), .B2(new_n756_), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n738_), .A2(new_n468_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n708_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n625_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n758_), .B1(new_n682_), .B2(new_n687_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n763_), .A2(new_n625_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n764_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g564(.A(G92gat), .B1(new_n761_), .B2(new_n416_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n763_), .A2(G92gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(new_n416_), .ZN(G1337gat));
  AOI21_X1  g567(.A(new_n495_), .B1(new_n763_), .B2(new_n375_), .ZN(new_n769_));
  AND2_X1   g568(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n760_), .A2(new_n508_), .A3(new_n376_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n769_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(G1338gat));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n408_), .B(new_n758_), .C1(new_n682_), .C2(new_n687_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n496_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n763_), .A2(new_n662_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(KEYINPUT114), .A3(G106gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n777_), .A2(new_n779_), .A3(KEYINPUT52), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n761_), .A2(new_n496_), .A3(new_n662_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n775_), .B(new_n782_), .C1(new_n776_), .C2(new_n496_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(new_n781_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT53), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n780_), .A2(new_n786_), .A3(new_n781_), .A4(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1339gat));
  OAI21_X1  g587(.A(new_n571_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n564_), .A2(KEYINPUT117), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n561_), .A2(new_n556_), .A3(new_n563_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n562_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n793_), .B1(new_n564_), .B2(KEYINPUT117), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n795_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n792_), .B1(new_n799_), .B2(new_n570_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n570_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n794_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT56), .B(new_n801_), .C1(new_n803_), .C2(new_n797_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT116), .B(new_n571_), .C1(new_n614_), .C2(new_n616_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n791_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n593_), .A2(new_n577_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n605_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n810_), .A2(new_n609_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n600_), .B2(new_n610_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n574_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n791_), .A2(new_n805_), .A3(KEYINPUT118), .A4(new_n806_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n809_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n630_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(KEYINPUT57), .A3(new_n630_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n805_), .A2(KEYINPUT119), .ZN(new_n821_));
  INV_X1    g620(.A(new_n800_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n572_), .B1(new_n822_), .B2(KEYINPUT119), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n823_), .A3(new_n813_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n825_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n821_), .A2(new_n823_), .A3(new_n813_), .A4(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n676_), .A3(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n819_), .A2(new_n820_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n468_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n622_), .A2(new_n575_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n468_), .B1(new_n547_), .B2(new_n552_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n835_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n832_), .A2(new_n837_), .A3(new_n833_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n836_), .A2(new_n838_), .B1(KEYINPUT115), .B2(KEYINPUT54), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n417_), .B1(new_n831_), .B2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n420_), .A2(new_n416_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n839_), .B1(new_n830_), .B2(new_n468_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  INV_X1    g644(.A(new_n842_), .ZN(new_n846_));
  NOR4_X1   g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n417_), .A4(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(G113gat), .B(new_n622_), .C1(new_n843_), .C2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n841_), .A2(new_n842_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n619_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n848_), .A2(KEYINPUT121), .A3(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1340gat));
  XNOR2_X1  g655(.A(KEYINPUT122), .B(G120gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n841_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n575_), .B2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(KEYINPUT123), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n859_), .A2(new_n864_), .A3(new_n861_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n843_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n847_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n737_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n863_), .A2(new_n865_), .B1(new_n868_), .B2(new_n858_), .ZN(G1341gat));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n850_), .B2(new_n468_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n872_), .ZN(new_n874_));
  OAI211_X1 g673(.A(G127gat), .B(new_n709_), .C1(new_n843_), .C2(new_n847_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(G1342gat));
  INV_X1    g675(.A(new_n850_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G134gat), .B1(new_n877_), .B2(new_n631_), .ZN(new_n878_));
  INV_X1    g677(.A(G134gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n880_), .B2(new_n676_), .ZN(G1343gat));
  NOR3_X1   g680(.A1(new_n844_), .A2(new_n418_), .A3(new_n846_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n617_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT125), .B(G141gat), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n883_), .B(new_n884_), .Z(G1344gat));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n575_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g686(.A1(new_n882_), .A2(new_n709_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1346gat));
  AOI21_X1  g689(.A(G162gat), .B1(new_n882_), .B2(new_n631_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n882_), .A2(G162gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n676_), .B2(new_n892_), .ZN(G1347gat));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n841_), .A2(new_n420_), .A3(new_n416_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n619_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n896_), .B2(new_n596_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n286_), .ZN(new_n898_));
  OAI211_X1 g697(.A(KEYINPUT62), .B(G169gat), .C1(new_n895_), .C2(new_n619_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(G1348gat));
  INV_X1    g699(.A(new_n895_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n575_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n569_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n285_), .B2(new_n902_), .ZN(G1349gat));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n709_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n268_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(new_n300_), .B2(new_n905_), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n895_), .B2(new_n553_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n631_), .A2(new_n267_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n895_), .B2(new_n909_), .ZN(G1351gat));
  NAND2_X1  g709(.A1(new_n831_), .A2(new_n840_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n625_), .A2(KEYINPUT126), .A3(new_n418_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n636_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT126), .B1(new_n625_), .B2(new_n418_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n911_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n911_), .A2(KEYINPUT127), .A3(new_n913_), .A4(new_n914_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n619_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(new_n598_), .ZN(G1352gat));
  AOI21_X1  g719(.A(new_n737_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n566_), .ZN(G1353gat));
  XNOR2_X1  g721(.A(KEYINPUT63), .B(G211gat), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n468_), .B(new_n923_), .C1(new_n917_), .C2(new_n918_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n917_), .A2(new_n918_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n709_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n924_), .B1(new_n926_), .B2(new_n927_), .ZN(G1354gat));
  AOI21_X1  g727(.A(G218gat), .B1(new_n925_), .B2(new_n631_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n925_), .A2(G218gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n676_), .B2(new_n930_), .ZN(G1355gat));
endmodule


