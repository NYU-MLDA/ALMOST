//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n959_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n997_, new_n998_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1011_,
    new_n1012_, new_n1013_, new_n1015_, new_n1016_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT36), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT72), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT73), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT8), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT67), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT7), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n211_), .A2(new_n213_), .A3(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G85gat), .B(G92gat), .Z(new_n221_));
  AOI21_X1  g020(.A(new_n209_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n209_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(KEYINPUT9), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(G85gat), .A3(G92gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n228_), .A3(new_n214_), .ZN(new_n229_));
  INV_X1    g028(.A(G106gat), .ZN(new_n230_));
  OR2_X1    g029(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(KEYINPUT65), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT65), .B1(new_n231_), .B2(new_n232_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n230_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT10), .B(G99gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n233_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(KEYINPUT66), .A3(new_n230_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n229_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n208_), .B1(new_n225_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n229_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT66), .B1(new_n242_), .B2(new_n230_), .ZN(new_n247_));
  AOI211_X1 g046(.A(new_n237_), .B(G106gat), .C1(new_n241_), .C2(new_n233_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n249_), .B(KEYINPUT68), .C1(new_n222_), .C2(new_n224_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G29gat), .B(G36gat), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT70), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(KEYINPUT70), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G43gat), .B(G50gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n252_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT15), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(KEYINPUT15), .A3(new_n258_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n245_), .A2(new_n250_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n245_), .A2(new_n250_), .A3(new_n263_), .A4(KEYINPUT71), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n249_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G232gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT34), .ZN(new_n271_));
  OAI22_X1  g070(.A1(new_n269_), .A2(new_n259_), .B1(KEYINPUT35), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n271_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT35), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n268_), .A2(new_n279_), .A3(new_n273_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n207_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n268_), .B2(new_n273_), .ZN(new_n282_));
  AOI211_X1 g081(.A(new_n277_), .B(new_n272_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT37), .B1(new_n281_), .B2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n278_), .A2(new_n284_), .A3(new_n280_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n206_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT37), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G127gat), .B(G155gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT16), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G183gat), .B(G211gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT74), .B(G1gat), .ZN(new_n300_));
  INV_X1    g099(.A(G8gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT14), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT75), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G15gat), .B(G22gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n303_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n299_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(new_n304_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT75), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(new_n305_), .A3(new_n298_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G231gat), .A2(G233gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(KEYINPUT76), .Z(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n314_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n308_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G57gat), .B(G64gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT11), .ZN(new_n320_));
  XOR2_X1   g119(.A(G71gat), .B(G78gat), .Z(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n319_), .A2(KEYINPUT11), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n320_), .A2(new_n321_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n318_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n315_), .A2(new_n326_), .A3(new_n317_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n297_), .B1(new_n330_), .B2(KEYINPUT17), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n297_), .A2(KEYINPUT17), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(KEYINPUT77), .A3(new_n329_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n331_), .A2(new_n334_), .A3(new_n332_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n293_), .A2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n339_), .A2(KEYINPUT78), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(KEYINPUT78), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n225_), .A2(new_n244_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n327_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n326_), .B1(new_n225_), .B2(new_n244_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G230gat), .A2(G233gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT64), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n326_), .A2(KEYINPUT12), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n245_), .A2(new_n250_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n348_), .B1(new_n342_), .B2(new_n327_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT12), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n344_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n349_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G120gat), .B(G148gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT5), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G176gat), .B(G204gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  NOR2_X1   g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n361_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT13), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n363_), .B(new_n364_), .C1(KEYINPUT69), .C2(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n367_));
  INV_X1    g166(.A(new_n364_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(new_n362_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n340_), .A2(new_n341_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT91), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G141gat), .A2(G148gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT89), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT89), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(G141gat), .A3(G148gat), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n375_), .B(new_n377_), .C1(G141gat), .C2(G148gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(KEYINPUT1), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT1), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n381_), .B1(G155gat), .B2(G162gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n379_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n383_), .B2(KEYINPUT90), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT90), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n385_), .A3(new_n379_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n378_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G155gat), .B(G162gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n389_));
  INV_X1    g188(.A(G141gat), .ZN(new_n390_));
  INV_X1    g189(.A(G148gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT2), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n375_), .A2(new_n377_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n388_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n373_), .B1(new_n387_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n388_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n397_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n400_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n382_), .A2(new_n385_), .A3(new_n379_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n385_), .B1(new_n382_), .B2(new_n379_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n404_), .A2(new_n405_), .A3(new_n380_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n403_), .B(KEYINPUT91), .C1(new_n406_), .C2(new_n378_), .ZN(new_n407_));
  INV_X1    g206(.A(G134gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G127gat), .ZN(new_n409_));
  INV_X1    g208(.A(G127gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G134gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G113gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(G120gat), .ZN(new_n414_));
  INV_X1    g213(.A(G120gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(G113gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n412_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G113gat), .B(G120gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n417_), .A2(new_n419_), .A3(KEYINPUT87), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT87), .B1(new_n417_), .B2(new_n419_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n399_), .A2(new_n407_), .A3(new_n422_), .A4(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G225gat), .A2(G233gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n399_), .A2(new_n407_), .A3(new_n422_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT98), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n387_), .A2(new_n398_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n417_), .A2(new_n419_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n429_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  NOR4_X1   g232(.A1(new_n387_), .A2(new_n431_), .A3(new_n398_), .A4(KEYINPUT98), .ZN(new_n434_));
  OAI211_X1 g233(.A(KEYINPUT4), .B(new_n428_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n427_), .A2(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n428_), .B(new_n425_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G1gat), .B(G29gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(G85gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT0), .B(G57gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n442_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n436_), .A2(new_n437_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G8gat), .B(G36gat), .Z(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G64gat), .B(G92gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n451_), .A2(KEYINPUT32), .ZN(new_n452_));
  AND2_X1   g251(.A1(KEYINPUT93), .A2(G204gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(KEYINPUT93), .A2(G204gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(G197gat), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(G197gat), .A2(G204gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT21), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G211gat), .B(G218gat), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n453_), .A2(new_n454_), .A3(G197gat), .ZN(new_n462_));
  INV_X1    g261(.A(G197gat), .ZN(new_n463_));
  INV_X1    g262(.A(G204gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT21), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n460_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT94), .B1(new_n458_), .B2(new_n459_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT94), .ZN(new_n469_));
  AOI211_X1 g268(.A(new_n469_), .B(KEYINPUT21), .C1(new_n455_), .C2(new_n457_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n467_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT95), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT93), .B(G204gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n456_), .B1(new_n474_), .B2(G197gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n469_), .B1(new_n475_), .B2(KEYINPUT21), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n458_), .A2(KEYINPUT94), .A3(new_n459_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(KEYINPUT95), .A3(new_n467_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n461_), .B1(new_n473_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G183gat), .A2(G190gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT23), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT23), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(G183gat), .A3(G190gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT24), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G169gat), .A2(G176gat), .ZN(new_n486_));
  AOI22_X1  g285(.A1(new_n482_), .A2(new_n484_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT96), .ZN(new_n488_));
  AND2_X1   g287(.A1(G169gat), .A2(G176gat), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n489_), .A2(new_n486_), .A3(new_n485_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT25), .B(G183gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT26), .B(G190gat), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT85), .B(G176gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT22), .B(G169gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n489_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n481_), .A2(new_n483_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n497_), .B(new_n498_), .C1(G183gat), .C2(G190gat), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n488_), .A2(new_n493_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT20), .B1(new_n480_), .B2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT82), .B(G190gat), .ZN(new_n502_));
  INV_X1    g301(.A(G183gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n496_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n482_), .A2(new_n484_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n486_), .A2(new_n485_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n487_), .A2(KEYINPUT84), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n490_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT81), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT80), .B(KEYINPUT25), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n515_), .B1(new_n516_), .B2(new_n503_), .ZN(new_n517_));
  INV_X1    g316(.A(G190gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT83), .B1(new_n518_), .B2(KEYINPUT26), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT26), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(G190gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n503_), .A2(KEYINPUT25), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n519_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n525_), .A2(KEYINPUT80), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(KEYINPUT80), .ZN(new_n527_));
  OAI211_X1 g326(.A(KEYINPUT81), .B(G183gat), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n502_), .A2(KEYINPUT26), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n517_), .A2(new_n524_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n507_), .B1(new_n514_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n461_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT95), .B1(new_n478_), .B2(new_n467_), .ZN(new_n533_));
  AOI211_X1 g332(.A(new_n472_), .B(new_n466_), .C1(new_n476_), .C2(new_n477_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n531_), .B(new_n532_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G226gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT19), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n501_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT20), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n480_), .B2(new_n500_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n490_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n487_), .A2(KEYINPUT84), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n530_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n506_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n540_), .B1(new_n542_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n452_), .B1(new_n539_), .B2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n538_), .B1(new_n501_), .B2(new_n536_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(new_n540_), .A3(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n446_), .B(new_n550_), .C1(new_n452_), .C2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n451_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n500_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n541_), .B1(new_n543_), .B2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n540_), .B1(new_n557_), .B2(new_n535_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n532_), .B(new_n500_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT20), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n473_), .A2(new_n479_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n531_), .B1(new_n561_), .B2(new_n532_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n560_), .A2(new_n562_), .A3(new_n538_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n555_), .B1(new_n558_), .B2(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n424_), .A2(new_n425_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT100), .B1(new_n565_), .B2(new_n435_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n428_), .B(new_n426_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n442_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n565_), .A2(new_n435_), .A3(KEYINPUT100), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n551_), .A2(new_n451_), .A3(new_n552_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n436_), .A2(new_n437_), .A3(KEYINPUT33), .A4(new_n444_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n564_), .A2(new_n571_), .A3(new_n572_), .A4(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT33), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n445_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT99), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n445_), .A2(new_n578_), .A3(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n554_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT29), .B1(new_n399_), .B2(new_n407_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT28), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n399_), .A2(new_n407_), .A3(KEYINPUT29), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G228gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT92), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n543_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT29), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n430_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n585_), .B1(new_n543_), .B2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n583_), .B1(new_n587_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n399_), .A2(new_n407_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n588_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT28), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT28), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n582_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(G228gat), .B(G233gat), .C1(new_n480_), .C2(new_n589_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n543_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G78gat), .B(G106gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G22gat), .B(G50gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  AND3_X1   g403(.A1(new_n592_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n592_), .B2(new_n601_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n581_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n572_), .A2(KEYINPUT27), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n538_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n557_), .A2(new_n540_), .A3(new_n535_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n451_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT27), .B1(new_n564_), .B2(new_n572_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n604_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n616_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n592_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n446_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n608_), .A2(new_n622_), .ZN(new_n623_));
  OR3_X1    g422(.A1(new_n420_), .A2(new_n421_), .A3(KEYINPUT31), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT31), .B1(new_n420_), .B2(new_n421_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n624_), .A2(KEYINPUT88), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT88), .B1(new_n624_), .B2(new_n625_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT86), .B(G43gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n546_), .A2(KEYINPUT30), .A3(new_n506_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT30), .B1(new_n546_), .B2(new_n506_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT30), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n547_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n546_), .A2(KEYINPUT30), .A3(new_n506_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n629_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G227gat), .A2(G233gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(G15gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(G71gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(G99gat), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n633_), .A2(new_n637_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n633_), .B2(new_n637_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n628_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n641_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n631_), .A2(new_n632_), .A3(new_n630_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n629_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n633_), .A2(new_n637_), .A3(new_n641_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n626_), .A3(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n644_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT27), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n551_), .A2(new_n451_), .A3(new_n552_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n451_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n654_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n555_), .B1(new_n539_), .B2(new_n549_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(KEYINPUT27), .A3(new_n572_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n443_), .A2(new_n445_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n651_), .A2(new_n661_), .A3(new_n620_), .A4(new_n619_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n653_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n644_), .A2(new_n443_), .A3(new_n650_), .A4(new_n445_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n664_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n665_), .A2(KEYINPUT101), .A3(new_n657_), .A4(new_n659_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n623_), .A2(new_n652_), .B1(new_n663_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n259_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n312_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(G229gat), .A2(G233gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT79), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n673_), .B(new_n259_), .C1(new_n308_), .C2(new_n311_), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT79), .B1(new_n312_), .B2(new_n668_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n670_), .B(new_n672_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n312_), .B1(new_n262_), .B2(new_n261_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n306_), .A2(new_n307_), .A3(new_n299_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n298_), .B1(new_n310_), .B2(new_n305_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n668_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n673_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n312_), .A2(KEYINPUT79), .A3(new_n668_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n677_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n676_), .B1(new_n683_), .B2(new_n672_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(G113gat), .B(G141gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(G169gat), .B(G197gat), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n685_), .B(new_n686_), .Z(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n687_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n676_), .B(new_n689_), .C1(new_n683_), .C2(new_n672_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n667_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n372_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n446_), .A2(new_n300_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT102), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n697_));
  INV_X1    g496(.A(new_n695_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n372_), .A2(new_n697_), .A3(new_n693_), .A4(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n696_), .A2(KEYINPUT38), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n288_), .A2(new_n289_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n607_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n655_), .A2(new_n656_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n445_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n705_), .A2(KEYINPUT33), .B1(new_n569_), .B2(new_n570_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n704_), .A2(new_n706_), .A3(new_n577_), .A4(new_n579_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n703_), .B1(new_n707_), .B2(new_n554_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n621_), .A2(new_n657_), .A3(new_n659_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n652_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n663_), .A2(new_n666_), .ZN(new_n711_));
  AOI211_X1 g510(.A(KEYINPUT103), .B(new_n702_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n581_), .A2(new_n607_), .B1(new_n615_), .B2(new_n621_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n711_), .B1(new_n714_), .B2(new_n651_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n713_), .B1(new_n715_), .B2(new_n701_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n712_), .A2(new_n716_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n371_), .A2(new_n692_), .A3(new_n338_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G1gat), .B1(new_n719_), .B2(new_n661_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n700_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT38), .B1(new_n696_), .B2(new_n699_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT104), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n722_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(new_n720_), .A4(new_n700_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1324gat));
  NAND4_X1  g526(.A1(new_n372_), .A2(new_n301_), .A3(new_n660_), .A4(new_n693_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n660_), .B(new_n718_), .C1(new_n712_), .C2(new_n716_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(G8gat), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n729_), .B2(G8gat), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(KEYINPUT39), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT39), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n729_), .A2(G8gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT105), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n737_), .B2(new_n731_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n728_), .B1(new_n734_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT40), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT40), .B(new_n728_), .C1(new_n734_), .C2(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1325gat));
  OR3_X1    g542(.A1(new_n694_), .A2(G15gat), .A3(new_n652_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G15gat), .B1(new_n719_), .B2(new_n652_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT41), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n746_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1326gat));
  OR3_X1    g548(.A1(new_n694_), .A2(G22gat), .A3(new_n607_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n717_), .A2(new_n703_), .A3(new_n718_), .ZN(new_n751_));
  XOR2_X1   g550(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n752_));
  AND3_X1   g551(.A1(new_n751_), .A2(G22gat), .A3(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n751_), .B2(G22gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(G1327gat));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n667_), .B2(new_n292_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n715_), .A2(new_n759_), .A3(new_n293_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n370_), .A2(new_n691_), .A3(new_n338_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT44), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n765_));
  AOI211_X1 g564(.A(new_n765_), .B(new_n762_), .C1(new_n758_), .C2(new_n760_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n446_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G29gat), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n702_), .A2(new_n338_), .ZN(new_n770_));
  NOR4_X1   g569(.A1(new_n667_), .A2(new_n692_), .A3(new_n371_), .A4(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n661_), .A2(G29gat), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT108), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n769_), .A2(new_n774_), .ZN(G1328gat));
  INV_X1    g574(.A(G36gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n771_), .A2(new_n776_), .A3(new_n660_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT45), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n767_), .B2(new_n660_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n667_), .A2(KEYINPUT43), .A3(new_n292_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n759_), .B1(new_n715_), .B2(new_n293_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n763_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n765_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n761_), .A2(KEYINPUT44), .A3(new_n763_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n784_), .A2(new_n779_), .A3(new_n660_), .A4(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(G36gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n778_), .B1(new_n780_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT46), .B(new_n778_), .C1(new_n780_), .C2(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1329gat));
  NAND2_X1  g591(.A1(new_n767_), .A2(new_n651_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(G43gat), .ZN(new_n794_));
  INV_X1    g593(.A(G43gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n771_), .A2(new_n795_), .A3(new_n651_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n794_), .A2(KEYINPUT47), .A3(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1330gat));
  AOI21_X1  g600(.A(G50gat), .B1(new_n771_), .B2(new_n703_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n703_), .A2(G50gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n767_), .B2(new_n803_), .ZN(G1331gat));
  INV_X1    g603(.A(new_n338_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n692_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(new_n370_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n717_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n717_), .A2(KEYINPUT111), .A3(new_n807_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n446_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G57gat), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n340_), .A2(new_n341_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n667_), .A2(new_n691_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n371_), .A3(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT110), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n661_), .A2(G57gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n813_), .B1(new_n817_), .B2(new_n818_), .ZN(G1332gat));
  NAND3_X1  g618(.A1(new_n810_), .A2(new_n660_), .A3(new_n811_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT48), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n820_), .A2(new_n821_), .A3(G64gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n820_), .B2(G64gat), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n615_), .A2(G64gat), .ZN(new_n824_));
  OAI22_X1  g623(.A1(new_n822_), .A2(new_n823_), .B1(new_n817_), .B2(new_n824_), .ZN(G1333gat));
  NAND3_X1  g624(.A1(new_n810_), .A2(new_n651_), .A3(new_n811_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n826_), .A2(G71gat), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n826_), .B2(G71gat), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n652_), .A2(G71gat), .ZN(new_n830_));
  OAI22_X1  g629(.A1(new_n828_), .A2(new_n829_), .B1(new_n817_), .B2(new_n830_), .ZN(G1334gat));
  NAND3_X1  g630(.A1(new_n810_), .A2(new_n703_), .A3(new_n811_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(G78gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(G78gat), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n607_), .A2(G78gat), .ZN(new_n836_));
  OAI22_X1  g635(.A1(new_n834_), .A2(new_n835_), .B1(new_n817_), .B2(new_n836_), .ZN(G1335gat));
  NOR3_X1   g636(.A1(new_n370_), .A2(new_n805_), .A3(new_n691_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n761_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G85gat), .B1(new_n840_), .B2(new_n661_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n770_), .A2(new_n370_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n815_), .A2(new_n842_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n661_), .A2(G85gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(G1336gat));
  OAI21_X1  g644(.A(G92gat), .B1(new_n840_), .B2(new_n615_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n615_), .A2(G92gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n843_), .B2(new_n847_), .ZN(G1337gat));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849_));
  INV_X1    g648(.A(new_n242_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n843_), .A2(new_n652_), .A3(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n761_), .A2(new_n651_), .A3(new_n838_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(G99gat), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n849_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT51), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n852_), .A2(G99gat), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n858_), .A2(KEYINPUT113), .A3(new_n851_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n855_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT113), .B1(new_n858_), .B2(new_n851_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n853_), .A2(new_n856_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n849_), .A4(KEYINPUT51), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n860_), .A2(new_n863_), .ZN(G1338gat));
  NAND4_X1  g663(.A1(new_n815_), .A2(new_n230_), .A3(new_n703_), .A4(new_n842_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n839_), .A2(new_n703_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(G106gat), .ZN(new_n868_));
  AOI211_X1 g667(.A(KEYINPUT52), .B(new_n230_), .C1(new_n839_), .C2(new_n703_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n865_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n865_), .B(new_n871_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1339gat));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n669_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT116), .B(new_n689_), .C1(new_n877_), .C2(new_n672_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n683_), .A2(new_n672_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n670_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n671_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT116), .B1(new_n882_), .B2(new_n689_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n688_), .B1(new_n880_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n688_), .B(KEYINPUT117), .C1(new_n880_), .C2(new_n883_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT55), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n356_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n352_), .A2(new_n343_), .A3(new_n355_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n348_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n352_), .A2(new_n353_), .A3(KEYINPUT55), .A4(new_n355_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n895_), .A3(new_n361_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n363_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n894_), .B2(new_n361_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n888_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n292_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n888_), .A2(new_n899_), .A3(KEYINPUT118), .A4(KEYINPUT58), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n888_), .A2(new_n899_), .A3(KEYINPUT58), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(new_n903_), .A3(new_n906_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n886_), .A2(new_n887_), .B1(new_n364_), .B2(new_n363_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n897_), .A2(new_n692_), .A3(new_n898_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n701_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  OAI211_X1 g711(.A(KEYINPUT57), .B(new_n701_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n907_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n338_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n806_), .A2(new_n371_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n292_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n338_), .A2(new_n691_), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n292_), .A2(new_n916_), .A3(new_n370_), .A4(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n918_), .A2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n703_), .B1(new_n915_), .B2(new_n923_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n660_), .A2(new_n661_), .A3(new_n652_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n876_), .B1(new_n926_), .B2(KEYINPUT119), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n924_), .A2(new_n928_), .A3(KEYINPUT59), .A4(new_n925_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n692_), .B1(new_n927_), .B2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n691_), .A2(new_n413_), .ZN(new_n931_));
  OAI22_X1  g730(.A1(new_n930_), .A2(new_n413_), .B1(new_n926_), .B2(new_n931_), .ZN(G1340gat));
  AOI21_X1  g731(.A(new_n370_), .B1(new_n927_), .B2(new_n929_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n415_), .B1(new_n370_), .B2(KEYINPUT60), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n415_), .A2(KEYINPUT60), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(KEYINPUT120), .B2(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(KEYINPUT120), .B2(new_n934_), .ZN(new_n937_));
  OAI22_X1  g736(.A1(new_n933_), .A2(new_n415_), .B1(new_n926_), .B2(new_n937_), .ZN(G1341gat));
  AOI21_X1  g737(.A(new_n338_), .B1(new_n927_), .B2(new_n929_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n805_), .A2(new_n410_), .ZN(new_n940_));
  OAI22_X1  g739(.A1(new_n939_), .A2(new_n410_), .B1(new_n926_), .B2(new_n940_), .ZN(G1342gat));
  AOI21_X1  g740(.A(new_n292_), .B1(new_n927_), .B2(new_n929_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n702_), .A2(new_n408_), .ZN(new_n943_));
  OAI22_X1  g742(.A1(new_n942_), .A2(new_n408_), .B1(new_n926_), .B2(new_n943_), .ZN(G1343gat));
  NAND2_X1  g743(.A1(new_n915_), .A2(new_n923_), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n660_), .A2(new_n607_), .A3(new_n661_), .A4(new_n651_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n692_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n390_), .ZN(G1344gat));
  NOR2_X1   g748(.A1(new_n947_), .A2(new_n370_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT121), .B(G148gat), .Z(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1345gat));
  OR3_X1    g751(.A1(new_n947_), .A2(KEYINPUT122), .A3(new_n338_), .ZN(new_n953_));
  OAI21_X1  g752(.A(KEYINPUT122), .B1(new_n947_), .B2(new_n338_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(KEYINPUT61), .B(G155gat), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n953_), .A2(new_n954_), .A3(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(new_n953_), .B2(new_n954_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1346gat));
  OR3_X1    g757(.A1(new_n947_), .A2(G162gat), .A3(new_n701_), .ZN(new_n959_));
  OAI21_X1  g758(.A(G162gat), .B1(new_n947_), .B2(new_n292_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(G1347gat));
  NOR2_X1   g760(.A1(new_n615_), .A2(new_n664_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(new_n691_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(KEYINPUT123), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n924_), .A2(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n965_), .A2(G169gat), .ZN(new_n966_));
  AND2_X1   g765(.A1(new_n966_), .A2(KEYINPUT62), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n966_), .A2(KEYINPUT62), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n945_), .A2(new_n660_), .A3(new_n665_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n691_), .A2(new_n495_), .ZN(new_n970_));
  OAI22_X1  g769(.A1(new_n967_), .A2(new_n968_), .B1(new_n969_), .B2(new_n970_), .ZN(G1348gat));
  OAI21_X1  g770(.A(new_n494_), .B1(new_n969_), .B2(new_n370_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n922_), .B1(new_n914_), .B2(new_n338_), .ZN(new_n973_));
  OAI21_X1  g772(.A(KEYINPUT124), .B1(new_n973_), .B2(new_n703_), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n975_));
  AND2_X1   g774(.A1(new_n912_), .A2(new_n913_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n805_), .B1(new_n976_), .B2(new_n907_), .ZN(new_n977_));
  OAI211_X1 g776(.A(new_n975_), .B(new_n607_), .C1(new_n977_), .C2(new_n922_), .ZN(new_n978_));
  AND2_X1   g777(.A1(new_n371_), .A2(G176gat), .ZN(new_n979_));
  NAND4_X1  g778(.A1(new_n974_), .A2(new_n978_), .A3(new_n962_), .A4(new_n979_), .ZN(new_n980_));
  AND2_X1   g779(.A1(new_n972_), .A2(new_n980_), .ZN(G1349gat));
  NAND2_X1  g780(.A1(new_n962_), .A2(new_n805_), .ZN(new_n982_));
  INV_X1    g781(.A(new_n982_), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n974_), .A2(new_n978_), .A3(new_n983_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n984_), .A2(new_n503_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n982_), .A2(new_n491_), .ZN(new_n986_));
  AOI21_X1  g785(.A(KEYINPUT125), .B1(new_n924_), .B2(new_n986_), .ZN(new_n987_));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n988_));
  INV_X1    g787(.A(new_n986_), .ZN(new_n989_));
  NOR4_X1   g788(.A1(new_n973_), .A2(new_n988_), .A3(new_n703_), .A4(new_n989_), .ZN(new_n990_));
  NOR2_X1   g789(.A1(new_n987_), .A2(new_n990_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n985_), .A2(new_n991_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n992_), .A2(KEYINPUT126), .ZN(new_n993_));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n994_));
  NAND3_X1  g793(.A1(new_n985_), .A2(new_n991_), .A3(new_n994_), .ZN(new_n995_));
  NAND2_X1  g794(.A1(new_n993_), .A2(new_n995_), .ZN(G1350gat));
  OAI21_X1  g795(.A(G190gat), .B1(new_n969_), .B2(new_n292_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n702_), .A2(new_n492_), .ZN(new_n998_));
  OAI21_X1  g797(.A(new_n997_), .B1(new_n969_), .B2(new_n998_), .ZN(G1351gat));
  NAND2_X1  g798(.A1(new_n621_), .A2(new_n652_), .ZN(new_n1000_));
  INV_X1    g799(.A(new_n1000_), .ZN(new_n1001_));
  NAND3_X1  g800(.A1(new_n945_), .A2(new_n660_), .A3(new_n1001_), .ZN(new_n1002_));
  NOR2_X1   g801(.A1(new_n1002_), .A2(new_n692_), .ZN(new_n1003_));
  XNOR2_X1  g802(.A(new_n1003_), .B(new_n463_), .ZN(G1352gat));
  NOR3_X1   g803(.A1(new_n1002_), .A2(new_n474_), .A3(new_n370_), .ZN(new_n1005_));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n1006_));
  AND2_X1   g805(.A1(new_n1005_), .A2(new_n1006_), .ZN(new_n1007_));
  NOR2_X1   g806(.A1(new_n1005_), .A2(new_n1006_), .ZN(new_n1008_));
  OAI21_X1  g807(.A(G204gat), .B1(new_n1002_), .B2(new_n370_), .ZN(new_n1009_));
  AOI21_X1  g808(.A(new_n1007_), .B1(new_n1008_), .B2(new_n1009_), .ZN(G1353gat));
  NOR2_X1   g809(.A1(new_n1002_), .A2(new_n338_), .ZN(new_n1011_));
  NOR3_X1   g810(.A1(new_n1011_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1012_));
  XOR2_X1   g811(.A(KEYINPUT63), .B(G211gat), .Z(new_n1013_));
  AOI21_X1  g812(.A(new_n1012_), .B1(new_n1011_), .B2(new_n1013_), .ZN(G1354gat));
  OAI21_X1  g813(.A(G218gat), .B1(new_n1002_), .B2(new_n292_), .ZN(new_n1015_));
  OR2_X1    g814(.A1(new_n701_), .A2(G218gat), .ZN(new_n1016_));
  OAI21_X1  g815(.A(new_n1015_), .B1(new_n1002_), .B2(new_n1016_), .ZN(G1355gat));
endmodule


