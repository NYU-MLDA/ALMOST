//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_;
  XOR2_X1   g000(.A(G155gat), .B(G162gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT85), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT85), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G141gat), .A3(G148gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n206_), .A2(new_n208_), .A3(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(KEYINPUT3), .ZN(new_n216_));
  OR3_X1    g015(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n218_), .A2(new_n219_), .A3(new_n202_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(new_n218_), .B2(new_n202_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n212_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI211_X1 g023(.A(KEYINPUT87), .B(new_n212_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OR3_X1    g025(.A1(new_n226_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n227_));
  INV_X1    g026(.A(G78gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT28), .B1(new_n226_), .B2(KEYINPUT29), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n228_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n232_));
  OAI21_X1  g031(.A(G106gat), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n232_), .ZN(new_n234_));
  INV_X1    g033(.A(G106gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n230_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n226_), .A2(KEYINPUT29), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT89), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G211gat), .B(G218gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(G197gat), .B(G204gat), .Z(new_n242_));
  OAI21_X1  g041(.A(new_n241_), .B1(new_n242_), .B2(KEYINPUT21), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(KEYINPUT21), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n238_), .A2(new_n239_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT90), .B(G233gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n248_), .A2(G228gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(KEYINPUT91), .Z(new_n250_));
  NAND4_X1  g049(.A1(new_n240_), .A2(new_n246_), .A3(new_n247_), .A4(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G22gat), .B(G50gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT88), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n222_), .A2(KEYINPUT92), .A3(KEYINPUT29), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n246_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT92), .B1(new_n222_), .B2(KEYINPUT29), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n249_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n254_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n237_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n251_), .A2(new_n258_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n253_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n264_), .A2(new_n233_), .A3(new_n236_), .A4(new_n259_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G169gat), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(KEYINPUT24), .A3(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(KEYINPUT25), .B(G183gat), .Z(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT26), .B(G190gat), .Z(new_n273_));
  OAI221_X1 g072(.A(new_n271_), .B1(KEYINPUT24), .B2(new_n269_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT23), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT22), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(KEYINPUT80), .ZN(new_n280_));
  OAI21_X1  g079(.A(G169gat), .B1(new_n280_), .B2(G176gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT81), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n282_), .B1(new_n275_), .B2(KEYINPUT23), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(new_n276_), .B2(new_n282_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285_));
  OAI221_X1 g084(.A(new_n281_), .B1(new_n269_), .B2(new_n280_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n278_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT82), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n278_), .A2(new_n286_), .A3(KEYINPUT82), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n245_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n270_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT22), .B(G169gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(new_n293_), .B2(new_n268_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT93), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(new_n277_), .B2(new_n285_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(new_n284_), .B2(new_n274_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n246_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n291_), .A2(KEYINPUT20), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT19), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n297_), .A2(new_n246_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n290_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT82), .B1(new_n278_), .B2(new_n286_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n246_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n301_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n303_), .A2(new_n306_), .A3(KEYINPUT20), .A4(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G8gat), .B(G36gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(G64gat), .B(G92gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n302_), .A2(new_n308_), .A3(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n299_), .A2(new_n301_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n303_), .A2(new_n306_), .A3(KEYINPUT20), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(new_n301_), .B2(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(KEYINPUT27), .B(new_n317_), .C1(new_n323_), .C2(new_n314_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n266_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT101), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT97), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT96), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n332_), .A2(G113gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(G113gat), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n333_), .A2(G120gat), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(G120gat), .B1(new_n333_), .B2(new_n334_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n218_), .A2(new_n202_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT86), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n218_), .A2(new_n219_), .A3(new_n202_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT87), .B1(new_n342_), .B2(new_n212_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n225_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n338_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n337_), .A3(new_n212_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n331_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n346_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(KEYINPUT96), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT4), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n337_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(KEYINPUT4), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n330_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n347_), .A2(new_n329_), .A3(new_n349_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G1gat), .B(G29gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G57gat), .B(G85gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  NOR3_X1   g159(.A1(new_n354_), .A2(new_n355_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n360_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT96), .B1(new_n351_), .B2(new_n348_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n349_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n329_), .B1(new_n366_), .B2(new_n352_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n355_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n362_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n327_), .B1(new_n361_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n360_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n368_), .A3(new_n362_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(KEYINPUT101), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT30), .B1(new_n304_), .B2(new_n305_), .ZN(new_n376_));
  INV_X1    g175(.A(G43gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n289_), .A2(new_n378_), .A3(new_n290_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n377_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G15gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G71gat), .B(G99gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n384_), .B(new_n385_), .Z(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n381_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n376_), .A2(new_n379_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G43gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n390_), .B2(new_n380_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n375_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT84), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n387_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n380_), .A3(new_n386_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(KEYINPUT83), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n337_), .B(KEYINPUT31), .Z(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n395_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n375_), .A3(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n393_), .A2(new_n396_), .A3(new_n397_), .A4(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n397_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n399_), .B1(new_n398_), .B2(new_n375_), .ZN(new_n403_));
  AOI211_X1 g202(.A(KEYINPUT83), .B(KEYINPUT84), .C1(new_n394_), .C2(new_n395_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n326_), .A2(new_n374_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n325_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n361_), .A2(new_n369_), .A3(new_n327_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT101), .B1(new_n371_), .B2(new_n372_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n406_), .B1(new_n411_), .B2(new_n266_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n364_), .A2(new_n329_), .A3(new_n365_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n360_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT99), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n330_), .B1(new_n366_), .B2(new_n352_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT99), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n417_), .A3(new_n360_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT100), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n415_), .A2(new_n416_), .A3(KEYINPUT100), .A4(new_n418_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT95), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n318_), .B(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n361_), .A2(KEYINPUT33), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n372_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .A4(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n262_), .A2(new_n265_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n314_), .A2(KEYINPUT32), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n302_), .A2(new_n308_), .A3(new_n431_), .ZN(new_n432_));
  OAI221_X1 g231(.A(new_n432_), .B1(new_n323_), .B2(new_n431_), .C1(new_n361_), .C2(new_n369_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT102), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n412_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n412_), .B2(new_n434_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n407_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G1gat), .B(G8gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT73), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G15gat), .ZN(new_n442_));
  INV_X1    g241(.A(G22gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G15gat), .A2(G22gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G1gat), .A2(G8gat), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n444_), .A2(new_n445_), .B1(KEYINPUT14), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n441_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT71), .B(G43gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G50gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(G29gat), .B(G36gat), .Z(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G50gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n449_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n451_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n452_), .A2(new_n456_), .A3(KEYINPUT15), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT15), .B1(new_n452_), .B2(new_n456_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n448_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT77), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G229gat), .A2(G233gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n452_), .A2(new_n456_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n448_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT77), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n448_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n460_), .A2(new_n461_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n441_), .A2(new_n447_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n441_), .A2(new_n447_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n452_), .A2(new_n456_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(new_n463_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT76), .B1(new_n473_), .B2(new_n461_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT76), .ZN(new_n475_));
  INV_X1    g274(.A(new_n461_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n475_), .B(new_n476_), .C1(new_n472_), .C2(new_n463_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n467_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G169gat), .B(G197gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT78), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(G113gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(G141gat), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n467_), .A2(new_n474_), .A3(new_n477_), .A4(new_n482_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT79), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT12), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT7), .ZN(new_n490_));
  INV_X1    g289(.A(G99gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n235_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n492_), .A2(new_n495_), .A3(new_n496_), .A4(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G85gat), .A2(G92gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n498_), .A2(KEYINPUT8), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT8), .B1(new_n498_), .B2(new_n502_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n495_), .A2(new_n496_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT9), .B1(new_n500_), .B2(new_n501_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT9), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT65), .B1(new_n499_), .B2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n506_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n500_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT64), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT10), .B(G99gat), .Z(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n513_), .B2(new_n235_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT10), .B(G99gat), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n515_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n510_), .B(new_n511_), .C1(new_n514_), .C2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n489_), .B1(new_n505_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G57gat), .ZN(new_n519_));
  INV_X1    g318(.A(G64gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT11), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G57gat), .A2(G64gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n525_));
  INV_X1    g324(.A(G71gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(G78gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n228_), .A2(G71gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n524_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n525_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n522_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n530_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(G57gat), .A2(G64gat), .ZN(new_n535_));
  NOR2_X1   g334(.A1(G57gat), .A2(G64gat), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n535_), .A2(new_n536_), .A3(KEYINPUT11), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G71gat), .B(G78gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT66), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n524_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n532_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT68), .B1(new_n534_), .B2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n533_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n539_), .A2(new_n540_), .A3(new_n532_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n518_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n505_), .A2(new_n517_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n545_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n551_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n489_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n518_), .A2(new_n542_), .A3(KEYINPUT69), .A4(new_n546_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n549_), .A2(new_n555_), .A3(new_n557_), .A4(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G120gat), .B(G148gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G204gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT5), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(new_n268_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n550_), .A2(new_n551_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n556_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT67), .B1(new_n565_), .B2(new_n554_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT67), .ZN(new_n567_));
  AOI211_X1 g366(.A(new_n567_), .B(new_n553_), .C1(new_n564_), .C2(new_n556_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n559_), .B(new_n563_), .C1(new_n566_), .C2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n556_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n554_), .B1(new_n572_), .B2(new_n552_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n567_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n565_), .A2(KEYINPUT67), .A3(new_n554_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n576_), .A2(KEYINPUT70), .A3(new_n559_), .A4(new_n563_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n559_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n563_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n582_), .A2(KEYINPUT13), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(KEYINPUT13), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n551_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n470_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT16), .B(G183gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G127gat), .B(G155gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT74), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n588_), .B(KEYINPUT68), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n595_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT15), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n462_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n452_), .A2(new_n456_), .A3(KEYINPUT15), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT72), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n550_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n605_), .B2(new_n550_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT34), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n471_), .A2(new_n517_), .A3(new_n505_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n610_), .A2(KEYINPUT35), .A3(new_n612_), .A4(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n609_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n612_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT35), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n615_), .A2(new_n618_), .A3(new_n613_), .A4(new_n607_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n616_), .A2(new_n617_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G190gat), .B(G218gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(G134gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(G162gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT36), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n614_), .A2(new_n622_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT36), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n614_), .B2(new_n622_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT37), .B1(new_n628_), .B2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n614_), .A2(new_n622_), .A3(new_n627_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT37), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n614_), .A2(new_n622_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n634_), .B(new_n635_), .C1(new_n636_), .C2(new_n631_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n585_), .A2(new_n601_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT75), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n488_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n438_), .B(new_n641_), .C1(new_n640_), .C2(new_n639_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT103), .ZN(new_n643_));
  INV_X1    g442(.A(G1gat), .ZN(new_n644_));
  INV_X1    g443(.A(new_n374_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT38), .ZN(new_n647_));
  INV_X1    g446(.A(new_n601_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n486_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n585_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n628_), .A2(new_n632_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n438_), .A2(new_n648_), .A3(new_n650_), .A4(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n374_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n647_), .A2(new_n653_), .ZN(G1324gat));
  OAI21_X1  g453(.A(G8gat), .B1(new_n652_), .B2(new_n408_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT39), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n408_), .A2(G8gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n643_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT104), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n656_), .A2(new_n661_), .A3(new_n658_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n660_), .A2(KEYINPUT40), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT40), .B1(new_n660_), .B2(new_n662_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1325gat));
  INV_X1    g464(.A(new_n406_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G15gat), .B1(new_n652_), .B2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT41), .Z(new_n668_));
  NAND3_X1  g467(.A1(new_n643_), .A2(new_n442_), .A3(new_n406_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1326gat));
  OAI21_X1  g469(.A(G22gat), .B1(new_n652_), .B2(new_n430_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT42), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n643_), .A2(new_n443_), .A3(new_n266_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1327gat));
  INV_X1    g473(.A(new_n407_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n429_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n325_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n666_), .B1(new_n677_), .B2(new_n430_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT102), .B1(new_n676_), .B2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n412_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n681_), .A2(new_n648_), .A3(new_n651_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n585_), .A2(new_n488_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(G29gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n686_), .A3(new_n645_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n638_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n681_), .A2(KEYINPUT43), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n438_), .B2(new_n638_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n601_), .B(new_n650_), .C1(new_n689_), .C2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n692_), .A2(new_n693_), .A3(KEYINPUT44), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n374_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n687_), .B1(new_n698_), .B2(new_n686_), .ZN(G1328gat));
  INV_X1    g498(.A(G36gat), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n325_), .A2(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n684_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n408_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n700_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n707_), .B(new_n704_), .C1(new_n705_), .C2(new_n700_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1329gat));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n692_), .A2(new_n693_), .A3(KEYINPUT44), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT44), .B1(new_n692_), .B2(new_n693_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n406_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G43gat), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n684_), .A2(G43gat), .A3(new_n666_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n712_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT47), .B(new_n717_), .C1(new_n715_), .C2(G43gat), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1330gat));
  NAND3_X1  g520(.A1(new_n685_), .A2(new_n453_), .A3(new_n266_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n430_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n453_), .ZN(G1331gat));
  NOR2_X1   g523(.A1(new_n487_), .A2(new_n601_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n438_), .A2(new_n585_), .A3(new_n651_), .A4(new_n725_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n726_), .A2(new_n519_), .A3(new_n374_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT107), .Z(new_n728_));
  INV_X1    g527(.A(new_n585_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n486_), .ZN(new_n730_));
  AND4_X1   g529(.A1(new_n648_), .A2(new_n438_), .A3(new_n688_), .A4(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G57gat), .B1(new_n731_), .B2(new_n645_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n728_), .A2(new_n732_), .ZN(G1332gat));
  OAI21_X1  g532(.A(G64gat), .B1(new_n726_), .B2(new_n408_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n520_), .A3(new_n325_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT108), .ZN(G1333gat));
  OAI21_X1  g537(.A(G71gat), .B1(new_n726_), .B2(new_n666_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT109), .Z(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT49), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n731_), .A2(new_n526_), .A3(new_n406_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1334gat));
  OAI21_X1  g542(.A(G78gat), .B1(new_n726_), .B2(new_n430_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT50), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n731_), .A2(new_n228_), .A3(new_n266_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1335gat));
  AND2_X1   g546(.A1(new_n682_), .A2(new_n730_), .ZN(new_n748_));
  INV_X1    g547(.A(G85gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n645_), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT43), .B1(new_n681_), .B2(new_n688_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n438_), .A2(new_n690_), .A3(new_n638_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n648_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n730_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n754_), .A2(KEYINPUT110), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(KEYINPUT110), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n374_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n750_), .B1(new_n757_), .B2(new_n749_), .ZN(G1336gat));
  INV_X1    g557(.A(G92gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n748_), .A2(new_n759_), .A3(new_n325_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n408_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n759_), .ZN(G1337gat));
  NOR2_X1   g561(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n763_));
  OAI21_X1  g562(.A(G99gat), .B1(new_n754_), .B2(new_n666_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n748_), .A2(new_n513_), .A3(new_n406_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n766_), .B(new_n767_), .Z(G1338gat));
  NAND3_X1  g567(.A1(new_n748_), .A2(new_n235_), .A3(new_n266_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n753_), .A2(new_n266_), .A3(new_n730_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(G106gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G106gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g574(.A1(new_n460_), .A2(new_n476_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n776_), .B(new_n483_), .C1(new_n476_), .C2(new_n473_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n485_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n582_), .A2(new_n779_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n571_), .A2(new_n577_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n549_), .A2(new_n558_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n782_), .A2(KEYINPUT55), .A3(new_n555_), .A4(new_n557_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n549_), .A2(new_n564_), .A3(new_n557_), .A4(new_n558_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n554_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n559_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n783_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT112), .B1(new_n788_), .B2(new_n580_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n781_), .B1(new_n789_), .B2(KEYINPUT56), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT112), .B(new_n791_), .C1(new_n788_), .C2(new_n580_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n780_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n651_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n788_), .A2(new_n580_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n778_), .B1(new_n798_), .B2(KEYINPUT56), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n788_), .A2(new_n791_), .A3(new_n580_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n799_), .A2(KEYINPUT58), .A3(new_n578_), .A4(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n638_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(new_n578_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n804_), .B1(new_n806_), .B2(new_n799_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n797_), .B1(new_n802_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n796_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n793_), .A2(KEYINPUT57), .A3(new_n651_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n559_), .B(KEYINPUT55), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n563_), .B1(new_n811_), .B2(new_n785_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n779_), .B1(new_n812_), .B2(new_n791_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n803_), .B1(new_n813_), .B2(new_n805_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(new_n801_), .A3(KEYINPUT114), .A4(new_n638_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n810_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT115), .B1(new_n809_), .B2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n810_), .A2(new_n815_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n796_), .A4(new_n808_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n601_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n639_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT54), .B1(new_n822_), .B2(new_n487_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n638_), .A2(KEYINPUT54), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n729_), .A2(new_n725_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n821_), .A2(KEYINPUT116), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT116), .B1(new_n821_), .B2(new_n826_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n326_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n829_), .A2(new_n374_), .A3(new_n666_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n827_), .A2(new_n828_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(new_n486_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n802_), .A2(new_n807_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n795_), .B2(new_n794_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT118), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n810_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n835_), .A2(KEYINPUT118), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n601_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n826_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n830_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n832_), .B2(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n821_), .A2(new_n826_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n821_), .A2(KEYINPUT116), .A3(new_n826_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n830_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(KEYINPUT117), .A3(KEYINPUT59), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n843_), .B1(new_n845_), .B2(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n852_), .A2(G113gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n833_), .B1(new_n853_), .B2(new_n487_), .ZN(G1340gat));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855_));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n852_), .B2(new_n585_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT60), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n729_), .B2(KEYINPUT60), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n832_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n855_), .B1(new_n857_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n851_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT117), .B1(new_n850_), .B2(KEYINPUT59), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n585_), .B(new_n842_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G120gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT119), .A3(new_n861_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n863_), .A2(new_n868_), .ZN(G1341gat));
  AOI21_X1  g668(.A(G127gat), .B1(new_n832_), .B2(new_n648_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n852_), .A2(G127gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n648_), .ZN(G1342gat));
  INV_X1    g671(.A(new_n651_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G134gat), .B1(new_n832_), .B2(new_n873_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n852_), .A2(new_n638_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g675(.A1(new_n827_), .A2(new_n828_), .A3(new_n430_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n374_), .A2(new_n325_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n877_), .A2(new_n878_), .A3(new_n666_), .A4(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n848_), .A2(new_n266_), .A3(new_n666_), .A4(new_n849_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n879_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT120), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n486_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n585_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT122), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT121), .B(G148gat), .Z(new_n889_));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n884_), .A2(new_n890_), .A3(new_n585_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n888_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n889_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n884_), .B2(new_n585_), .ZN(new_n894_));
  AOI211_X1 g693(.A(KEYINPUT122), .B(new_n729_), .C1(new_n880_), .C2(new_n883_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n892_), .A2(new_n896_), .ZN(G1345gat));
  NAND2_X1  g696(.A1(new_n884_), .A2(new_n648_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT123), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT61), .B(G155gat), .Z(new_n900_));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n884_), .A2(new_n901_), .A3(new_n648_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n899_), .A2(new_n900_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n900_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n901_), .B1(new_n884_), .B2(new_n648_), .ZN(new_n905_));
  AOI211_X1 g704(.A(KEYINPUT123), .B(new_n601_), .C1(new_n880_), .C2(new_n883_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n907_), .ZN(G1346gat));
  AOI21_X1  g707(.A(G162gat), .B1(new_n884_), .B2(new_n873_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n688_), .B1(new_n880_), .B2(new_n883_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(G162gat), .B2(new_n910_), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n645_), .A2(new_n408_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n913_), .A2(new_n266_), .A3(new_n666_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n840_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n649_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G169gat), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n920_), .A2(KEYINPUT62), .A3(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n916_), .A2(new_n293_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n918_), .A2(new_n919_), .A3(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n922_), .A2(new_n923_), .A3(new_n925_), .ZN(G1348gat));
  INV_X1    g725(.A(new_n915_), .ZN(new_n927_));
  AOI21_X1  g726(.A(G176gat), .B1(new_n927_), .B2(new_n585_), .ZN(new_n928_));
  AND4_X1   g727(.A1(G176gat), .A2(new_n848_), .A3(new_n849_), .A4(new_n914_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n585_), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n648_), .A2(new_n272_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n848_), .A2(new_n648_), .A3(new_n849_), .A4(new_n914_), .ZN(new_n933_));
  INV_X1    g732(.A(G183gat), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n927_), .A2(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n915_), .B2(new_n688_), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n651_), .A2(new_n273_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n915_), .B2(new_n937_), .ZN(G1351gat));
  NAND4_X1  g737(.A1(new_n877_), .A2(KEYINPUT125), .A3(new_n666_), .A4(new_n912_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n940_), .B1(new_n881_), .B2(new_n913_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n649_), .B1(new_n939_), .B2(new_n941_), .ZN(new_n942_));
  AND3_X1   g741(.A1(new_n942_), .A2(KEYINPUT126), .A3(G197gat), .ZN(new_n943_));
  AOI21_X1  g742(.A(KEYINPUT126), .B1(new_n942_), .B2(G197gat), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n942_), .A2(G197gat), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(G1352gat));
  NAND2_X1  g745(.A1(new_n939_), .A2(new_n941_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n585_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  NAND2_X1  g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  AND4_X1   g750(.A1(new_n648_), .A2(new_n947_), .A3(new_n950_), .A4(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n950_), .B1(new_n947_), .B2(new_n648_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1354gat));
  AOI21_X1  g753(.A(G218gat), .B1(new_n947_), .B2(new_n873_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n638_), .A2(G218gat), .ZN(new_n956_));
  XOR2_X1   g755(.A(new_n956_), .B(KEYINPUT127), .Z(new_n957_));
  AOI21_X1  g756(.A(new_n955_), .B1(new_n947_), .B2(new_n957_), .ZN(G1355gat));
endmodule


