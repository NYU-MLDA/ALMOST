// Benchmark "c6288" written by ABC on Wed Jul  6 02:18:53 2022

module c6288 ( 
    G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat,
    G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat  );
  input  G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat;
  output G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat;
  wire new_n65_, new_n66_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n86_, new_n87_, new_n88_,
    new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_,
    new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n144_, new_n145_,
    new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_,
    new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_,
    new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_,
    new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_,
    new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_,
    new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_,
    new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_,
    new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_,
    new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_,
    new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_,
    new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_,
    new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_,
    new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_,
    new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_,
    new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_,
    new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_,
    new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_,
    new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_,
    new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_,
    new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_,
    new_n2260_, new_n2261_, new_n2262_, new_n2264_, new_n2265_, new_n2266_,
    new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_,
    new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_,
    new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_,
    new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_,
    new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_,
    new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_,
    new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_,
    new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_,
    new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_,
    new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_,
    new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_,
    new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_,
    new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_,
    new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_,
    new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_,
    new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_,
    new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_,
    new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_,
    new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_,
    new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2718_, new_n2719_, new_n2720_,
    new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_,
    new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_,
    new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_,
    new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_,
    new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_,
    new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_,
    new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_,
    new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_,
    new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_,
    new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_,
    new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_,
    new_n2972_, new_n2973_, new_n2974_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2988_, new_n2989_, new_n2990_;
  INV_X1    g0000(.A(G1gat), .ZN(new_n65_));
  INV_X1    g0001(.A(G273gat), .ZN(new_n66_));
  NOR2_X1   g0002(.A1(new_n65_), .A2(new_n66_), .ZN(G545gat));
  INV_X1    g0003(.A(G18gat), .ZN(new_n68_));
  NOR2_X1   g0004(.A1(new_n68_), .A2(new_n66_), .ZN(new_n69_));
  INV_X1    g0005(.A(G290gat), .ZN(new_n70_));
  NOR2_X1   g0006(.A1(new_n65_), .A2(new_n70_), .ZN(new_n71_));
  NAND2_X1  g0007(.A1(new_n69_), .A2(new_n71_), .ZN(new_n72_));
  INV_X1    g0008(.A(new_n72_), .ZN(new_n73_));
  NOR2_X1   g0009(.A1(new_n69_), .A2(new_n71_), .ZN(new_n74_));
  NOR2_X1   g0010(.A1(new_n73_), .A2(new_n74_), .ZN(G1581gat));
  INV_X1    g0011(.A(G35gat), .ZN(new_n76_));
  OAI22_X1  g0012(.A1(new_n68_), .A2(new_n70_), .B1(new_n76_), .B2(new_n66_), .ZN(new_n77_));
  NAND4_X1  g0013(.A1(G18gat), .A2(G35gat), .A3(G273gat), .A4(G290gat), .ZN(new_n78_));
  NAND2_X1  g0014(.A1(new_n77_), .A2(new_n78_), .ZN(new_n79_));
  NOR2_X1   g0015(.A1(new_n73_), .A2(new_n79_), .ZN(new_n80_));
  INV_X1    g0016(.A(new_n80_), .ZN(new_n81_));
  NAND2_X1  g0017(.A1(new_n73_), .A2(new_n79_), .ZN(new_n82_));
  NAND2_X1  g0018(.A1(new_n81_), .A2(new_n82_), .ZN(new_n83_));
  NAND2_X1  g0019(.A1(G1gat), .A2(G307gat), .ZN(new_n84_));
  XNOR2_X1  g0020(.A(new_n83_), .B(new_n84_), .ZN(G1901gat));
  INV_X1    g0021(.A(G52gat), .ZN(new_n86_));
  OAI22_X1  g0022(.A1(new_n76_), .A2(new_n70_), .B1(new_n86_), .B2(new_n66_), .ZN(new_n87_));
  NAND4_X1  g0023(.A1(G35gat), .A2(G52gat), .A3(G273gat), .A4(G290gat), .ZN(new_n88_));
  NAND3_X1  g0024(.A1(new_n87_), .A2(new_n78_), .A3(new_n88_), .ZN(new_n89_));
  INV_X1    g0025(.A(new_n89_), .ZN(new_n90_));
  AOI21_X1  g0026(.A(new_n78_), .B1(new_n87_), .B2(new_n88_), .ZN(new_n91_));
  NOR2_X1   g0027(.A1(new_n90_), .A2(new_n91_), .ZN(new_n92_));
  NAND2_X1  g0028(.A1(G18gat), .A2(G307gat), .ZN(new_n93_));
  NOR2_X1   g0029(.A1(new_n92_), .A2(new_n93_), .ZN(new_n94_));
  INV_X1    g0030(.A(new_n94_), .ZN(new_n95_));
  NAND2_X1  g0031(.A1(new_n92_), .A2(new_n93_), .ZN(new_n96_));
  AOI22_X1  g0032(.A1(new_n81_), .A2(new_n82_), .B1(G1gat), .B2(G307gat), .ZN(new_n97_));
  NAND2_X1  g0033(.A1(new_n79_), .A2(new_n72_), .ZN(new_n98_));
  INV_X1    g0034(.A(new_n98_), .ZN(new_n99_));
  OAI211_X1 g0035(.A(new_n95_), .B(new_n96_), .C1(new_n97_), .C2(new_n99_), .ZN(new_n100_));
  NAND2_X1  g0036(.A1(new_n83_), .A2(new_n84_), .ZN(new_n101_));
  INV_X1    g0037(.A(new_n96_), .ZN(new_n102_));
  OAI211_X1 g0038(.A(new_n101_), .B(new_n98_), .C1(new_n102_), .C2(new_n94_), .ZN(new_n103_));
  NAND2_X1  g0039(.A1(new_n100_), .A2(new_n103_), .ZN(new_n104_));
  NAND2_X1  g0040(.A1(G1gat), .A2(G324gat), .ZN(new_n105_));
  XNOR2_X1  g0041(.A(new_n104_), .B(new_n105_), .ZN(G2223gat));
  NAND2_X1  g0042(.A1(G1gat), .A2(G341gat), .ZN(new_n107_));
  NAND2_X1  g0043(.A1(new_n104_), .A2(new_n105_), .ZN(new_n108_));
  OAI21_X1  g0044(.A(new_n93_), .B1(new_n90_), .B2(new_n91_), .ZN(new_n109_));
  NAND2_X1  g0045(.A1(new_n87_), .A2(new_n88_), .ZN(new_n110_));
  NAND2_X1  g0046(.A1(new_n110_), .A2(new_n78_), .ZN(new_n111_));
  NAND2_X1  g0047(.A1(new_n109_), .A2(new_n111_), .ZN(new_n112_));
  INV_X1    g0048(.A(G69gat), .ZN(new_n113_));
  OAI22_X1  g0049(.A1(new_n86_), .A2(new_n70_), .B1(new_n113_), .B2(new_n66_), .ZN(new_n114_));
  NAND4_X1  g0050(.A1(G52gat), .A2(G69gat), .A3(G273gat), .A4(G290gat), .ZN(new_n115_));
  NAND3_X1  g0051(.A1(new_n114_), .A2(new_n88_), .A3(new_n115_), .ZN(new_n116_));
  INV_X1    g0052(.A(new_n116_), .ZN(new_n117_));
  AOI21_X1  g0053(.A(new_n88_), .B1(new_n114_), .B2(new_n115_), .ZN(new_n118_));
  OAI211_X1 g0054(.A(G35gat), .B(G307gat), .C1(new_n117_), .C2(new_n118_), .ZN(new_n119_));
  NAND2_X1  g0055(.A1(new_n114_), .A2(new_n115_), .ZN(new_n120_));
  INV_X1    g0056(.A(new_n88_), .ZN(new_n121_));
  NAND2_X1  g0057(.A1(new_n120_), .A2(new_n121_), .ZN(new_n122_));
  NAND2_X1  g0058(.A1(G35gat), .A2(G307gat), .ZN(new_n123_));
  NAND3_X1  g0059(.A1(new_n122_), .A2(new_n116_), .A3(new_n123_), .ZN(new_n124_));
  NAND3_X1  g0060(.A1(new_n112_), .A2(new_n119_), .A3(new_n124_), .ZN(new_n125_));
  AND3_X1   g0061(.A1(new_n122_), .A2(new_n116_), .A3(new_n123_), .ZN(new_n126_));
  AOI21_X1  g0062(.A(new_n123_), .B1(new_n122_), .B2(new_n116_), .ZN(new_n127_));
  OAI211_X1 g0063(.A(new_n109_), .B(new_n111_), .C1(new_n126_), .C2(new_n127_), .ZN(new_n128_));
  NAND2_X1  g0064(.A1(new_n125_), .A2(new_n128_), .ZN(new_n129_));
  INV_X1    g0065(.A(G324gat), .ZN(new_n130_));
  NOR2_X1   g0066(.A1(new_n68_), .A2(new_n130_), .ZN(new_n131_));
  NAND2_X1  g0067(.A1(new_n129_), .A2(new_n131_), .ZN(new_n132_));
  OAI211_X1 g0068(.A(new_n125_), .B(new_n128_), .C1(new_n68_), .C2(new_n130_), .ZN(new_n133_));
  NAND2_X1  g0069(.A1(new_n132_), .A2(new_n133_), .ZN(new_n134_));
  AOI22_X1  g0070(.A1(new_n96_), .A2(new_n95_), .B1(new_n98_), .B2(new_n101_), .ZN(new_n135_));
  INV_X1    g0071(.A(new_n135_), .ZN(new_n136_));
  NAND3_X1  g0072(.A1(new_n108_), .A2(new_n134_), .A3(new_n136_), .ZN(new_n137_));
  AOI22_X1  g0073(.A1(new_n100_), .A2(new_n103_), .B1(G1gat), .B2(G324gat), .ZN(new_n138_));
  OAI211_X1 g0074(.A(new_n132_), .B(new_n133_), .C1(new_n138_), .C2(new_n135_), .ZN(new_n139_));
  AOI21_X1  g0075(.A(new_n107_), .B1(new_n137_), .B2(new_n139_), .ZN(new_n140_));
  AOI22_X1  g0076(.A1(new_n139_), .A2(new_n137_), .B1(G1gat), .B2(G341gat), .ZN(new_n141_));
  INV_X1    g0077(.A(new_n141_), .ZN(new_n142_));
  AOI21_X1  g0078(.A(new_n140_), .B1(new_n107_), .B2(new_n142_), .ZN(G2548gat));
  OAI21_X1  g0079(.A(new_n123_), .B1(new_n117_), .B2(new_n118_), .ZN(new_n144_));
  NAND2_X1  g0080(.A1(new_n120_), .A2(new_n88_), .ZN(new_n145_));
  INV_X1    g0081(.A(G86gat), .ZN(new_n146_));
  OAI22_X1  g0082(.A1(new_n113_), .A2(new_n70_), .B1(new_n146_), .B2(new_n66_), .ZN(new_n147_));
  NAND4_X1  g0083(.A1(G69gat), .A2(G86gat), .A3(G273gat), .A4(G290gat), .ZN(new_n148_));
  NAND3_X1  g0084(.A1(new_n147_), .A2(new_n115_), .A3(new_n148_), .ZN(new_n149_));
  INV_X1    g0085(.A(new_n149_), .ZN(new_n150_));
  AOI21_X1  g0086(.A(new_n115_), .B1(new_n147_), .B2(new_n148_), .ZN(new_n151_));
  NAND2_X1  g0087(.A1(G52gat), .A2(G307gat), .ZN(new_n152_));
  INV_X1    g0088(.A(new_n152_), .ZN(new_n153_));
  NOR3_X1   g0089(.A1(new_n150_), .A2(new_n151_), .A3(new_n153_), .ZN(new_n154_));
  NAND2_X1  g0090(.A1(new_n147_), .A2(new_n148_), .ZN(new_n155_));
  INV_X1    g0091(.A(new_n115_), .ZN(new_n156_));
  NAND2_X1  g0092(.A1(new_n155_), .A2(new_n156_), .ZN(new_n157_));
  AOI21_X1  g0093(.A(new_n152_), .B1(new_n157_), .B2(new_n149_), .ZN(new_n158_));
  OAI211_X1 g0094(.A(new_n144_), .B(new_n145_), .C1(new_n154_), .C2(new_n158_), .ZN(new_n159_));
  OAI21_X1  g0095(.A(new_n153_), .B1(new_n150_), .B2(new_n151_), .ZN(new_n160_));
  NAND3_X1  g0096(.A1(new_n157_), .A2(new_n149_), .A3(new_n152_), .ZN(new_n161_));
  AOI22_X1  g0097(.A1(new_n122_), .A2(new_n116_), .B1(G35gat), .B2(G307gat), .ZN(new_n162_));
  INV_X1    g0098(.A(new_n145_), .ZN(new_n163_));
  OAI211_X1 g0099(.A(new_n160_), .B(new_n161_), .C1(new_n162_), .C2(new_n163_), .ZN(new_n164_));
  NAND2_X1  g0100(.A1(new_n159_), .A2(new_n164_), .ZN(new_n165_));
  NOR2_X1   g0101(.A1(new_n76_), .A2(new_n130_), .ZN(new_n166_));
  NAND2_X1  g0102(.A1(new_n165_), .A2(new_n166_), .ZN(new_n167_));
  OAI211_X1 g0103(.A(new_n159_), .B(new_n164_), .C1(new_n76_), .C2(new_n130_), .ZN(new_n168_));
  NAND2_X1  g0104(.A1(new_n167_), .A2(new_n168_), .ZN(new_n169_));
  AOI21_X1  g0105(.A(new_n131_), .B1(new_n125_), .B2(new_n128_), .ZN(new_n170_));
  NAND2_X1  g0106(.A1(new_n119_), .A2(new_n124_), .ZN(new_n171_));
  NAND2_X1  g0107(.A1(new_n171_), .A2(new_n112_), .ZN(new_n172_));
  INV_X1    g0108(.A(new_n172_), .ZN(new_n173_));
  NOR2_X1   g0109(.A1(new_n170_), .A2(new_n173_), .ZN(new_n174_));
  NAND2_X1  g0110(.A1(new_n169_), .A2(new_n174_), .ZN(new_n175_));
  OAI211_X1 g0111(.A(new_n167_), .B(new_n168_), .C1(new_n170_), .C2(new_n173_), .ZN(new_n176_));
  NAND2_X1  g0112(.A1(new_n175_), .A2(new_n176_), .ZN(new_n177_));
  INV_X1    g0113(.A(G341gat), .ZN(new_n178_));
  NOR2_X1   g0114(.A1(new_n68_), .A2(new_n178_), .ZN(new_n179_));
  NAND2_X1  g0115(.A1(new_n177_), .A2(new_n179_), .ZN(new_n180_));
  INV_X1    g0116(.A(new_n179_), .ZN(new_n181_));
  NAND3_X1  g0117(.A1(new_n175_), .A2(new_n176_), .A3(new_n181_), .ZN(new_n182_));
  NAND2_X1  g0118(.A1(new_n180_), .A2(new_n182_), .ZN(new_n183_));
  NAND2_X1  g0119(.A1(new_n108_), .A2(new_n136_), .ZN(new_n184_));
  NAND2_X1  g0120(.A1(new_n184_), .A2(new_n134_), .ZN(new_n185_));
  NAND3_X1  g0121(.A1(new_n142_), .A2(new_n183_), .A3(new_n185_), .ZN(new_n186_));
  INV_X1    g0122(.A(new_n185_), .ZN(new_n187_));
  OAI211_X1 g0123(.A(new_n180_), .B(new_n182_), .C1(new_n141_), .C2(new_n187_), .ZN(new_n188_));
  NAND2_X1  g0124(.A1(new_n186_), .A2(new_n188_), .ZN(new_n189_));
  INV_X1    g0125(.A(G358gat), .ZN(new_n190_));
  NOR2_X1   g0126(.A1(new_n65_), .A2(new_n190_), .ZN(new_n191_));
  XOR2_X1   g0127(.A(new_n189_), .B(new_n191_), .Z(G2877gat));
  AOI21_X1  g0128(.A(new_n191_), .B1(new_n186_), .B2(new_n188_), .ZN(new_n193_));
  INV_X1    g0129(.A(new_n193_), .ZN(new_n194_));
  NAND2_X1  g0130(.A1(new_n177_), .A2(new_n181_), .ZN(new_n195_));
  INV_X1    g0131(.A(new_n174_), .ZN(new_n196_));
  NAND2_X1  g0132(.A1(new_n196_), .A2(new_n169_), .ZN(new_n197_));
  AOI21_X1  g0133(.A(new_n166_), .B1(new_n159_), .B2(new_n164_), .ZN(new_n198_));
  INV_X1    g0134(.A(new_n198_), .ZN(new_n199_));
  AOI22_X1  g0135(.A1(new_n145_), .A2(new_n144_), .B1(new_n160_), .B2(new_n161_), .ZN(new_n200_));
  INV_X1    g0136(.A(new_n200_), .ZN(new_n201_));
  NAND2_X1  g0137(.A1(new_n155_), .A2(new_n115_), .ZN(new_n202_));
  OAI21_X1  g0138(.A(new_n152_), .B1(new_n150_), .B2(new_n151_), .ZN(new_n203_));
  NAND2_X1  g0139(.A1(G69gat), .A2(G307gat), .ZN(new_n204_));
  INV_X1    g0140(.A(G103gat), .ZN(new_n205_));
  OAI22_X1  g0141(.A1(new_n146_), .A2(new_n70_), .B1(new_n205_), .B2(new_n66_), .ZN(new_n206_));
  NAND4_X1  g0142(.A1(G86gat), .A2(G103gat), .A3(G273gat), .A4(G290gat), .ZN(new_n207_));
  AOI21_X1  g0143(.A(new_n148_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g0144(.A(new_n208_), .ZN(new_n209_));
  NAND3_X1  g0145(.A1(new_n206_), .A2(new_n148_), .A3(new_n207_), .ZN(new_n210_));
  AOI21_X1  g0146(.A(new_n204_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g0147(.A(new_n210_), .ZN(new_n212_));
  INV_X1    g0148(.A(new_n204_), .ZN(new_n213_));
  NOR3_X1   g0149(.A1(new_n212_), .A2(new_n208_), .A3(new_n213_), .ZN(new_n214_));
  OAI211_X1 g0150(.A(new_n202_), .B(new_n203_), .C1(new_n211_), .C2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g0151(.A(new_n213_), .B1(new_n212_), .B2(new_n208_), .ZN(new_n216_));
  NAND3_X1  g0152(.A1(new_n209_), .A2(new_n210_), .A3(new_n204_), .ZN(new_n217_));
  AOI21_X1  g0153(.A(new_n153_), .B1(new_n157_), .B2(new_n149_), .ZN(new_n218_));
  INV_X1    g0154(.A(new_n202_), .ZN(new_n219_));
  OAI211_X1 g0155(.A(new_n216_), .B(new_n217_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g0156(.A1(new_n86_), .A2(new_n130_), .ZN(new_n221_));
  INV_X1    g0157(.A(new_n221_), .ZN(new_n222_));
  NAND3_X1  g0158(.A1(new_n215_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g0159(.A(new_n223_), .ZN(new_n224_));
  AOI21_X1  g0160(.A(new_n222_), .B1(new_n215_), .B2(new_n220_), .ZN(new_n225_));
  OAI211_X1 g0161(.A(new_n199_), .B(new_n201_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g0162(.A1(new_n215_), .A2(new_n220_), .ZN(new_n227_));
  NAND2_X1  g0163(.A1(new_n227_), .A2(new_n221_), .ZN(new_n228_));
  OAI211_X1 g0164(.A(new_n228_), .B(new_n223_), .C1(new_n198_), .C2(new_n200_), .ZN(new_n229_));
  NOR2_X1   g0165(.A1(new_n76_), .A2(new_n178_), .ZN(new_n230_));
  INV_X1    g0166(.A(new_n230_), .ZN(new_n231_));
  AND3_X1   g0167(.A1(new_n226_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g0168(.A(new_n231_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n233_));
  OAI211_X1 g0169(.A(new_n195_), .B(new_n197_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g0170(.A1(new_n226_), .A2(new_n229_), .ZN(new_n235_));
  NAND2_X1  g0171(.A1(new_n235_), .A2(new_n230_), .ZN(new_n236_));
  NAND3_X1  g0172(.A1(new_n226_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n237_));
  AOI21_X1  g0173(.A(new_n179_), .B1(new_n175_), .B2(new_n176_), .ZN(new_n238_));
  INV_X1    g0174(.A(new_n197_), .ZN(new_n239_));
  OAI211_X1 g0175(.A(new_n236_), .B(new_n237_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g0176(.A1(new_n234_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g0177(.A1(new_n68_), .A2(new_n190_), .ZN(new_n242_));
  NAND2_X1  g0178(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g0179(.A(new_n242_), .ZN(new_n244_));
  NAND3_X1  g0180(.A1(new_n234_), .A2(new_n240_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g0181(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g0182(.A1(new_n142_), .A2(new_n185_), .ZN(new_n247_));
  NAND2_X1  g0183(.A1(new_n247_), .A2(new_n183_), .ZN(new_n248_));
  NAND3_X1  g0184(.A1(new_n194_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g0185(.A(new_n248_), .ZN(new_n250_));
  OAI211_X1 g0186(.A(new_n243_), .B(new_n245_), .C1(new_n250_), .C2(new_n193_), .ZN(new_n251_));
  NAND2_X1  g0187(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g0188(.A(G375gat), .ZN(new_n253_));
  NOR2_X1   g0189(.A1(new_n65_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g0190(.A(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g0191(.A(new_n252_), .B(new_n255_), .ZN(G3211gat));
  NAND2_X1  g0192(.A1(new_n252_), .A2(new_n255_), .ZN(new_n257_));
  NAND2_X1  g0193(.A1(new_n194_), .A2(new_n248_), .ZN(new_n258_));
  NAND2_X1  g0194(.A1(new_n258_), .A2(new_n246_), .ZN(new_n259_));
  NAND2_X1  g0195(.A1(new_n241_), .A2(new_n244_), .ZN(new_n260_));
  NOR2_X1   g0196(.A1(new_n232_), .A2(new_n233_), .ZN(new_n261_));
  NOR2_X1   g0197(.A1(new_n238_), .A2(new_n239_), .ZN(new_n262_));
  NOR2_X1   g0198(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g0199(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g0200(.A1(new_n235_), .A2(new_n231_), .ZN(new_n265_));
  NOR2_X1   g0201(.A1(new_n224_), .A2(new_n225_), .ZN(new_n266_));
  NOR2_X1   g0202(.A1(new_n198_), .A2(new_n200_), .ZN(new_n267_));
  NOR2_X1   g0203(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g0204(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g0205(.A1(new_n227_), .A2(new_n222_), .ZN(new_n270_));
  AOI22_X1  g0206(.A1(new_n216_), .A2(new_n217_), .B1(new_n203_), .B2(new_n202_), .ZN(new_n271_));
  INV_X1    g0207(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g0208(.A1(new_n206_), .A2(new_n207_), .ZN(new_n273_));
  NAND2_X1  g0209(.A1(new_n273_), .A2(new_n148_), .ZN(new_n274_));
  OAI21_X1  g0210(.A(new_n204_), .B1(new_n212_), .B2(new_n208_), .ZN(new_n275_));
  INV_X1    g0211(.A(G120gat), .ZN(new_n276_));
  OAI22_X1  g0212(.A1(new_n205_), .A2(new_n70_), .B1(new_n276_), .B2(new_n66_), .ZN(new_n277_));
  NAND4_X1  g0213(.A1(G103gat), .A2(G120gat), .A3(G273gat), .A4(G290gat), .ZN(new_n278_));
  NAND3_X1  g0214(.A1(new_n277_), .A2(new_n207_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g0215(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g0216(.A(new_n207_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n281_));
  NAND2_X1  g0217(.A1(G86gat), .A2(G307gat), .ZN(new_n282_));
  INV_X1    g0218(.A(new_n282_), .ZN(new_n283_));
  NOR3_X1   g0219(.A1(new_n280_), .A2(new_n281_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g0220(.A1(new_n277_), .A2(new_n278_), .ZN(new_n285_));
  INV_X1    g0221(.A(new_n207_), .ZN(new_n286_));
  NAND2_X1  g0222(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g0223(.A(new_n282_), .B1(new_n287_), .B2(new_n279_), .ZN(new_n288_));
  OAI211_X1 g0224(.A(new_n274_), .B(new_n275_), .C1(new_n284_), .C2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g0225(.A(new_n283_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n290_));
  NAND3_X1  g0226(.A1(new_n287_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n291_));
  AOI21_X1  g0227(.A(new_n213_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n292_));
  INV_X1    g0228(.A(new_n274_), .ZN(new_n293_));
  OAI211_X1 g0229(.A(new_n290_), .B(new_n291_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g0230(.A1(new_n113_), .A2(new_n130_), .ZN(new_n295_));
  INV_X1    g0231(.A(new_n295_), .ZN(new_n296_));
  NAND3_X1  g0232(.A1(new_n289_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g0233(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g0234(.A(new_n296_), .B1(new_n289_), .B2(new_n294_), .ZN(new_n299_));
  OAI211_X1 g0235(.A(new_n270_), .B(new_n272_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g0236(.A1(new_n289_), .A2(new_n294_), .ZN(new_n301_));
  NAND2_X1  g0237(.A1(new_n301_), .A2(new_n295_), .ZN(new_n302_));
  AOI21_X1  g0238(.A(new_n221_), .B1(new_n215_), .B2(new_n220_), .ZN(new_n303_));
  OAI211_X1 g0239(.A(new_n302_), .B(new_n297_), .C1(new_n271_), .C2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g0240(.A1(new_n86_), .A2(new_n178_), .ZN(new_n305_));
  INV_X1    g0241(.A(new_n305_), .ZN(new_n306_));
  NAND3_X1  g0242(.A1(new_n300_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g0243(.A(new_n307_), .ZN(new_n308_));
  AOI21_X1  g0244(.A(new_n306_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n309_));
  OAI211_X1 g0245(.A(new_n265_), .B(new_n269_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g0246(.A1(new_n300_), .A2(new_n304_), .ZN(new_n311_));
  NAND2_X1  g0247(.A1(new_n311_), .A2(new_n305_), .ZN(new_n312_));
  AOI21_X1  g0248(.A(new_n230_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n313_));
  OAI211_X1 g0249(.A(new_n312_), .B(new_n307_), .C1(new_n268_), .C2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g0250(.A1(new_n76_), .A2(new_n190_), .ZN(new_n315_));
  INV_X1    g0251(.A(new_n315_), .ZN(new_n316_));
  AND3_X1   g0252(.A1(new_n310_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g0253(.A(new_n316_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n318_));
  OAI211_X1 g0254(.A(new_n260_), .B(new_n264_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g0255(.A1(new_n310_), .A2(new_n314_), .ZN(new_n320_));
  NAND2_X1  g0256(.A1(new_n320_), .A2(new_n315_), .ZN(new_n321_));
  NAND3_X1  g0257(.A1(new_n310_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n322_));
  AOI21_X1  g0258(.A(new_n242_), .B1(new_n234_), .B2(new_n240_), .ZN(new_n323_));
  OAI211_X1 g0259(.A(new_n321_), .B(new_n322_), .C1(new_n323_), .C2(new_n263_), .ZN(new_n324_));
  NOR2_X1   g0260(.A1(new_n68_), .A2(new_n253_), .ZN(new_n325_));
  INV_X1    g0261(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g0262(.A1(new_n319_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g0263(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g0264(.A(new_n326_), .B1(new_n319_), .B2(new_n324_), .ZN(new_n329_));
  OAI211_X1 g0265(.A(new_n257_), .B(new_n259_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n330_));
  INV_X1    g0266(.A(new_n329_), .ZN(new_n331_));
  AOI21_X1  g0267(.A(new_n254_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n332_));
  INV_X1    g0268(.A(new_n259_), .ZN(new_n333_));
  OAI211_X1 g0269(.A(new_n331_), .B(new_n327_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g0270(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g0271(.A(G392gat), .ZN(new_n336_));
  NOR2_X1   g0272(.A1(new_n65_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g0273(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g0274(.A(new_n335_), .B(new_n338_), .ZN(G3552gat));
  NAND2_X1  g0275(.A1(new_n335_), .A2(new_n338_), .ZN(new_n340_));
  NOR2_X1   g0276(.A1(new_n332_), .A2(new_n333_), .ZN(new_n341_));
  NOR2_X1   g0277(.A1(new_n328_), .A2(new_n329_), .ZN(new_n342_));
  NOR2_X1   g0278(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g0279(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g0280(.A1(new_n319_), .A2(new_n324_), .ZN(new_n345_));
  NAND2_X1  g0281(.A1(new_n345_), .A2(new_n326_), .ZN(new_n346_));
  NOR2_X1   g0282(.A1(new_n317_), .A2(new_n318_), .ZN(new_n347_));
  NOR2_X1   g0283(.A1(new_n323_), .A2(new_n263_), .ZN(new_n348_));
  NOR2_X1   g0284(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g0285(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g0286(.A1(new_n320_), .A2(new_n316_), .ZN(new_n351_));
  NOR2_X1   g0287(.A1(new_n308_), .A2(new_n309_), .ZN(new_n352_));
  NOR2_X1   g0288(.A1(new_n313_), .A2(new_n268_), .ZN(new_n353_));
  NOR2_X1   g0289(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g0290(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g0291(.A1(new_n311_), .A2(new_n306_), .ZN(new_n356_));
  NOR2_X1   g0292(.A1(new_n298_), .A2(new_n299_), .ZN(new_n357_));
  NOR2_X1   g0293(.A1(new_n303_), .A2(new_n271_), .ZN(new_n358_));
  NOR2_X1   g0294(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g0295(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g0296(.A1(new_n301_), .A2(new_n296_), .ZN(new_n361_));
  AOI22_X1  g0297(.A1(new_n274_), .A2(new_n275_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n362_));
  INV_X1    g0298(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g0299(.A1(new_n146_), .A2(new_n130_), .ZN(new_n364_));
  INV_X1    g0300(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g0301(.A1(G103gat), .A2(G307gat), .ZN(new_n366_));
  AOI22_X1  g0302(.A1(G120gat), .A2(G290gat), .B1(G137gat), .B2(G273gat), .ZN(new_n367_));
  INV_X1    g0303(.A(new_n367_), .ZN(new_n368_));
  NAND4_X1  g0304(.A1(G120gat), .A2(G137gat), .A3(G273gat), .A4(G290gat), .ZN(new_n369_));
  NAND3_X1  g0305(.A1(new_n368_), .A2(new_n278_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g0306(.A(new_n278_), .ZN(new_n371_));
  INV_X1    g0307(.A(new_n369_), .ZN(new_n372_));
  OAI21_X1  g0308(.A(new_n371_), .B1(new_n372_), .B2(new_n367_), .ZN(new_n373_));
  AOI21_X1  g0309(.A(new_n366_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g0310(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g0311(.A1(new_n370_), .A2(new_n373_), .A3(new_n366_), .ZN(new_n376_));
  AOI21_X1  g0312(.A(new_n283_), .B1(new_n287_), .B2(new_n279_), .ZN(new_n377_));
  NAND2_X1  g0313(.A1(new_n285_), .A2(new_n207_), .ZN(new_n378_));
  INV_X1    g0314(.A(new_n378_), .ZN(new_n379_));
  OAI211_X1 g0315(.A(new_n375_), .B(new_n376_), .C1(new_n377_), .C2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g0316(.A(new_n282_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n381_));
  INV_X1    g0317(.A(new_n376_), .ZN(new_n382_));
  OAI211_X1 g0318(.A(new_n381_), .B(new_n378_), .C1(new_n382_), .C2(new_n374_), .ZN(new_n383_));
  AOI21_X1  g0319(.A(new_n365_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n384_));
  AND3_X1   g0320(.A1(new_n380_), .A2(new_n383_), .A3(new_n365_), .ZN(new_n385_));
  OAI211_X1 g0321(.A(new_n361_), .B(new_n363_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g0322(.A1(new_n380_), .A2(new_n383_), .ZN(new_n387_));
  NAND2_X1  g0323(.A1(new_n387_), .A2(new_n364_), .ZN(new_n388_));
  NAND3_X1  g0324(.A1(new_n380_), .A2(new_n383_), .A3(new_n365_), .ZN(new_n389_));
  AOI21_X1  g0325(.A(new_n295_), .B1(new_n289_), .B2(new_n294_), .ZN(new_n390_));
  OAI211_X1 g0326(.A(new_n388_), .B(new_n389_), .C1(new_n390_), .C2(new_n362_), .ZN(new_n391_));
  NOR2_X1   g0327(.A1(new_n113_), .A2(new_n178_), .ZN(new_n392_));
  INV_X1    g0328(.A(new_n392_), .ZN(new_n393_));
  NAND3_X1  g0329(.A1(new_n386_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g0330(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g0331(.A(new_n393_), .B1(new_n386_), .B2(new_n391_), .ZN(new_n396_));
  OAI211_X1 g0332(.A(new_n356_), .B(new_n360_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g0333(.A1(new_n386_), .A2(new_n391_), .ZN(new_n398_));
  NAND2_X1  g0334(.A1(new_n398_), .A2(new_n392_), .ZN(new_n399_));
  AOI21_X1  g0335(.A(new_n305_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n400_));
  OAI211_X1 g0336(.A(new_n399_), .B(new_n394_), .C1(new_n400_), .C2(new_n359_), .ZN(new_n401_));
  NOR2_X1   g0337(.A1(new_n86_), .A2(new_n190_), .ZN(new_n402_));
  INV_X1    g0338(.A(new_n402_), .ZN(new_n403_));
  NAND3_X1  g0339(.A1(new_n397_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g0340(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g0341(.A(new_n403_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n406_));
  OAI211_X1 g0342(.A(new_n351_), .B(new_n355_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g0343(.A1(new_n397_), .A2(new_n401_), .ZN(new_n408_));
  NAND2_X1  g0344(.A1(new_n408_), .A2(new_n402_), .ZN(new_n409_));
  AOI21_X1  g0345(.A(new_n315_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n410_));
  OAI211_X1 g0346(.A(new_n409_), .B(new_n404_), .C1(new_n410_), .C2(new_n354_), .ZN(new_n411_));
  NOR2_X1   g0347(.A1(new_n76_), .A2(new_n253_), .ZN(new_n412_));
  INV_X1    g0348(.A(new_n412_), .ZN(new_n413_));
  AND3_X1   g0349(.A1(new_n407_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g0350(.A(new_n413_), .B1(new_n407_), .B2(new_n411_), .ZN(new_n415_));
  OAI211_X1 g0351(.A(new_n346_), .B(new_n350_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g0352(.A1(new_n407_), .A2(new_n411_), .ZN(new_n417_));
  NAND2_X1  g0353(.A1(new_n417_), .A2(new_n412_), .ZN(new_n418_));
  NAND3_X1  g0354(.A1(new_n407_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n419_));
  AOI21_X1  g0355(.A(new_n325_), .B1(new_n319_), .B2(new_n324_), .ZN(new_n420_));
  OAI211_X1 g0356(.A(new_n418_), .B(new_n419_), .C1(new_n420_), .C2(new_n349_), .ZN(new_n421_));
  NOR2_X1   g0357(.A1(new_n68_), .A2(new_n336_), .ZN(new_n422_));
  INV_X1    g0358(.A(new_n422_), .ZN(new_n423_));
  NAND3_X1  g0359(.A1(new_n416_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g0360(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g0361(.A(new_n423_), .B1(new_n416_), .B2(new_n421_), .ZN(new_n426_));
  OAI211_X1 g0362(.A(new_n340_), .B(new_n344_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  INV_X1    g0363(.A(new_n426_), .ZN(new_n428_));
  AOI21_X1  g0364(.A(new_n337_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n429_));
  OAI211_X1 g0365(.A(new_n428_), .B(new_n424_), .C1(new_n429_), .C2(new_n343_), .ZN(new_n430_));
  NAND2_X1  g0366(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g0367(.A(G409gat), .ZN(new_n432_));
  NOR2_X1   g0368(.A1(new_n65_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g0369(.A(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g0370(.A(new_n431_), .B(new_n434_), .ZN(G3895gat));
  NAND2_X1  g0371(.A1(new_n431_), .A2(new_n434_), .ZN(new_n436_));
  NOR2_X1   g0372(.A1(new_n429_), .A2(new_n343_), .ZN(new_n437_));
  NOR2_X1   g0373(.A1(new_n425_), .A2(new_n426_), .ZN(new_n438_));
  NOR2_X1   g0374(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g0375(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g0376(.A1(new_n416_), .A2(new_n421_), .ZN(new_n441_));
  NAND2_X1  g0377(.A1(new_n441_), .A2(new_n423_), .ZN(new_n442_));
  NOR2_X1   g0378(.A1(new_n414_), .A2(new_n415_), .ZN(new_n443_));
  NOR2_X1   g0379(.A1(new_n420_), .A2(new_n349_), .ZN(new_n444_));
  NOR2_X1   g0380(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g0381(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g0382(.A1(new_n417_), .A2(new_n413_), .ZN(new_n447_));
  NOR2_X1   g0383(.A1(new_n405_), .A2(new_n406_), .ZN(new_n448_));
  NOR2_X1   g0384(.A1(new_n410_), .A2(new_n354_), .ZN(new_n449_));
  NOR2_X1   g0385(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g0386(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g0387(.A1(new_n408_), .A2(new_n403_), .ZN(new_n452_));
  NOR2_X1   g0388(.A1(new_n395_), .A2(new_n396_), .ZN(new_n453_));
  NOR2_X1   g0389(.A1(new_n400_), .A2(new_n359_), .ZN(new_n454_));
  NOR2_X1   g0390(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g0391(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g0392(.A1(new_n398_), .A2(new_n393_), .ZN(new_n457_));
  NOR2_X1   g0393(.A1(new_n390_), .A2(new_n362_), .ZN(new_n458_));
  NOR2_X1   g0394(.A1(new_n385_), .A2(new_n384_), .ZN(new_n459_));
  NOR2_X1   g0395(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g0396(.A(new_n460_), .ZN(new_n461_));
  NOR2_X1   g0397(.A1(new_n146_), .A2(new_n178_), .ZN(new_n462_));
  INV_X1    g0398(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g0399(.A1(new_n387_), .A2(new_n365_), .ZN(new_n464_));
  AOI22_X1  g0400(.A1(new_n378_), .A2(new_n381_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n465_));
  INV_X1    g0401(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g0402(.A1(G120gat), .A2(G307gat), .ZN(new_n467_));
  AOI22_X1  g0403(.A1(G137gat), .A2(G290gat), .B1(G154gat), .B2(G273gat), .ZN(new_n468_));
  INV_X1    g0404(.A(new_n468_), .ZN(new_n469_));
  NAND4_X1  g0405(.A1(G137gat), .A2(G154gat), .A3(G273gat), .A4(G290gat), .ZN(new_n470_));
  NAND3_X1  g0406(.A1(new_n469_), .A2(new_n369_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g0407(.A(new_n470_), .ZN(new_n472_));
  OAI21_X1  g0408(.A(new_n372_), .B1(new_n472_), .B2(new_n468_), .ZN(new_n473_));
  AOI21_X1  g0409(.A(new_n467_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g0410(.A(new_n474_), .ZN(new_n475_));
  NAND3_X1  g0411(.A1(new_n471_), .A2(new_n473_), .A3(new_n467_), .ZN(new_n476_));
  AOI21_X1  g0412(.A(new_n371_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n477_));
  AOI22_X1  g0413(.A1(new_n370_), .A2(new_n373_), .B1(G103gat), .B2(G307gat), .ZN(new_n478_));
  OAI211_X1 g0414(.A(new_n475_), .B(new_n476_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  NOR3_X1   g0415(.A1(new_n371_), .A2(new_n372_), .A3(new_n367_), .ZN(new_n480_));
  AOI21_X1  g0416(.A(new_n278_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n481_));
  OAI21_X1  g0417(.A(new_n366_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g0418(.A(new_n477_), .ZN(new_n483_));
  INV_X1    g0419(.A(new_n476_), .ZN(new_n484_));
  OAI211_X1 g0420(.A(new_n482_), .B(new_n483_), .C1(new_n484_), .C2(new_n474_), .ZN(new_n485_));
  NOR2_X1   g0421(.A1(new_n205_), .A2(new_n130_), .ZN(new_n486_));
  INV_X1    g0422(.A(new_n486_), .ZN(new_n487_));
  AND3_X1   g0423(.A1(new_n479_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g0424(.A(new_n487_), .B1(new_n479_), .B2(new_n485_), .ZN(new_n489_));
  OAI211_X1 g0425(.A(new_n464_), .B(new_n466_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g0426(.A1(new_n479_), .A2(new_n485_), .ZN(new_n491_));
  NAND2_X1  g0427(.A1(new_n491_), .A2(new_n486_), .ZN(new_n492_));
  NAND3_X1  g0428(.A1(new_n479_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n493_));
  AOI21_X1  g0429(.A(new_n364_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n494_));
  OAI211_X1 g0430(.A(new_n492_), .B(new_n493_), .C1(new_n494_), .C2(new_n465_), .ZN(new_n495_));
  AOI21_X1  g0431(.A(new_n463_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n496_));
  AND3_X1   g0432(.A1(new_n490_), .A2(new_n495_), .A3(new_n463_), .ZN(new_n497_));
  OAI211_X1 g0433(.A(new_n457_), .B(new_n461_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g0434(.A1(new_n490_), .A2(new_n495_), .ZN(new_n499_));
  NAND2_X1  g0435(.A1(new_n499_), .A2(new_n462_), .ZN(new_n500_));
  NAND3_X1  g0436(.A1(new_n490_), .A2(new_n495_), .A3(new_n463_), .ZN(new_n501_));
  AOI21_X1  g0437(.A(new_n392_), .B1(new_n386_), .B2(new_n391_), .ZN(new_n502_));
  OAI211_X1 g0438(.A(new_n500_), .B(new_n501_), .C1(new_n502_), .C2(new_n460_), .ZN(new_n503_));
  NOR2_X1   g0439(.A1(new_n113_), .A2(new_n190_), .ZN(new_n504_));
  INV_X1    g0440(.A(new_n504_), .ZN(new_n505_));
  NAND3_X1  g0441(.A1(new_n498_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g0442(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g0443(.A(new_n505_), .B1(new_n498_), .B2(new_n503_), .ZN(new_n508_));
  OAI211_X1 g0444(.A(new_n452_), .B(new_n456_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g0445(.A1(new_n498_), .A2(new_n503_), .ZN(new_n510_));
  NAND2_X1  g0446(.A1(new_n510_), .A2(new_n504_), .ZN(new_n511_));
  AOI21_X1  g0447(.A(new_n402_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n512_));
  OAI211_X1 g0448(.A(new_n511_), .B(new_n506_), .C1(new_n512_), .C2(new_n455_), .ZN(new_n513_));
  NOR2_X1   g0449(.A1(new_n86_), .A2(new_n253_), .ZN(new_n514_));
  INV_X1    g0450(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g0451(.A1(new_n509_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g0452(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g0453(.A(new_n515_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n518_));
  OAI211_X1 g0454(.A(new_n447_), .B(new_n451_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g0455(.A1(new_n509_), .A2(new_n513_), .ZN(new_n520_));
  NAND2_X1  g0456(.A1(new_n520_), .A2(new_n514_), .ZN(new_n521_));
  AOI21_X1  g0457(.A(new_n412_), .B1(new_n407_), .B2(new_n411_), .ZN(new_n522_));
  OAI211_X1 g0458(.A(new_n521_), .B(new_n516_), .C1(new_n522_), .C2(new_n450_), .ZN(new_n523_));
  NOR2_X1   g0459(.A1(new_n76_), .A2(new_n336_), .ZN(new_n524_));
  INV_X1    g0460(.A(new_n524_), .ZN(new_n525_));
  AND3_X1   g0461(.A1(new_n519_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g0462(.A(new_n525_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n527_));
  OAI211_X1 g0463(.A(new_n442_), .B(new_n446_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g0464(.A1(new_n519_), .A2(new_n523_), .ZN(new_n529_));
  NAND2_X1  g0465(.A1(new_n529_), .A2(new_n524_), .ZN(new_n530_));
  NAND3_X1  g0466(.A1(new_n519_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n531_));
  AOI21_X1  g0467(.A(new_n422_), .B1(new_n416_), .B2(new_n421_), .ZN(new_n532_));
  OAI211_X1 g0468(.A(new_n530_), .B(new_n531_), .C1(new_n532_), .C2(new_n445_), .ZN(new_n533_));
  NOR2_X1   g0469(.A1(new_n68_), .A2(new_n432_), .ZN(new_n534_));
  INV_X1    g0470(.A(new_n534_), .ZN(new_n535_));
  NAND3_X1  g0471(.A1(new_n528_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g0472(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g0473(.A(new_n535_), .B1(new_n528_), .B2(new_n533_), .ZN(new_n538_));
  OAI211_X1 g0474(.A(new_n436_), .B(new_n440_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n539_));
  INV_X1    g0475(.A(new_n538_), .ZN(new_n540_));
  AOI21_X1  g0476(.A(new_n433_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n541_));
  OAI211_X1 g0477(.A(new_n540_), .B(new_n536_), .C1(new_n541_), .C2(new_n439_), .ZN(new_n542_));
  NAND2_X1  g0478(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g0479(.A(G426gat), .ZN(new_n544_));
  NOR2_X1   g0480(.A1(new_n65_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g0481(.A(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g0482(.A(new_n543_), .B(new_n546_), .ZN(G4241gat));
  NAND2_X1  g0483(.A1(new_n543_), .A2(new_n546_), .ZN(new_n548_));
  NOR2_X1   g0484(.A1(new_n541_), .A2(new_n439_), .ZN(new_n549_));
  NOR2_X1   g0485(.A1(new_n537_), .A2(new_n538_), .ZN(new_n550_));
  NOR2_X1   g0486(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g0487(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g0488(.A1(new_n528_), .A2(new_n533_), .ZN(new_n553_));
  NAND2_X1  g0489(.A1(new_n553_), .A2(new_n535_), .ZN(new_n554_));
  NOR2_X1   g0490(.A1(new_n526_), .A2(new_n527_), .ZN(new_n555_));
  NOR2_X1   g0491(.A1(new_n532_), .A2(new_n445_), .ZN(new_n556_));
  NOR2_X1   g0492(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g0493(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g0494(.A1(new_n529_), .A2(new_n525_), .ZN(new_n559_));
  NOR2_X1   g0495(.A1(new_n517_), .A2(new_n518_), .ZN(new_n560_));
  NOR2_X1   g0496(.A1(new_n522_), .A2(new_n450_), .ZN(new_n561_));
  NOR2_X1   g0497(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g0498(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g0499(.A1(new_n520_), .A2(new_n515_), .ZN(new_n564_));
  NOR2_X1   g0500(.A1(new_n507_), .A2(new_n508_), .ZN(new_n565_));
  NOR2_X1   g0501(.A1(new_n512_), .A2(new_n455_), .ZN(new_n566_));
  NOR2_X1   g0502(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g0503(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g0504(.A1(new_n510_), .A2(new_n505_), .ZN(new_n569_));
  NOR2_X1   g0505(.A1(new_n497_), .A2(new_n496_), .ZN(new_n570_));
  NOR2_X1   g0506(.A1(new_n502_), .A2(new_n460_), .ZN(new_n571_));
  NOR2_X1   g0507(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g0508(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g0509(.A1(new_n146_), .A2(new_n190_), .ZN(new_n574_));
  INV_X1    g0510(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g0511(.A1(new_n499_), .A2(new_n463_), .ZN(new_n576_));
  NOR2_X1   g0512(.A1(new_n488_), .A2(new_n489_), .ZN(new_n577_));
  NOR2_X1   g0513(.A1(new_n494_), .A2(new_n465_), .ZN(new_n578_));
  NOR2_X1   g0514(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g0515(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g0516(.A1(new_n491_), .A2(new_n487_), .ZN(new_n581_));
  AOI22_X1  g0517(.A1(new_n475_), .A2(new_n476_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n582_));
  INV_X1    g0518(.A(new_n582_), .ZN(new_n583_));
  AOI22_X1  g0519(.A1(G154gat), .A2(G290gat), .B1(G171gat), .B2(G273gat), .ZN(new_n584_));
  INV_X1    g0520(.A(new_n584_), .ZN(new_n585_));
  NAND4_X1  g0521(.A1(G154gat), .A2(G171gat), .A3(G273gat), .A4(G290gat), .ZN(new_n586_));
  NAND3_X1  g0522(.A1(new_n585_), .A2(new_n470_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g0523(.A(new_n586_), .ZN(new_n588_));
  OAI21_X1  g0524(.A(new_n472_), .B1(new_n588_), .B2(new_n584_), .ZN(new_n589_));
  NAND2_X1  g0525(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g0526(.A1(G137gat), .A2(G307gat), .ZN(new_n591_));
  INV_X1    g0527(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g0528(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g0529(.A1(new_n587_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n594_));
  AOI22_X1  g0530(.A1(new_n471_), .A2(new_n473_), .B1(G120gat), .B2(G307gat), .ZN(new_n595_));
  AOI21_X1  g0531(.A(new_n372_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n596_));
  OAI211_X1 g0532(.A(new_n593_), .B(new_n594_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n597_));
  NOR3_X1   g0533(.A1(new_n372_), .A2(new_n472_), .A3(new_n468_), .ZN(new_n598_));
  AOI21_X1  g0534(.A(new_n369_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n599_));
  OAI21_X1  g0535(.A(new_n467_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g0536(.A(new_n596_), .ZN(new_n601_));
  AND3_X1   g0537(.A1(new_n587_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n602_));
  AOI21_X1  g0538(.A(new_n591_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n603_));
  OAI211_X1 g0539(.A(new_n600_), .B(new_n601_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g0540(.A1(new_n276_), .A2(new_n130_), .ZN(new_n605_));
  INV_X1    g0541(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g0542(.A1(new_n597_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g0543(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g0544(.A(new_n606_), .B1(new_n597_), .B2(new_n604_), .ZN(new_n609_));
  OAI211_X1 g0545(.A(new_n581_), .B(new_n583_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g0546(.A1(new_n597_), .A2(new_n604_), .ZN(new_n611_));
  NAND2_X1  g0547(.A1(new_n611_), .A2(new_n605_), .ZN(new_n612_));
  AOI21_X1  g0548(.A(new_n486_), .B1(new_n479_), .B2(new_n485_), .ZN(new_n613_));
  OAI211_X1 g0549(.A(new_n612_), .B(new_n607_), .C1(new_n613_), .C2(new_n582_), .ZN(new_n614_));
  NOR2_X1   g0550(.A1(new_n205_), .A2(new_n178_), .ZN(new_n615_));
  INV_X1    g0551(.A(new_n615_), .ZN(new_n616_));
  AND3_X1   g0552(.A1(new_n610_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g0553(.A(new_n616_), .B1(new_n610_), .B2(new_n614_), .ZN(new_n618_));
  OAI211_X1 g0554(.A(new_n576_), .B(new_n580_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g0555(.A1(new_n610_), .A2(new_n614_), .ZN(new_n620_));
  NAND2_X1  g0556(.A1(new_n620_), .A2(new_n615_), .ZN(new_n621_));
  NAND3_X1  g0557(.A1(new_n610_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n622_));
  AOI21_X1  g0558(.A(new_n462_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n623_));
  OAI211_X1 g0559(.A(new_n621_), .B(new_n622_), .C1(new_n623_), .C2(new_n579_), .ZN(new_n624_));
  AOI21_X1  g0560(.A(new_n575_), .B1(new_n619_), .B2(new_n624_), .ZN(new_n625_));
  AND3_X1   g0561(.A1(new_n619_), .A2(new_n624_), .A3(new_n575_), .ZN(new_n626_));
  OAI211_X1 g0562(.A(new_n569_), .B(new_n573_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g0563(.A1(new_n619_), .A2(new_n624_), .ZN(new_n628_));
  NAND2_X1  g0564(.A1(new_n628_), .A2(new_n574_), .ZN(new_n629_));
  NAND3_X1  g0565(.A1(new_n619_), .A2(new_n624_), .A3(new_n575_), .ZN(new_n630_));
  AOI21_X1  g0566(.A(new_n504_), .B1(new_n498_), .B2(new_n503_), .ZN(new_n631_));
  OAI211_X1 g0567(.A(new_n629_), .B(new_n630_), .C1(new_n631_), .C2(new_n572_), .ZN(new_n632_));
  NOR2_X1   g0568(.A1(new_n113_), .A2(new_n253_), .ZN(new_n633_));
  INV_X1    g0569(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g0570(.A1(new_n627_), .A2(new_n632_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g0571(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g0572(.A(new_n634_), .B1(new_n627_), .B2(new_n632_), .ZN(new_n637_));
  OAI211_X1 g0573(.A(new_n564_), .B(new_n568_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g0574(.A1(new_n627_), .A2(new_n632_), .ZN(new_n639_));
  NAND2_X1  g0575(.A1(new_n639_), .A2(new_n633_), .ZN(new_n640_));
  AOI21_X1  g0576(.A(new_n514_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n641_));
  OAI211_X1 g0577(.A(new_n640_), .B(new_n635_), .C1(new_n641_), .C2(new_n567_), .ZN(new_n642_));
  NOR2_X1   g0578(.A1(new_n86_), .A2(new_n336_), .ZN(new_n643_));
  INV_X1    g0579(.A(new_n643_), .ZN(new_n644_));
  NAND3_X1  g0580(.A1(new_n638_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g0581(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g0582(.A(new_n644_), .B1(new_n638_), .B2(new_n642_), .ZN(new_n647_));
  OAI211_X1 g0583(.A(new_n559_), .B(new_n563_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g0584(.A1(new_n638_), .A2(new_n642_), .ZN(new_n649_));
  NAND2_X1  g0585(.A1(new_n649_), .A2(new_n643_), .ZN(new_n650_));
  AOI21_X1  g0586(.A(new_n524_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n651_));
  OAI211_X1 g0587(.A(new_n650_), .B(new_n645_), .C1(new_n651_), .C2(new_n562_), .ZN(new_n652_));
  NOR2_X1   g0588(.A1(new_n76_), .A2(new_n432_), .ZN(new_n653_));
  INV_X1    g0589(.A(new_n653_), .ZN(new_n654_));
  AND3_X1   g0590(.A1(new_n648_), .A2(new_n652_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g0591(.A(new_n654_), .B1(new_n648_), .B2(new_n652_), .ZN(new_n656_));
  OAI211_X1 g0592(.A(new_n554_), .B(new_n558_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g0593(.A1(new_n648_), .A2(new_n652_), .ZN(new_n658_));
  NAND2_X1  g0594(.A1(new_n658_), .A2(new_n653_), .ZN(new_n659_));
  NAND3_X1  g0595(.A1(new_n648_), .A2(new_n652_), .A3(new_n654_), .ZN(new_n660_));
  AOI21_X1  g0596(.A(new_n534_), .B1(new_n528_), .B2(new_n533_), .ZN(new_n661_));
  OAI211_X1 g0597(.A(new_n659_), .B(new_n660_), .C1(new_n661_), .C2(new_n557_), .ZN(new_n662_));
  NOR2_X1   g0598(.A1(new_n68_), .A2(new_n544_), .ZN(new_n663_));
  INV_X1    g0599(.A(new_n663_), .ZN(new_n664_));
  NAND3_X1  g0600(.A1(new_n657_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g0601(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g0602(.A(new_n664_), .B1(new_n657_), .B2(new_n662_), .ZN(new_n667_));
  OAI211_X1 g0603(.A(new_n548_), .B(new_n552_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n668_));
  INV_X1    g0604(.A(new_n667_), .ZN(new_n669_));
  AOI21_X1  g0605(.A(new_n545_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n670_));
  OAI211_X1 g0606(.A(new_n669_), .B(new_n665_), .C1(new_n670_), .C2(new_n551_), .ZN(new_n671_));
  NAND2_X1  g0607(.A1(new_n668_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g0608(.A(G443gat), .ZN(new_n673_));
  NOR2_X1   g0609(.A1(new_n65_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g0610(.A(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g0611(.A(new_n672_), .B(new_n675_), .ZN(G4591gat));
  NAND2_X1  g0612(.A1(new_n672_), .A2(new_n675_), .ZN(new_n677_));
  NOR2_X1   g0613(.A1(new_n670_), .A2(new_n551_), .ZN(new_n678_));
  NOR2_X1   g0614(.A1(new_n666_), .A2(new_n667_), .ZN(new_n679_));
  NOR2_X1   g0615(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g0616(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g0617(.A1(new_n657_), .A2(new_n662_), .ZN(new_n682_));
  NAND2_X1  g0618(.A1(new_n682_), .A2(new_n664_), .ZN(new_n683_));
  NOR2_X1   g0619(.A1(new_n655_), .A2(new_n656_), .ZN(new_n684_));
  NOR2_X1   g0620(.A1(new_n661_), .A2(new_n557_), .ZN(new_n685_));
  NOR2_X1   g0621(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g0622(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g0623(.A1(new_n658_), .A2(new_n654_), .ZN(new_n688_));
  NOR2_X1   g0624(.A1(new_n646_), .A2(new_n647_), .ZN(new_n689_));
  NOR2_X1   g0625(.A1(new_n651_), .A2(new_n562_), .ZN(new_n690_));
  NOR2_X1   g0626(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g0627(.A(new_n691_), .ZN(new_n692_));
  NAND2_X1  g0628(.A1(new_n649_), .A2(new_n644_), .ZN(new_n693_));
  NOR2_X1   g0629(.A1(new_n636_), .A2(new_n637_), .ZN(new_n694_));
  NOR2_X1   g0630(.A1(new_n641_), .A2(new_n567_), .ZN(new_n695_));
  NOR2_X1   g0631(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g0632(.A(new_n696_), .ZN(new_n697_));
  NAND2_X1  g0633(.A1(new_n639_), .A2(new_n634_), .ZN(new_n698_));
  NOR2_X1   g0634(.A1(new_n626_), .A2(new_n625_), .ZN(new_n699_));
  NOR2_X1   g0635(.A1(new_n631_), .A2(new_n572_), .ZN(new_n700_));
  NOR2_X1   g0636(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g0637(.A(new_n701_), .ZN(new_n702_));
  NAND2_X1  g0638(.A1(new_n628_), .A2(new_n575_), .ZN(new_n703_));
  NOR2_X1   g0639(.A1(new_n617_), .A2(new_n618_), .ZN(new_n704_));
  NOR2_X1   g0640(.A1(new_n623_), .A2(new_n579_), .ZN(new_n705_));
  NOR2_X1   g0641(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g0642(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g0643(.A1(new_n620_), .A2(new_n616_), .ZN(new_n708_));
  NOR2_X1   g0644(.A1(new_n608_), .A2(new_n609_), .ZN(new_n709_));
  NOR2_X1   g0645(.A1(new_n613_), .A2(new_n582_), .ZN(new_n710_));
  NOR2_X1   g0646(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g0647(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g0648(.A(new_n592_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n713_));
  AOI21_X1  g0649(.A(new_n472_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n714_));
  NOR2_X1   g0650(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g0651(.A1(G154gat), .A2(G307gat), .ZN(new_n716_));
  INV_X1    g0652(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g0653(.A1(G171gat), .A2(G290gat), .ZN(new_n718_));
  INV_X1    g0654(.A(G188gat), .ZN(new_n719_));
  OAI21_X1  g0655(.A(new_n718_), .B1(new_n719_), .B2(new_n66_), .ZN(new_n720_));
  NAND4_X1  g0656(.A1(G171gat), .A2(G188gat), .A3(G273gat), .A4(G290gat), .ZN(new_n721_));
  AND3_X1   g0657(.A1(new_n720_), .A2(new_n586_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g0658(.A(new_n586_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n723_));
  OAI21_X1  g0659(.A(new_n717_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g0660(.A1(new_n720_), .A2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g0661(.A1(new_n725_), .A2(new_n588_), .ZN(new_n726_));
  NAND3_X1  g0662(.A1(new_n720_), .A2(new_n586_), .A3(new_n721_), .ZN(new_n727_));
  NAND3_X1  g0663(.A1(new_n726_), .A2(new_n727_), .A3(new_n716_), .ZN(new_n728_));
  NAND2_X1  g0664(.A1(new_n724_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g0665(.A1(new_n715_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g0666(.A(new_n724_), .B(new_n728_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n731_));
  NAND2_X1  g0667(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g0668(.A(G137gat), .ZN(new_n733_));
  NOR2_X1   g0669(.A1(new_n733_), .A2(new_n130_), .ZN(new_n734_));
  NAND2_X1  g0670(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g0671(.A(new_n734_), .ZN(new_n736_));
  NAND3_X1  g0672(.A1(new_n730_), .A2(new_n731_), .A3(new_n736_), .ZN(new_n737_));
  AOI22_X1  g0673(.A1(new_n601_), .A2(new_n600_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n738_));
  AOI21_X1  g0674(.A(new_n605_), .B1(new_n597_), .B2(new_n604_), .ZN(new_n739_));
  OAI211_X1 g0675(.A(new_n735_), .B(new_n737_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g0676(.A1(new_n611_), .A2(new_n606_), .ZN(new_n741_));
  INV_X1    g0677(.A(new_n738_), .ZN(new_n742_));
  AND3_X1   g0678(.A1(new_n730_), .A2(new_n731_), .A3(new_n736_), .ZN(new_n743_));
  AOI21_X1  g0679(.A(new_n736_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n744_));
  OAI211_X1 g0680(.A(new_n741_), .B(new_n742_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g0681(.A1(new_n276_), .A2(new_n178_), .ZN(new_n746_));
  INV_X1    g0682(.A(new_n746_), .ZN(new_n747_));
  NAND3_X1  g0683(.A1(new_n740_), .A2(new_n745_), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g0684(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g0685(.A(new_n747_), .B1(new_n740_), .B2(new_n745_), .ZN(new_n750_));
  OAI211_X1 g0686(.A(new_n708_), .B(new_n712_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g0687(.A1(new_n740_), .A2(new_n745_), .ZN(new_n752_));
  NAND2_X1  g0688(.A1(new_n752_), .A2(new_n746_), .ZN(new_n753_));
  AOI21_X1  g0689(.A(new_n615_), .B1(new_n610_), .B2(new_n614_), .ZN(new_n754_));
  OAI211_X1 g0690(.A(new_n753_), .B(new_n748_), .C1(new_n711_), .C2(new_n754_), .ZN(new_n755_));
  NOR2_X1   g0691(.A1(new_n205_), .A2(new_n190_), .ZN(new_n756_));
  INV_X1    g0692(.A(new_n756_), .ZN(new_n757_));
  NAND3_X1  g0693(.A1(new_n751_), .A2(new_n755_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g0694(.A(new_n758_), .ZN(new_n759_));
  AOI21_X1  g0695(.A(new_n757_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n760_));
  OAI211_X1 g0696(.A(new_n703_), .B(new_n707_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g0697(.A1(new_n751_), .A2(new_n755_), .ZN(new_n762_));
  NAND2_X1  g0698(.A1(new_n762_), .A2(new_n756_), .ZN(new_n763_));
  AOI21_X1  g0699(.A(new_n574_), .B1(new_n619_), .B2(new_n624_), .ZN(new_n764_));
  OAI211_X1 g0700(.A(new_n763_), .B(new_n758_), .C1(new_n706_), .C2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g0701(.A1(new_n146_), .A2(new_n253_), .ZN(new_n766_));
  INV_X1    g0702(.A(new_n766_), .ZN(new_n767_));
  NAND3_X1  g0703(.A1(new_n761_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g0704(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g0705(.A(new_n767_), .B1(new_n761_), .B2(new_n765_), .ZN(new_n770_));
  OAI211_X1 g0706(.A(new_n698_), .B(new_n702_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g0707(.A1(new_n761_), .A2(new_n765_), .ZN(new_n772_));
  NAND2_X1  g0708(.A1(new_n772_), .A2(new_n766_), .ZN(new_n773_));
  AOI21_X1  g0709(.A(new_n633_), .B1(new_n627_), .B2(new_n632_), .ZN(new_n774_));
  OAI211_X1 g0710(.A(new_n773_), .B(new_n768_), .C1(new_n701_), .C2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g0711(.A1(new_n113_), .A2(new_n336_), .ZN(new_n776_));
  INV_X1    g0712(.A(new_n776_), .ZN(new_n777_));
  NAND3_X1  g0713(.A1(new_n771_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g0714(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g0715(.A(new_n777_), .B1(new_n771_), .B2(new_n775_), .ZN(new_n780_));
  OAI211_X1 g0716(.A(new_n693_), .B(new_n697_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g0717(.A1(new_n771_), .A2(new_n775_), .ZN(new_n782_));
  NAND2_X1  g0718(.A1(new_n782_), .A2(new_n776_), .ZN(new_n783_));
  AOI21_X1  g0719(.A(new_n643_), .B1(new_n638_), .B2(new_n642_), .ZN(new_n784_));
  OAI211_X1 g0720(.A(new_n783_), .B(new_n778_), .C1(new_n784_), .C2(new_n696_), .ZN(new_n785_));
  NOR2_X1   g0721(.A1(new_n86_), .A2(new_n432_), .ZN(new_n786_));
  INV_X1    g0722(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g0723(.A1(new_n781_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g0724(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g0725(.A(new_n787_), .B1(new_n781_), .B2(new_n785_), .ZN(new_n790_));
  OAI211_X1 g0726(.A(new_n688_), .B(new_n692_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g0727(.A1(new_n781_), .A2(new_n785_), .ZN(new_n792_));
  NAND2_X1  g0728(.A1(new_n792_), .A2(new_n786_), .ZN(new_n793_));
  AOI21_X1  g0729(.A(new_n653_), .B1(new_n648_), .B2(new_n652_), .ZN(new_n794_));
  OAI211_X1 g0730(.A(new_n793_), .B(new_n788_), .C1(new_n794_), .C2(new_n691_), .ZN(new_n795_));
  NOR2_X1   g0731(.A1(new_n76_), .A2(new_n544_), .ZN(new_n796_));
  INV_X1    g0732(.A(new_n796_), .ZN(new_n797_));
  NAND3_X1  g0733(.A1(new_n791_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g0734(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g0735(.A(new_n797_), .B1(new_n791_), .B2(new_n795_), .ZN(new_n800_));
  OAI211_X1 g0736(.A(new_n683_), .B(new_n687_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g0737(.A1(new_n791_), .A2(new_n795_), .ZN(new_n802_));
  NAND2_X1  g0738(.A1(new_n802_), .A2(new_n796_), .ZN(new_n803_));
  AOI21_X1  g0739(.A(new_n663_), .B1(new_n657_), .B2(new_n662_), .ZN(new_n804_));
  OAI211_X1 g0740(.A(new_n803_), .B(new_n798_), .C1(new_n804_), .C2(new_n686_), .ZN(new_n805_));
  NOR2_X1   g0741(.A1(new_n68_), .A2(new_n673_), .ZN(new_n806_));
  INV_X1    g0742(.A(new_n806_), .ZN(new_n807_));
  NAND3_X1  g0743(.A1(new_n801_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g0744(.A(new_n808_), .ZN(new_n809_));
  AOI21_X1  g0745(.A(new_n807_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n810_));
  OAI211_X1 g0746(.A(new_n677_), .B(new_n681_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n811_));
  INV_X1    g0747(.A(new_n810_), .ZN(new_n812_));
  AOI21_X1  g0748(.A(new_n674_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n813_));
  OAI211_X1 g0749(.A(new_n812_), .B(new_n808_), .C1(new_n813_), .C2(new_n680_), .ZN(new_n814_));
  NAND2_X1  g0750(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g0751(.A(G460gat), .ZN(new_n816_));
  NOR2_X1   g0752(.A1(new_n65_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g0753(.A(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g0754(.A(new_n815_), .B(new_n818_), .ZN(G4946gat));
  NAND2_X1  g0755(.A1(new_n815_), .A2(new_n818_), .ZN(new_n820_));
  NOR2_X1   g0756(.A1(new_n813_), .A2(new_n680_), .ZN(new_n821_));
  NOR2_X1   g0757(.A1(new_n809_), .A2(new_n810_), .ZN(new_n822_));
  NOR2_X1   g0758(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g0759(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g0760(.A1(new_n801_), .A2(new_n805_), .ZN(new_n825_));
  NAND2_X1  g0761(.A1(new_n825_), .A2(new_n807_), .ZN(new_n826_));
  NOR2_X1   g0762(.A1(new_n799_), .A2(new_n800_), .ZN(new_n827_));
  NOR2_X1   g0763(.A1(new_n804_), .A2(new_n686_), .ZN(new_n828_));
  NOR2_X1   g0764(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g0765(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g0766(.A1(new_n802_), .A2(new_n797_), .ZN(new_n831_));
  NOR2_X1   g0767(.A1(new_n789_), .A2(new_n790_), .ZN(new_n832_));
  NOR2_X1   g0768(.A1(new_n794_), .A2(new_n691_), .ZN(new_n833_));
  NOR2_X1   g0769(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g0770(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g0771(.A1(new_n792_), .A2(new_n787_), .ZN(new_n836_));
  NOR2_X1   g0772(.A1(new_n779_), .A2(new_n780_), .ZN(new_n837_));
  NOR2_X1   g0773(.A1(new_n784_), .A2(new_n696_), .ZN(new_n838_));
  NOR2_X1   g0774(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g0775(.A(new_n839_), .ZN(new_n840_));
  NAND2_X1  g0776(.A1(new_n782_), .A2(new_n777_), .ZN(new_n841_));
  NOR2_X1   g0777(.A1(new_n769_), .A2(new_n770_), .ZN(new_n842_));
  NOR2_X1   g0778(.A1(new_n774_), .A2(new_n701_), .ZN(new_n843_));
  NOR2_X1   g0779(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g0780(.A(new_n844_), .ZN(new_n845_));
  NAND2_X1  g0781(.A1(new_n772_), .A2(new_n767_), .ZN(new_n846_));
  NOR2_X1   g0782(.A1(new_n759_), .A2(new_n760_), .ZN(new_n847_));
  NOR2_X1   g0783(.A1(new_n764_), .A2(new_n706_), .ZN(new_n848_));
  NOR2_X1   g0784(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g0785(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g0786(.A1(new_n762_), .A2(new_n757_), .ZN(new_n851_));
  NOR2_X1   g0787(.A1(new_n749_), .A2(new_n750_), .ZN(new_n852_));
  NOR2_X1   g0788(.A1(new_n754_), .A2(new_n711_), .ZN(new_n853_));
  NOR2_X1   g0789(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g0790(.A(new_n854_), .ZN(new_n855_));
  NAND2_X1  g0791(.A1(new_n752_), .A2(new_n747_), .ZN(new_n856_));
  NOR2_X1   g0792(.A1(new_n743_), .A2(new_n744_), .ZN(new_n857_));
  NOR2_X1   g0793(.A1(new_n739_), .A2(new_n738_), .ZN(new_n858_));
  NOR2_X1   g0794(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g0795(.A(new_n859_), .ZN(new_n860_));
  NAND2_X1  g0796(.A1(new_n732_), .A2(new_n736_), .ZN(new_n861_));
  AOI21_X1  g0797(.A(new_n715_), .B1(new_n724_), .B2(new_n728_), .ZN(new_n862_));
  INV_X1    g0798(.A(new_n862_), .ZN(new_n863_));
  AOI21_X1  g0799(.A(new_n588_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n864_));
  INV_X1    g0800(.A(new_n864_), .ZN(new_n865_));
  OAI21_X1  g0801(.A(new_n716_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n866_));
  INV_X1    g0802(.A(new_n721_), .ZN(new_n867_));
  NAND4_X1  g0803(.A1(G188gat), .A2(G205gat), .A3(G273gat), .A4(G290gat), .ZN(new_n868_));
  INV_X1    g0804(.A(new_n868_), .ZN(new_n869_));
  AOI22_X1  g0805(.A1(G188gat), .A2(G290gat), .B1(G205gat), .B2(G273gat), .ZN(new_n870_));
  OAI21_X1  g0806(.A(new_n867_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g0807(.A1(G188gat), .A2(G290gat), .ZN(new_n872_));
  INV_X1    g0808(.A(G205gat), .ZN(new_n873_));
  OAI21_X1  g0809(.A(new_n872_), .B1(new_n873_), .B2(new_n66_), .ZN(new_n874_));
  NAND3_X1  g0810(.A1(new_n874_), .A2(new_n721_), .A3(new_n868_), .ZN(new_n875_));
  INV_X1    g0811(.A(G171gat), .ZN(new_n876_));
  INV_X1    g0812(.A(G307gat), .ZN(new_n877_));
  NOR2_X1   g0813(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g0814(.A(new_n878_), .ZN(new_n879_));
  NAND3_X1  g0815(.A1(new_n871_), .A2(new_n875_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g0816(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g0817(.A(new_n879_), .B1(new_n871_), .B2(new_n875_), .ZN(new_n882_));
  OAI211_X1 g0818(.A(new_n865_), .B(new_n866_), .C1(new_n881_), .C2(new_n882_), .ZN(new_n883_));
  AND3_X1   g0819(.A1(new_n874_), .A2(new_n721_), .A3(new_n868_), .ZN(new_n884_));
  AOI21_X1  g0820(.A(new_n721_), .B1(new_n874_), .B2(new_n868_), .ZN(new_n885_));
  OAI21_X1  g0821(.A(new_n878_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g0822(.A(new_n717_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n887_));
  OAI211_X1 g0823(.A(new_n886_), .B(new_n880_), .C1(new_n887_), .C2(new_n864_), .ZN(new_n888_));
  INV_X1    g0824(.A(G154gat), .ZN(new_n889_));
  NOR2_X1   g0825(.A1(new_n889_), .A2(new_n130_), .ZN(new_n890_));
  INV_X1    g0826(.A(new_n890_), .ZN(new_n891_));
  NAND3_X1  g0827(.A1(new_n883_), .A2(new_n888_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g0828(.A(new_n892_), .ZN(new_n893_));
  AOI21_X1  g0829(.A(new_n891_), .B1(new_n883_), .B2(new_n888_), .ZN(new_n894_));
  OAI211_X1 g0830(.A(new_n861_), .B(new_n863_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g0831(.A1(new_n883_), .A2(new_n888_), .ZN(new_n896_));
  NAND2_X1  g0832(.A1(new_n896_), .A2(new_n890_), .ZN(new_n897_));
  AOI21_X1  g0833(.A(new_n734_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n898_));
  OAI211_X1 g0834(.A(new_n897_), .B(new_n892_), .C1(new_n862_), .C2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g0835(.A1(new_n733_), .A2(new_n178_), .ZN(new_n900_));
  INV_X1    g0836(.A(new_n900_), .ZN(new_n901_));
  NAND3_X1  g0837(.A1(new_n895_), .A2(new_n899_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g0838(.A(new_n902_), .ZN(new_n903_));
  AOI21_X1  g0839(.A(new_n901_), .B1(new_n895_), .B2(new_n899_), .ZN(new_n904_));
  OAI211_X1 g0840(.A(new_n856_), .B(new_n860_), .C1(new_n903_), .C2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g0841(.A1(new_n895_), .A2(new_n899_), .ZN(new_n906_));
  NAND2_X1  g0842(.A1(new_n906_), .A2(new_n900_), .ZN(new_n907_));
  AOI21_X1  g0843(.A(new_n746_), .B1(new_n740_), .B2(new_n745_), .ZN(new_n908_));
  OAI211_X1 g0844(.A(new_n907_), .B(new_n902_), .C1(new_n859_), .C2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g0845(.A1(new_n276_), .A2(new_n190_), .ZN(new_n910_));
  INV_X1    g0846(.A(new_n910_), .ZN(new_n911_));
  NAND3_X1  g0847(.A1(new_n905_), .A2(new_n909_), .A3(new_n911_), .ZN(new_n912_));
  INV_X1    g0848(.A(new_n912_), .ZN(new_n913_));
  AOI21_X1  g0849(.A(new_n911_), .B1(new_n905_), .B2(new_n909_), .ZN(new_n914_));
  OAI211_X1 g0850(.A(new_n851_), .B(new_n855_), .C1(new_n913_), .C2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g0851(.A1(new_n905_), .A2(new_n909_), .ZN(new_n916_));
  NAND2_X1  g0852(.A1(new_n916_), .A2(new_n910_), .ZN(new_n917_));
  AOI21_X1  g0853(.A(new_n756_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n918_));
  OAI211_X1 g0854(.A(new_n917_), .B(new_n912_), .C1(new_n854_), .C2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g0855(.A1(new_n205_), .A2(new_n253_), .ZN(new_n920_));
  INV_X1    g0856(.A(new_n920_), .ZN(new_n921_));
  NAND3_X1  g0857(.A1(new_n915_), .A2(new_n919_), .A3(new_n921_), .ZN(new_n922_));
  INV_X1    g0858(.A(new_n922_), .ZN(new_n923_));
  AOI21_X1  g0859(.A(new_n921_), .B1(new_n915_), .B2(new_n919_), .ZN(new_n924_));
  OAI211_X1 g0860(.A(new_n846_), .B(new_n850_), .C1(new_n923_), .C2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g0861(.A1(new_n915_), .A2(new_n919_), .ZN(new_n926_));
  NAND2_X1  g0862(.A1(new_n926_), .A2(new_n920_), .ZN(new_n927_));
  AOI21_X1  g0863(.A(new_n766_), .B1(new_n761_), .B2(new_n765_), .ZN(new_n928_));
  OAI211_X1 g0864(.A(new_n927_), .B(new_n922_), .C1(new_n849_), .C2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g0865(.A1(new_n146_), .A2(new_n336_), .ZN(new_n930_));
  INV_X1    g0866(.A(new_n930_), .ZN(new_n931_));
  NAND3_X1  g0867(.A1(new_n925_), .A2(new_n929_), .A3(new_n931_), .ZN(new_n932_));
  INV_X1    g0868(.A(new_n932_), .ZN(new_n933_));
  AOI21_X1  g0869(.A(new_n931_), .B1(new_n925_), .B2(new_n929_), .ZN(new_n934_));
  OAI211_X1 g0870(.A(new_n841_), .B(new_n845_), .C1(new_n933_), .C2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g0871(.A1(new_n925_), .A2(new_n929_), .ZN(new_n936_));
  NAND2_X1  g0872(.A1(new_n936_), .A2(new_n930_), .ZN(new_n937_));
  AOI21_X1  g0873(.A(new_n776_), .B1(new_n771_), .B2(new_n775_), .ZN(new_n938_));
  OAI211_X1 g0874(.A(new_n937_), .B(new_n932_), .C1(new_n844_), .C2(new_n938_), .ZN(new_n939_));
  NOR2_X1   g0875(.A1(new_n113_), .A2(new_n432_), .ZN(new_n940_));
  INV_X1    g0876(.A(new_n940_), .ZN(new_n941_));
  NAND3_X1  g0877(.A1(new_n935_), .A2(new_n939_), .A3(new_n941_), .ZN(new_n942_));
  INV_X1    g0878(.A(new_n942_), .ZN(new_n943_));
  AOI21_X1  g0879(.A(new_n941_), .B1(new_n935_), .B2(new_n939_), .ZN(new_n944_));
  OAI211_X1 g0880(.A(new_n836_), .B(new_n840_), .C1(new_n943_), .C2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g0881(.A1(new_n935_), .A2(new_n939_), .ZN(new_n946_));
  NAND2_X1  g0882(.A1(new_n946_), .A2(new_n940_), .ZN(new_n947_));
  AOI21_X1  g0883(.A(new_n786_), .B1(new_n781_), .B2(new_n785_), .ZN(new_n948_));
  OAI211_X1 g0884(.A(new_n947_), .B(new_n942_), .C1(new_n948_), .C2(new_n839_), .ZN(new_n949_));
  NOR2_X1   g0885(.A1(new_n86_), .A2(new_n544_), .ZN(new_n950_));
  INV_X1    g0886(.A(new_n950_), .ZN(new_n951_));
  NAND3_X1  g0887(.A1(new_n945_), .A2(new_n949_), .A3(new_n951_), .ZN(new_n952_));
  INV_X1    g0888(.A(new_n952_), .ZN(new_n953_));
  AOI21_X1  g0889(.A(new_n951_), .B1(new_n945_), .B2(new_n949_), .ZN(new_n954_));
  OAI211_X1 g0890(.A(new_n831_), .B(new_n835_), .C1(new_n953_), .C2(new_n954_), .ZN(new_n955_));
  NAND2_X1  g0891(.A1(new_n945_), .A2(new_n949_), .ZN(new_n956_));
  NAND2_X1  g0892(.A1(new_n956_), .A2(new_n950_), .ZN(new_n957_));
  AOI21_X1  g0893(.A(new_n796_), .B1(new_n791_), .B2(new_n795_), .ZN(new_n958_));
  OAI211_X1 g0894(.A(new_n957_), .B(new_n952_), .C1(new_n958_), .C2(new_n834_), .ZN(new_n959_));
  NOR2_X1   g0895(.A1(new_n76_), .A2(new_n673_), .ZN(new_n960_));
  INV_X1    g0896(.A(new_n960_), .ZN(new_n961_));
  NAND3_X1  g0897(.A1(new_n955_), .A2(new_n959_), .A3(new_n961_), .ZN(new_n962_));
  INV_X1    g0898(.A(new_n962_), .ZN(new_n963_));
  AOI21_X1  g0899(.A(new_n961_), .B1(new_n955_), .B2(new_n959_), .ZN(new_n964_));
  OAI211_X1 g0900(.A(new_n826_), .B(new_n830_), .C1(new_n963_), .C2(new_n964_), .ZN(new_n965_));
  NAND2_X1  g0901(.A1(new_n955_), .A2(new_n959_), .ZN(new_n966_));
  NAND2_X1  g0902(.A1(new_n966_), .A2(new_n960_), .ZN(new_n967_));
  AOI21_X1  g0903(.A(new_n806_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n968_));
  OAI211_X1 g0904(.A(new_n967_), .B(new_n962_), .C1(new_n968_), .C2(new_n829_), .ZN(new_n969_));
  NOR2_X1   g0905(.A1(new_n68_), .A2(new_n816_), .ZN(new_n970_));
  INV_X1    g0906(.A(new_n970_), .ZN(new_n971_));
  NAND3_X1  g0907(.A1(new_n965_), .A2(new_n969_), .A3(new_n971_), .ZN(new_n972_));
  INV_X1    g0908(.A(new_n972_), .ZN(new_n973_));
  AOI21_X1  g0909(.A(new_n971_), .B1(new_n965_), .B2(new_n969_), .ZN(new_n974_));
  OAI211_X1 g0910(.A(new_n820_), .B(new_n824_), .C1(new_n973_), .C2(new_n974_), .ZN(new_n975_));
  INV_X1    g0911(.A(new_n974_), .ZN(new_n976_));
  AOI21_X1  g0912(.A(new_n817_), .B1(new_n811_), .B2(new_n814_), .ZN(new_n977_));
  OAI211_X1 g0913(.A(new_n976_), .B(new_n972_), .C1(new_n977_), .C2(new_n823_), .ZN(new_n978_));
  NAND2_X1  g0914(.A1(new_n975_), .A2(new_n978_), .ZN(new_n979_));
  INV_X1    g0915(.A(G477gat), .ZN(new_n980_));
  NOR2_X1   g0916(.A1(new_n65_), .A2(new_n980_), .ZN(new_n981_));
  INV_X1    g0917(.A(new_n981_), .ZN(new_n982_));
  XNOR2_X1  g0918(.A(new_n979_), .B(new_n982_), .ZN(G5308gat));
  NAND2_X1  g0919(.A1(new_n979_), .A2(new_n982_), .ZN(new_n984_));
  NOR2_X1   g0920(.A1(new_n977_), .A2(new_n823_), .ZN(new_n985_));
  NOR2_X1   g0921(.A1(new_n973_), .A2(new_n974_), .ZN(new_n986_));
  NOR2_X1   g0922(.A1(new_n985_), .A2(new_n986_), .ZN(new_n987_));
  INV_X1    g0923(.A(new_n987_), .ZN(new_n988_));
  NAND2_X1  g0924(.A1(new_n965_), .A2(new_n969_), .ZN(new_n989_));
  NAND2_X1  g0925(.A1(new_n989_), .A2(new_n971_), .ZN(new_n990_));
  NOR2_X1   g0926(.A1(new_n963_), .A2(new_n964_), .ZN(new_n991_));
  NOR2_X1   g0927(.A1(new_n968_), .A2(new_n829_), .ZN(new_n992_));
  NOR2_X1   g0928(.A1(new_n991_), .A2(new_n992_), .ZN(new_n993_));
  INV_X1    g0929(.A(new_n993_), .ZN(new_n994_));
  NAND2_X1  g0930(.A1(new_n966_), .A2(new_n961_), .ZN(new_n995_));
  NOR2_X1   g0931(.A1(new_n953_), .A2(new_n954_), .ZN(new_n996_));
  NOR2_X1   g0932(.A1(new_n958_), .A2(new_n834_), .ZN(new_n997_));
  NOR2_X1   g0933(.A1(new_n996_), .A2(new_n997_), .ZN(new_n998_));
  INV_X1    g0934(.A(new_n998_), .ZN(new_n999_));
  NAND2_X1  g0935(.A1(new_n956_), .A2(new_n951_), .ZN(new_n1000_));
  NOR2_X1   g0936(.A1(new_n943_), .A2(new_n944_), .ZN(new_n1001_));
  NOR2_X1   g0937(.A1(new_n948_), .A2(new_n839_), .ZN(new_n1002_));
  NOR2_X1   g0938(.A1(new_n1001_), .A2(new_n1002_), .ZN(new_n1003_));
  INV_X1    g0939(.A(new_n1003_), .ZN(new_n1004_));
  NAND2_X1  g0940(.A1(new_n946_), .A2(new_n941_), .ZN(new_n1005_));
  NOR2_X1   g0941(.A1(new_n933_), .A2(new_n934_), .ZN(new_n1006_));
  NOR2_X1   g0942(.A1(new_n938_), .A2(new_n844_), .ZN(new_n1007_));
  NOR2_X1   g0943(.A1(new_n1006_), .A2(new_n1007_), .ZN(new_n1008_));
  INV_X1    g0944(.A(new_n1008_), .ZN(new_n1009_));
  NAND2_X1  g0945(.A1(new_n936_), .A2(new_n931_), .ZN(new_n1010_));
  NOR2_X1   g0946(.A1(new_n923_), .A2(new_n924_), .ZN(new_n1011_));
  NOR2_X1   g0947(.A1(new_n928_), .A2(new_n849_), .ZN(new_n1012_));
  NOR2_X1   g0948(.A1(new_n1011_), .A2(new_n1012_), .ZN(new_n1013_));
  INV_X1    g0949(.A(new_n1013_), .ZN(new_n1014_));
  NAND2_X1  g0950(.A1(new_n926_), .A2(new_n921_), .ZN(new_n1015_));
  NOR2_X1   g0951(.A1(new_n913_), .A2(new_n914_), .ZN(new_n1016_));
  NOR2_X1   g0952(.A1(new_n918_), .A2(new_n854_), .ZN(new_n1017_));
  NOR2_X1   g0953(.A1(new_n1016_), .A2(new_n1017_), .ZN(new_n1018_));
  INV_X1    g0954(.A(new_n1018_), .ZN(new_n1019_));
  NAND2_X1  g0955(.A1(new_n916_), .A2(new_n911_), .ZN(new_n1020_));
  NOR2_X1   g0956(.A1(new_n903_), .A2(new_n904_), .ZN(new_n1021_));
  NOR2_X1   g0957(.A1(new_n908_), .A2(new_n859_), .ZN(new_n1022_));
  NOR2_X1   g0958(.A1(new_n1021_), .A2(new_n1022_), .ZN(new_n1023_));
  INV_X1    g0959(.A(new_n1023_), .ZN(new_n1024_));
  NAND2_X1  g0960(.A1(new_n906_), .A2(new_n901_), .ZN(new_n1025_));
  NOR2_X1   g0961(.A1(new_n893_), .A2(new_n894_), .ZN(new_n1026_));
  NOR2_X1   g0962(.A1(new_n898_), .A2(new_n862_), .ZN(new_n1027_));
  NOR2_X1   g0963(.A1(new_n1026_), .A2(new_n1027_), .ZN(new_n1028_));
  INV_X1    g0964(.A(new_n1028_), .ZN(new_n1029_));
  NAND2_X1  g0965(.A1(new_n896_), .A2(new_n891_), .ZN(new_n1030_));
  AOI22_X1  g0966(.A1(new_n865_), .A2(new_n866_), .B1(new_n886_), .B2(new_n880_), .ZN(new_n1031_));
  INV_X1    g0967(.A(new_n1031_), .ZN(new_n1032_));
  NOR2_X1   g0968(.A1(new_n876_), .A2(new_n130_), .ZN(new_n1033_));
  INV_X1    g0969(.A(new_n1033_), .ZN(new_n1034_));
  NAND2_X1  g0970(.A1(G188gat), .A2(G307gat), .ZN(new_n1035_));
  INV_X1    g0971(.A(new_n1035_), .ZN(new_n1036_));
  AND4_X1   g0972(.A1(G205gat), .A2(G222gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1037_));
  AOI22_X1  g0973(.A1(G205gat), .A2(G290gat), .B1(G222gat), .B2(G273gat), .ZN(new_n1038_));
  NOR3_X1   g0974(.A1(new_n869_), .A2(new_n1037_), .A3(new_n1038_), .ZN(new_n1039_));
  NAND2_X1  g0975(.A1(G205gat), .A2(G290gat), .ZN(new_n1040_));
  INV_X1    g0976(.A(G222gat), .ZN(new_n1041_));
  OAI21_X1  g0977(.A(new_n1040_), .B1(new_n1041_), .B2(new_n66_), .ZN(new_n1042_));
  NAND4_X1  g0978(.A1(G205gat), .A2(G222gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1043_));
  AOI21_X1  g0979(.A(new_n868_), .B1(new_n1042_), .B2(new_n1043_), .ZN(new_n1044_));
  OAI21_X1  g0980(.A(new_n1036_), .B1(new_n1039_), .B2(new_n1044_), .ZN(new_n1045_));
  OAI21_X1  g0981(.A(new_n869_), .B1(new_n1037_), .B2(new_n1038_), .ZN(new_n1046_));
  NAND3_X1  g0982(.A1(new_n1042_), .A2(new_n868_), .A3(new_n1043_), .ZN(new_n1047_));
  NAND3_X1  g0983(.A1(new_n1046_), .A2(new_n1047_), .A3(new_n1035_), .ZN(new_n1048_));
  AOI21_X1  g0984(.A(new_n878_), .B1(new_n871_), .B2(new_n875_), .ZN(new_n1049_));
  AOI21_X1  g0985(.A(new_n867_), .B1(new_n868_), .B2(new_n874_), .ZN(new_n1050_));
  OAI211_X1 g0986(.A(new_n1045_), .B(new_n1048_), .C1(new_n1049_), .C2(new_n1050_), .ZN(new_n1051_));
  OAI21_X1  g0987(.A(new_n879_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n1052_));
  INV_X1    g0988(.A(new_n1050_), .ZN(new_n1053_));
  AND3_X1   g0989(.A1(new_n1046_), .A2(new_n1047_), .A3(new_n1035_), .ZN(new_n1054_));
  AOI21_X1  g0990(.A(new_n1035_), .B1(new_n1046_), .B2(new_n1047_), .ZN(new_n1055_));
  OAI211_X1 g0991(.A(new_n1052_), .B(new_n1053_), .C1(new_n1054_), .C2(new_n1055_), .ZN(new_n1056_));
  AOI21_X1  g0992(.A(new_n1034_), .B1(new_n1051_), .B2(new_n1056_), .ZN(new_n1057_));
  AND3_X1   g0993(.A1(new_n1051_), .A2(new_n1056_), .A3(new_n1034_), .ZN(new_n1058_));
  OAI211_X1 g0994(.A(new_n1030_), .B(new_n1032_), .C1(new_n1057_), .C2(new_n1058_), .ZN(new_n1059_));
  NAND2_X1  g0995(.A1(new_n1051_), .A2(new_n1056_), .ZN(new_n1060_));
  NAND2_X1  g0996(.A1(new_n1060_), .A2(new_n1033_), .ZN(new_n1061_));
  NAND3_X1  g0997(.A1(new_n1051_), .A2(new_n1056_), .A3(new_n1034_), .ZN(new_n1062_));
  AOI21_X1  g0998(.A(new_n890_), .B1(new_n883_), .B2(new_n888_), .ZN(new_n1063_));
  OAI211_X1 g0999(.A(new_n1061_), .B(new_n1062_), .C1(new_n1063_), .C2(new_n1031_), .ZN(new_n1064_));
  NOR2_X1   g1000(.A1(new_n889_), .A2(new_n178_), .ZN(new_n1065_));
  INV_X1    g1001(.A(new_n1065_), .ZN(new_n1066_));
  NAND3_X1  g1002(.A1(new_n1059_), .A2(new_n1064_), .A3(new_n1066_), .ZN(new_n1067_));
  INV_X1    g1003(.A(new_n1067_), .ZN(new_n1068_));
  AOI21_X1  g1004(.A(new_n1066_), .B1(new_n1059_), .B2(new_n1064_), .ZN(new_n1069_));
  OAI211_X1 g1005(.A(new_n1025_), .B(new_n1029_), .C1(new_n1068_), .C2(new_n1069_), .ZN(new_n1070_));
  NAND2_X1  g1006(.A1(new_n1059_), .A2(new_n1064_), .ZN(new_n1071_));
  NAND2_X1  g1007(.A1(new_n1071_), .A2(new_n1065_), .ZN(new_n1072_));
  AOI21_X1  g1008(.A(new_n900_), .B1(new_n895_), .B2(new_n899_), .ZN(new_n1073_));
  OAI211_X1 g1009(.A(new_n1072_), .B(new_n1067_), .C1(new_n1073_), .C2(new_n1028_), .ZN(new_n1074_));
  NOR2_X1   g1010(.A1(new_n733_), .A2(new_n190_), .ZN(new_n1075_));
  INV_X1    g1011(.A(new_n1075_), .ZN(new_n1076_));
  NAND3_X1  g1012(.A1(new_n1070_), .A2(new_n1074_), .A3(new_n1076_), .ZN(new_n1077_));
  INV_X1    g1013(.A(new_n1077_), .ZN(new_n1078_));
  AOI21_X1  g1014(.A(new_n1076_), .B1(new_n1070_), .B2(new_n1074_), .ZN(new_n1079_));
  OAI211_X1 g1015(.A(new_n1020_), .B(new_n1024_), .C1(new_n1078_), .C2(new_n1079_), .ZN(new_n1080_));
  NAND2_X1  g1016(.A1(new_n1070_), .A2(new_n1074_), .ZN(new_n1081_));
  NAND2_X1  g1017(.A1(new_n1081_), .A2(new_n1075_), .ZN(new_n1082_));
  AOI21_X1  g1018(.A(new_n910_), .B1(new_n905_), .B2(new_n909_), .ZN(new_n1083_));
  OAI211_X1 g1019(.A(new_n1082_), .B(new_n1077_), .C1(new_n1083_), .C2(new_n1023_), .ZN(new_n1084_));
  NOR2_X1   g1020(.A1(new_n276_), .A2(new_n253_), .ZN(new_n1085_));
  INV_X1    g1021(.A(new_n1085_), .ZN(new_n1086_));
  NAND3_X1  g1022(.A1(new_n1080_), .A2(new_n1084_), .A3(new_n1086_), .ZN(new_n1087_));
  INV_X1    g1023(.A(new_n1087_), .ZN(new_n1088_));
  AOI21_X1  g1024(.A(new_n1086_), .B1(new_n1080_), .B2(new_n1084_), .ZN(new_n1089_));
  OAI211_X1 g1025(.A(new_n1015_), .B(new_n1019_), .C1(new_n1088_), .C2(new_n1089_), .ZN(new_n1090_));
  NAND2_X1  g1026(.A1(new_n1080_), .A2(new_n1084_), .ZN(new_n1091_));
  NAND2_X1  g1027(.A1(new_n1091_), .A2(new_n1085_), .ZN(new_n1092_));
  AOI21_X1  g1028(.A(new_n920_), .B1(new_n915_), .B2(new_n919_), .ZN(new_n1093_));
  OAI211_X1 g1029(.A(new_n1092_), .B(new_n1087_), .C1(new_n1093_), .C2(new_n1018_), .ZN(new_n1094_));
  NOR2_X1   g1030(.A1(new_n205_), .A2(new_n336_), .ZN(new_n1095_));
  INV_X1    g1031(.A(new_n1095_), .ZN(new_n1096_));
  NAND3_X1  g1032(.A1(new_n1090_), .A2(new_n1094_), .A3(new_n1096_), .ZN(new_n1097_));
  INV_X1    g1033(.A(new_n1097_), .ZN(new_n1098_));
  AOI21_X1  g1034(.A(new_n1096_), .B1(new_n1090_), .B2(new_n1094_), .ZN(new_n1099_));
  OAI211_X1 g1035(.A(new_n1010_), .B(new_n1014_), .C1(new_n1098_), .C2(new_n1099_), .ZN(new_n1100_));
  NAND2_X1  g1036(.A1(new_n1090_), .A2(new_n1094_), .ZN(new_n1101_));
  NAND2_X1  g1037(.A1(new_n1101_), .A2(new_n1095_), .ZN(new_n1102_));
  AOI21_X1  g1038(.A(new_n930_), .B1(new_n925_), .B2(new_n929_), .ZN(new_n1103_));
  OAI211_X1 g1039(.A(new_n1102_), .B(new_n1097_), .C1(new_n1103_), .C2(new_n1013_), .ZN(new_n1104_));
  NOR2_X1   g1040(.A1(new_n146_), .A2(new_n432_), .ZN(new_n1105_));
  INV_X1    g1041(.A(new_n1105_), .ZN(new_n1106_));
  NAND3_X1  g1042(.A1(new_n1100_), .A2(new_n1104_), .A3(new_n1106_), .ZN(new_n1107_));
  INV_X1    g1043(.A(new_n1107_), .ZN(new_n1108_));
  AOI21_X1  g1044(.A(new_n1106_), .B1(new_n1100_), .B2(new_n1104_), .ZN(new_n1109_));
  OAI211_X1 g1045(.A(new_n1005_), .B(new_n1009_), .C1(new_n1108_), .C2(new_n1109_), .ZN(new_n1110_));
  NAND2_X1  g1046(.A1(new_n1100_), .A2(new_n1104_), .ZN(new_n1111_));
  NAND2_X1  g1047(.A1(new_n1111_), .A2(new_n1105_), .ZN(new_n1112_));
  AOI21_X1  g1048(.A(new_n940_), .B1(new_n935_), .B2(new_n939_), .ZN(new_n1113_));
  OAI211_X1 g1049(.A(new_n1112_), .B(new_n1107_), .C1(new_n1113_), .C2(new_n1008_), .ZN(new_n1114_));
  NOR2_X1   g1050(.A1(new_n113_), .A2(new_n544_), .ZN(new_n1115_));
  INV_X1    g1051(.A(new_n1115_), .ZN(new_n1116_));
  NAND3_X1  g1052(.A1(new_n1110_), .A2(new_n1114_), .A3(new_n1116_), .ZN(new_n1117_));
  INV_X1    g1053(.A(new_n1117_), .ZN(new_n1118_));
  AOI21_X1  g1054(.A(new_n1116_), .B1(new_n1110_), .B2(new_n1114_), .ZN(new_n1119_));
  OAI211_X1 g1055(.A(new_n1000_), .B(new_n1004_), .C1(new_n1118_), .C2(new_n1119_), .ZN(new_n1120_));
  NAND2_X1  g1056(.A1(new_n1110_), .A2(new_n1114_), .ZN(new_n1121_));
  NAND2_X1  g1057(.A1(new_n1121_), .A2(new_n1115_), .ZN(new_n1122_));
  AOI21_X1  g1058(.A(new_n950_), .B1(new_n945_), .B2(new_n949_), .ZN(new_n1123_));
  OAI211_X1 g1059(.A(new_n1122_), .B(new_n1117_), .C1(new_n1123_), .C2(new_n1003_), .ZN(new_n1124_));
  NOR2_X1   g1060(.A1(new_n86_), .A2(new_n673_), .ZN(new_n1125_));
  INV_X1    g1061(.A(new_n1125_), .ZN(new_n1126_));
  NAND3_X1  g1062(.A1(new_n1120_), .A2(new_n1124_), .A3(new_n1126_), .ZN(new_n1127_));
  INV_X1    g1063(.A(new_n1127_), .ZN(new_n1128_));
  AOI21_X1  g1064(.A(new_n1126_), .B1(new_n1120_), .B2(new_n1124_), .ZN(new_n1129_));
  OAI211_X1 g1065(.A(new_n995_), .B(new_n999_), .C1(new_n1128_), .C2(new_n1129_), .ZN(new_n1130_));
  NAND2_X1  g1066(.A1(new_n1120_), .A2(new_n1124_), .ZN(new_n1131_));
  NAND2_X1  g1067(.A1(new_n1131_), .A2(new_n1125_), .ZN(new_n1132_));
  AOI21_X1  g1068(.A(new_n960_), .B1(new_n955_), .B2(new_n959_), .ZN(new_n1133_));
  OAI211_X1 g1069(.A(new_n1132_), .B(new_n1127_), .C1(new_n1133_), .C2(new_n998_), .ZN(new_n1134_));
  NOR2_X1   g1070(.A1(new_n76_), .A2(new_n816_), .ZN(new_n1135_));
  INV_X1    g1071(.A(new_n1135_), .ZN(new_n1136_));
  NAND3_X1  g1072(.A1(new_n1130_), .A2(new_n1134_), .A3(new_n1136_), .ZN(new_n1137_));
  INV_X1    g1073(.A(new_n1137_), .ZN(new_n1138_));
  AOI21_X1  g1074(.A(new_n1136_), .B1(new_n1130_), .B2(new_n1134_), .ZN(new_n1139_));
  OAI211_X1 g1075(.A(new_n990_), .B(new_n994_), .C1(new_n1138_), .C2(new_n1139_), .ZN(new_n1140_));
  NAND2_X1  g1076(.A1(new_n1130_), .A2(new_n1134_), .ZN(new_n1141_));
  NAND2_X1  g1077(.A1(new_n1141_), .A2(new_n1135_), .ZN(new_n1142_));
  AOI21_X1  g1078(.A(new_n970_), .B1(new_n965_), .B2(new_n969_), .ZN(new_n1143_));
  OAI211_X1 g1079(.A(new_n1142_), .B(new_n1137_), .C1(new_n1143_), .C2(new_n993_), .ZN(new_n1144_));
  NOR2_X1   g1080(.A1(new_n68_), .A2(new_n980_), .ZN(new_n1145_));
  INV_X1    g1081(.A(new_n1145_), .ZN(new_n1146_));
  NAND3_X1  g1082(.A1(new_n1140_), .A2(new_n1144_), .A3(new_n1146_), .ZN(new_n1147_));
  INV_X1    g1083(.A(new_n1147_), .ZN(new_n1148_));
  AOI21_X1  g1084(.A(new_n1146_), .B1(new_n1140_), .B2(new_n1144_), .ZN(new_n1149_));
  OAI211_X1 g1085(.A(new_n984_), .B(new_n988_), .C1(new_n1148_), .C2(new_n1149_), .ZN(new_n1150_));
  INV_X1    g1086(.A(new_n1149_), .ZN(new_n1151_));
  AOI21_X1  g1087(.A(new_n981_), .B1(new_n975_), .B2(new_n978_), .ZN(new_n1152_));
  OAI211_X1 g1088(.A(new_n1151_), .B(new_n1147_), .C1(new_n1152_), .C2(new_n987_), .ZN(new_n1153_));
  NAND2_X1  g1089(.A1(new_n1150_), .A2(new_n1153_), .ZN(new_n1154_));
  INV_X1    g1090(.A(G494gat), .ZN(new_n1155_));
  NOR2_X1   g1091(.A1(new_n65_), .A2(new_n1155_), .ZN(new_n1156_));
  INV_X1    g1092(.A(new_n1156_), .ZN(new_n1157_));
  XNOR2_X1  g1093(.A(new_n1154_), .B(new_n1157_), .ZN(G5672gat));
  NAND2_X1  g1094(.A1(new_n1154_), .A2(new_n1157_), .ZN(new_n1159_));
  NOR2_X1   g1095(.A1(new_n1152_), .A2(new_n987_), .ZN(new_n1160_));
  NOR2_X1   g1096(.A1(new_n1148_), .A2(new_n1149_), .ZN(new_n1161_));
  NOR2_X1   g1097(.A1(new_n1160_), .A2(new_n1161_), .ZN(new_n1162_));
  INV_X1    g1098(.A(new_n1162_), .ZN(new_n1163_));
  NAND2_X1  g1099(.A1(new_n1140_), .A2(new_n1144_), .ZN(new_n1164_));
  NAND2_X1  g1100(.A1(new_n1164_), .A2(new_n1146_), .ZN(new_n1165_));
  NOR2_X1   g1101(.A1(new_n1138_), .A2(new_n1139_), .ZN(new_n1166_));
  NOR2_X1   g1102(.A1(new_n1143_), .A2(new_n993_), .ZN(new_n1167_));
  NOR2_X1   g1103(.A1(new_n1166_), .A2(new_n1167_), .ZN(new_n1168_));
  INV_X1    g1104(.A(new_n1168_), .ZN(new_n1169_));
  NAND2_X1  g1105(.A1(new_n1141_), .A2(new_n1136_), .ZN(new_n1170_));
  NOR2_X1   g1106(.A1(new_n1128_), .A2(new_n1129_), .ZN(new_n1171_));
  NOR2_X1   g1107(.A1(new_n1133_), .A2(new_n998_), .ZN(new_n1172_));
  NOR2_X1   g1108(.A1(new_n1171_), .A2(new_n1172_), .ZN(new_n1173_));
  INV_X1    g1109(.A(new_n1173_), .ZN(new_n1174_));
  NAND2_X1  g1110(.A1(new_n1131_), .A2(new_n1126_), .ZN(new_n1175_));
  NOR2_X1   g1111(.A1(new_n1118_), .A2(new_n1119_), .ZN(new_n1176_));
  NOR2_X1   g1112(.A1(new_n1123_), .A2(new_n1003_), .ZN(new_n1177_));
  NOR2_X1   g1113(.A1(new_n1176_), .A2(new_n1177_), .ZN(new_n1178_));
  INV_X1    g1114(.A(new_n1178_), .ZN(new_n1179_));
  NAND2_X1  g1115(.A1(new_n1121_), .A2(new_n1116_), .ZN(new_n1180_));
  NOR2_X1   g1116(.A1(new_n1108_), .A2(new_n1109_), .ZN(new_n1181_));
  NOR2_X1   g1117(.A1(new_n1113_), .A2(new_n1008_), .ZN(new_n1182_));
  NOR2_X1   g1118(.A1(new_n1181_), .A2(new_n1182_), .ZN(new_n1183_));
  INV_X1    g1119(.A(new_n1183_), .ZN(new_n1184_));
  NAND2_X1  g1120(.A1(new_n1111_), .A2(new_n1106_), .ZN(new_n1185_));
  NOR2_X1   g1121(.A1(new_n1098_), .A2(new_n1099_), .ZN(new_n1186_));
  NOR2_X1   g1122(.A1(new_n1103_), .A2(new_n1013_), .ZN(new_n1187_));
  NOR2_X1   g1123(.A1(new_n1186_), .A2(new_n1187_), .ZN(new_n1188_));
  INV_X1    g1124(.A(new_n1188_), .ZN(new_n1189_));
  NAND2_X1  g1125(.A1(new_n1101_), .A2(new_n1096_), .ZN(new_n1190_));
  NOR2_X1   g1126(.A1(new_n1088_), .A2(new_n1089_), .ZN(new_n1191_));
  NOR2_X1   g1127(.A1(new_n1093_), .A2(new_n1018_), .ZN(new_n1192_));
  NOR2_X1   g1128(.A1(new_n1191_), .A2(new_n1192_), .ZN(new_n1193_));
  INV_X1    g1129(.A(new_n1193_), .ZN(new_n1194_));
  NAND2_X1  g1130(.A1(new_n1091_), .A2(new_n1086_), .ZN(new_n1195_));
  NOR2_X1   g1131(.A1(new_n1078_), .A2(new_n1079_), .ZN(new_n1196_));
  NOR2_X1   g1132(.A1(new_n1083_), .A2(new_n1023_), .ZN(new_n1197_));
  NOR2_X1   g1133(.A1(new_n1196_), .A2(new_n1197_), .ZN(new_n1198_));
  INV_X1    g1134(.A(new_n1198_), .ZN(new_n1199_));
  NAND2_X1  g1135(.A1(new_n1081_), .A2(new_n1076_), .ZN(new_n1200_));
  NOR2_X1   g1136(.A1(new_n1068_), .A2(new_n1069_), .ZN(new_n1201_));
  NOR2_X1   g1137(.A1(new_n1073_), .A2(new_n1028_), .ZN(new_n1202_));
  NOR2_X1   g1138(.A1(new_n1201_), .A2(new_n1202_), .ZN(new_n1203_));
  INV_X1    g1139(.A(new_n1203_), .ZN(new_n1204_));
  NAND2_X1  g1140(.A1(new_n1071_), .A2(new_n1066_), .ZN(new_n1205_));
  NOR2_X1   g1141(.A1(new_n1058_), .A2(new_n1057_), .ZN(new_n1206_));
  NOR2_X1   g1142(.A1(new_n1063_), .A2(new_n1031_), .ZN(new_n1207_));
  NOR2_X1   g1143(.A1(new_n1206_), .A2(new_n1207_), .ZN(new_n1208_));
  INV_X1    g1144(.A(new_n1208_), .ZN(new_n1209_));
  NAND2_X1  g1145(.A1(new_n1060_), .A2(new_n1034_), .ZN(new_n1210_));
  AOI22_X1  g1146(.A1(new_n1053_), .A2(new_n1052_), .B1(new_n1045_), .B2(new_n1048_), .ZN(new_n1211_));
  INV_X1    g1147(.A(new_n1211_), .ZN(new_n1212_));
  OAI21_X1  g1148(.A(new_n1035_), .B1(new_n1039_), .B2(new_n1044_), .ZN(new_n1213_));
  AOI21_X1  g1149(.A(new_n869_), .B1(new_n1042_), .B2(new_n1043_), .ZN(new_n1214_));
  INV_X1    g1150(.A(new_n1214_), .ZN(new_n1215_));
  AND4_X1   g1151(.A1(G222gat), .A2(G239gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1216_));
  AOI22_X1  g1152(.A1(G222gat), .A2(G290gat), .B1(G239gat), .B2(G273gat), .ZN(new_n1217_));
  OAI21_X1  g1153(.A(new_n1037_), .B1(new_n1216_), .B2(new_n1217_), .ZN(new_n1218_));
  NAND2_X1  g1154(.A1(G222gat), .A2(G290gat), .ZN(new_n1219_));
  INV_X1    g1155(.A(G239gat), .ZN(new_n1220_));
  OAI21_X1  g1156(.A(new_n1219_), .B1(new_n1220_), .B2(new_n66_), .ZN(new_n1221_));
  NAND4_X1  g1157(.A1(G222gat), .A2(G239gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1222_));
  NAND3_X1  g1158(.A1(new_n1221_), .A2(new_n1043_), .A3(new_n1222_), .ZN(new_n1223_));
  NAND2_X1  g1159(.A1(G205gat), .A2(G307gat), .ZN(new_n1224_));
  AND3_X1   g1160(.A1(new_n1218_), .A2(new_n1223_), .A3(new_n1224_), .ZN(new_n1225_));
  AOI21_X1  g1161(.A(new_n1224_), .B1(new_n1218_), .B2(new_n1223_), .ZN(new_n1226_));
  OAI211_X1 g1162(.A(new_n1213_), .B(new_n1215_), .C1(new_n1225_), .C2(new_n1226_), .ZN(new_n1227_));
  INV_X1    g1163(.A(new_n1224_), .ZN(new_n1228_));
  AND3_X1   g1164(.A1(new_n1221_), .A2(new_n1043_), .A3(new_n1222_), .ZN(new_n1229_));
  AOI21_X1  g1165(.A(new_n1043_), .B1(new_n1221_), .B2(new_n1222_), .ZN(new_n1230_));
  OAI21_X1  g1166(.A(new_n1228_), .B1(new_n1229_), .B2(new_n1230_), .ZN(new_n1231_));
  NAND3_X1  g1167(.A1(new_n1218_), .A2(new_n1223_), .A3(new_n1224_), .ZN(new_n1232_));
  AOI21_X1  g1168(.A(new_n1036_), .B1(new_n1046_), .B2(new_n1047_), .ZN(new_n1233_));
  OAI211_X1 g1169(.A(new_n1231_), .B(new_n1232_), .C1(new_n1233_), .C2(new_n1214_), .ZN(new_n1234_));
  NOR2_X1   g1170(.A1(new_n719_), .A2(new_n130_), .ZN(new_n1235_));
  INV_X1    g1171(.A(new_n1235_), .ZN(new_n1236_));
  NAND3_X1  g1172(.A1(new_n1227_), .A2(new_n1234_), .A3(new_n1236_), .ZN(new_n1237_));
  INV_X1    g1173(.A(new_n1237_), .ZN(new_n1238_));
  AOI21_X1  g1174(.A(new_n1236_), .B1(new_n1227_), .B2(new_n1234_), .ZN(new_n1239_));
  OAI211_X1 g1175(.A(new_n1210_), .B(new_n1212_), .C1(new_n1238_), .C2(new_n1239_), .ZN(new_n1240_));
  NAND2_X1  g1176(.A1(new_n1227_), .A2(new_n1234_), .ZN(new_n1241_));
  NAND2_X1  g1177(.A1(new_n1241_), .A2(new_n1235_), .ZN(new_n1242_));
  AOI21_X1  g1178(.A(new_n1033_), .B1(new_n1051_), .B2(new_n1056_), .ZN(new_n1243_));
  OAI211_X1 g1179(.A(new_n1242_), .B(new_n1237_), .C1(new_n1211_), .C2(new_n1243_), .ZN(new_n1244_));
  NOR2_X1   g1180(.A1(new_n876_), .A2(new_n178_), .ZN(new_n1245_));
  INV_X1    g1181(.A(new_n1245_), .ZN(new_n1246_));
  NAND3_X1  g1182(.A1(new_n1240_), .A2(new_n1244_), .A3(new_n1246_), .ZN(new_n1247_));
  INV_X1    g1183(.A(new_n1247_), .ZN(new_n1248_));
  AOI21_X1  g1184(.A(new_n1246_), .B1(new_n1240_), .B2(new_n1244_), .ZN(new_n1249_));
  OAI211_X1 g1185(.A(new_n1205_), .B(new_n1209_), .C1(new_n1248_), .C2(new_n1249_), .ZN(new_n1250_));
  NAND2_X1  g1186(.A1(new_n1240_), .A2(new_n1244_), .ZN(new_n1251_));
  NAND2_X1  g1187(.A1(new_n1251_), .A2(new_n1245_), .ZN(new_n1252_));
  AOI21_X1  g1188(.A(new_n1065_), .B1(new_n1059_), .B2(new_n1064_), .ZN(new_n1253_));
  OAI211_X1 g1189(.A(new_n1252_), .B(new_n1247_), .C1(new_n1208_), .C2(new_n1253_), .ZN(new_n1254_));
  NOR2_X1   g1190(.A1(new_n889_), .A2(new_n190_), .ZN(new_n1255_));
  INV_X1    g1191(.A(new_n1255_), .ZN(new_n1256_));
  NAND3_X1  g1192(.A1(new_n1250_), .A2(new_n1254_), .A3(new_n1256_), .ZN(new_n1257_));
  INV_X1    g1193(.A(new_n1257_), .ZN(new_n1258_));
  AOI21_X1  g1194(.A(new_n1256_), .B1(new_n1250_), .B2(new_n1254_), .ZN(new_n1259_));
  OAI211_X1 g1195(.A(new_n1200_), .B(new_n1204_), .C1(new_n1258_), .C2(new_n1259_), .ZN(new_n1260_));
  NAND2_X1  g1196(.A1(new_n1250_), .A2(new_n1254_), .ZN(new_n1261_));
  NAND2_X1  g1197(.A1(new_n1261_), .A2(new_n1255_), .ZN(new_n1262_));
  AOI21_X1  g1198(.A(new_n1075_), .B1(new_n1070_), .B2(new_n1074_), .ZN(new_n1263_));
  OAI211_X1 g1199(.A(new_n1262_), .B(new_n1257_), .C1(new_n1263_), .C2(new_n1203_), .ZN(new_n1264_));
  NOR2_X1   g1200(.A1(new_n733_), .A2(new_n253_), .ZN(new_n1265_));
  INV_X1    g1201(.A(new_n1265_), .ZN(new_n1266_));
  NAND3_X1  g1202(.A1(new_n1260_), .A2(new_n1264_), .A3(new_n1266_), .ZN(new_n1267_));
  INV_X1    g1203(.A(new_n1267_), .ZN(new_n1268_));
  AOI21_X1  g1204(.A(new_n1266_), .B1(new_n1260_), .B2(new_n1264_), .ZN(new_n1269_));
  OAI211_X1 g1205(.A(new_n1195_), .B(new_n1199_), .C1(new_n1268_), .C2(new_n1269_), .ZN(new_n1270_));
  NAND2_X1  g1206(.A1(new_n1260_), .A2(new_n1264_), .ZN(new_n1271_));
  NAND2_X1  g1207(.A1(new_n1271_), .A2(new_n1265_), .ZN(new_n1272_));
  AOI21_X1  g1208(.A(new_n1085_), .B1(new_n1080_), .B2(new_n1084_), .ZN(new_n1273_));
  OAI211_X1 g1209(.A(new_n1272_), .B(new_n1267_), .C1(new_n1273_), .C2(new_n1198_), .ZN(new_n1274_));
  NOR2_X1   g1210(.A1(new_n276_), .A2(new_n336_), .ZN(new_n1275_));
  INV_X1    g1211(.A(new_n1275_), .ZN(new_n1276_));
  NAND3_X1  g1212(.A1(new_n1270_), .A2(new_n1274_), .A3(new_n1276_), .ZN(new_n1277_));
  INV_X1    g1213(.A(new_n1277_), .ZN(new_n1278_));
  AOI21_X1  g1214(.A(new_n1276_), .B1(new_n1270_), .B2(new_n1274_), .ZN(new_n1279_));
  OAI211_X1 g1215(.A(new_n1190_), .B(new_n1194_), .C1(new_n1278_), .C2(new_n1279_), .ZN(new_n1280_));
  NAND2_X1  g1216(.A1(new_n1270_), .A2(new_n1274_), .ZN(new_n1281_));
  NAND2_X1  g1217(.A1(new_n1281_), .A2(new_n1275_), .ZN(new_n1282_));
  AOI21_X1  g1218(.A(new_n1095_), .B1(new_n1090_), .B2(new_n1094_), .ZN(new_n1283_));
  OAI211_X1 g1219(.A(new_n1282_), .B(new_n1277_), .C1(new_n1283_), .C2(new_n1193_), .ZN(new_n1284_));
  NOR2_X1   g1220(.A1(new_n205_), .A2(new_n432_), .ZN(new_n1285_));
  INV_X1    g1221(.A(new_n1285_), .ZN(new_n1286_));
  NAND3_X1  g1222(.A1(new_n1280_), .A2(new_n1284_), .A3(new_n1286_), .ZN(new_n1287_));
  INV_X1    g1223(.A(new_n1287_), .ZN(new_n1288_));
  AOI21_X1  g1224(.A(new_n1286_), .B1(new_n1280_), .B2(new_n1284_), .ZN(new_n1289_));
  OAI211_X1 g1225(.A(new_n1185_), .B(new_n1189_), .C1(new_n1288_), .C2(new_n1289_), .ZN(new_n1290_));
  NAND2_X1  g1226(.A1(new_n1280_), .A2(new_n1284_), .ZN(new_n1291_));
  NAND2_X1  g1227(.A1(new_n1291_), .A2(new_n1285_), .ZN(new_n1292_));
  AOI21_X1  g1228(.A(new_n1105_), .B1(new_n1100_), .B2(new_n1104_), .ZN(new_n1293_));
  OAI211_X1 g1229(.A(new_n1292_), .B(new_n1287_), .C1(new_n1293_), .C2(new_n1188_), .ZN(new_n1294_));
  NOR2_X1   g1230(.A1(new_n146_), .A2(new_n544_), .ZN(new_n1295_));
  INV_X1    g1231(.A(new_n1295_), .ZN(new_n1296_));
  NAND3_X1  g1232(.A1(new_n1290_), .A2(new_n1294_), .A3(new_n1296_), .ZN(new_n1297_));
  INV_X1    g1233(.A(new_n1297_), .ZN(new_n1298_));
  AOI21_X1  g1234(.A(new_n1296_), .B1(new_n1290_), .B2(new_n1294_), .ZN(new_n1299_));
  OAI211_X1 g1235(.A(new_n1180_), .B(new_n1184_), .C1(new_n1298_), .C2(new_n1299_), .ZN(new_n1300_));
  NAND2_X1  g1236(.A1(new_n1290_), .A2(new_n1294_), .ZN(new_n1301_));
  NAND2_X1  g1237(.A1(new_n1301_), .A2(new_n1295_), .ZN(new_n1302_));
  AOI21_X1  g1238(.A(new_n1115_), .B1(new_n1110_), .B2(new_n1114_), .ZN(new_n1303_));
  OAI211_X1 g1239(.A(new_n1302_), .B(new_n1297_), .C1(new_n1303_), .C2(new_n1183_), .ZN(new_n1304_));
  NOR2_X1   g1240(.A1(new_n113_), .A2(new_n673_), .ZN(new_n1305_));
  INV_X1    g1241(.A(new_n1305_), .ZN(new_n1306_));
  NAND3_X1  g1242(.A1(new_n1300_), .A2(new_n1304_), .A3(new_n1306_), .ZN(new_n1307_));
  INV_X1    g1243(.A(new_n1307_), .ZN(new_n1308_));
  AOI21_X1  g1244(.A(new_n1306_), .B1(new_n1300_), .B2(new_n1304_), .ZN(new_n1309_));
  OAI211_X1 g1245(.A(new_n1175_), .B(new_n1179_), .C1(new_n1308_), .C2(new_n1309_), .ZN(new_n1310_));
  NAND2_X1  g1246(.A1(new_n1300_), .A2(new_n1304_), .ZN(new_n1311_));
  NAND2_X1  g1247(.A1(new_n1311_), .A2(new_n1305_), .ZN(new_n1312_));
  AOI21_X1  g1248(.A(new_n1125_), .B1(new_n1120_), .B2(new_n1124_), .ZN(new_n1313_));
  OAI211_X1 g1249(.A(new_n1312_), .B(new_n1307_), .C1(new_n1313_), .C2(new_n1178_), .ZN(new_n1314_));
  NOR2_X1   g1250(.A1(new_n86_), .A2(new_n816_), .ZN(new_n1315_));
  INV_X1    g1251(.A(new_n1315_), .ZN(new_n1316_));
  NAND3_X1  g1252(.A1(new_n1310_), .A2(new_n1314_), .A3(new_n1316_), .ZN(new_n1317_));
  INV_X1    g1253(.A(new_n1317_), .ZN(new_n1318_));
  AOI21_X1  g1254(.A(new_n1316_), .B1(new_n1310_), .B2(new_n1314_), .ZN(new_n1319_));
  OAI211_X1 g1255(.A(new_n1170_), .B(new_n1174_), .C1(new_n1318_), .C2(new_n1319_), .ZN(new_n1320_));
  NAND2_X1  g1256(.A1(new_n1310_), .A2(new_n1314_), .ZN(new_n1321_));
  NAND2_X1  g1257(.A1(new_n1321_), .A2(new_n1315_), .ZN(new_n1322_));
  AOI21_X1  g1258(.A(new_n1135_), .B1(new_n1130_), .B2(new_n1134_), .ZN(new_n1323_));
  OAI211_X1 g1259(.A(new_n1322_), .B(new_n1317_), .C1(new_n1323_), .C2(new_n1173_), .ZN(new_n1324_));
  NOR2_X1   g1260(.A1(new_n76_), .A2(new_n980_), .ZN(new_n1325_));
  INV_X1    g1261(.A(new_n1325_), .ZN(new_n1326_));
  NAND3_X1  g1262(.A1(new_n1320_), .A2(new_n1324_), .A3(new_n1326_), .ZN(new_n1327_));
  INV_X1    g1263(.A(new_n1327_), .ZN(new_n1328_));
  AOI21_X1  g1264(.A(new_n1326_), .B1(new_n1320_), .B2(new_n1324_), .ZN(new_n1329_));
  OAI211_X1 g1265(.A(new_n1165_), .B(new_n1169_), .C1(new_n1328_), .C2(new_n1329_), .ZN(new_n1330_));
  NAND2_X1  g1266(.A1(new_n1320_), .A2(new_n1324_), .ZN(new_n1331_));
  NAND2_X1  g1267(.A1(new_n1331_), .A2(new_n1325_), .ZN(new_n1332_));
  AOI21_X1  g1268(.A(new_n1145_), .B1(new_n1140_), .B2(new_n1144_), .ZN(new_n1333_));
  OAI211_X1 g1269(.A(new_n1332_), .B(new_n1327_), .C1(new_n1333_), .C2(new_n1168_), .ZN(new_n1334_));
  NOR2_X1   g1270(.A1(new_n68_), .A2(new_n1155_), .ZN(new_n1335_));
  INV_X1    g1271(.A(new_n1335_), .ZN(new_n1336_));
  NAND3_X1  g1272(.A1(new_n1330_), .A2(new_n1334_), .A3(new_n1336_), .ZN(new_n1337_));
  INV_X1    g1273(.A(new_n1337_), .ZN(new_n1338_));
  AOI21_X1  g1274(.A(new_n1336_), .B1(new_n1330_), .B2(new_n1334_), .ZN(new_n1339_));
  OAI211_X1 g1275(.A(new_n1159_), .B(new_n1163_), .C1(new_n1338_), .C2(new_n1339_), .ZN(new_n1340_));
  INV_X1    g1276(.A(new_n1339_), .ZN(new_n1341_));
  AOI21_X1  g1277(.A(new_n1156_), .B1(new_n1150_), .B2(new_n1153_), .ZN(new_n1342_));
  OAI211_X1 g1278(.A(new_n1341_), .B(new_n1337_), .C1(new_n1342_), .C2(new_n1162_), .ZN(new_n1343_));
  NAND2_X1  g1279(.A1(new_n1340_), .A2(new_n1343_), .ZN(new_n1344_));
  INV_X1    g1280(.A(G511gat), .ZN(new_n1345_));
  NOR2_X1   g1281(.A1(new_n65_), .A2(new_n1345_), .ZN(new_n1346_));
  INV_X1    g1282(.A(new_n1346_), .ZN(new_n1347_));
  XNOR2_X1  g1283(.A(new_n1344_), .B(new_n1347_), .ZN(G5971gat));
  NAND2_X1  g1284(.A1(new_n1330_), .A2(new_n1334_), .ZN(new_n1349_));
  NAND2_X1  g1285(.A1(new_n1349_), .A2(new_n1336_), .ZN(new_n1350_));
  NOR2_X1   g1286(.A1(new_n1328_), .A2(new_n1329_), .ZN(new_n1351_));
  NOR2_X1   g1287(.A1(new_n1333_), .A2(new_n1168_), .ZN(new_n1352_));
  NOR2_X1   g1288(.A1(new_n1351_), .A2(new_n1352_), .ZN(new_n1353_));
  INV_X1    g1289(.A(new_n1353_), .ZN(new_n1354_));
  NAND2_X1  g1290(.A1(new_n1331_), .A2(new_n1326_), .ZN(new_n1355_));
  NOR2_X1   g1291(.A1(new_n1318_), .A2(new_n1319_), .ZN(new_n1356_));
  NOR2_X1   g1292(.A1(new_n1323_), .A2(new_n1173_), .ZN(new_n1357_));
  NOR2_X1   g1293(.A1(new_n1356_), .A2(new_n1357_), .ZN(new_n1358_));
  INV_X1    g1294(.A(new_n1358_), .ZN(new_n1359_));
  NAND2_X1  g1295(.A1(new_n1321_), .A2(new_n1316_), .ZN(new_n1360_));
  NOR2_X1   g1296(.A1(new_n1308_), .A2(new_n1309_), .ZN(new_n1361_));
  NOR2_X1   g1297(.A1(new_n1313_), .A2(new_n1178_), .ZN(new_n1362_));
  NOR2_X1   g1298(.A1(new_n1361_), .A2(new_n1362_), .ZN(new_n1363_));
  INV_X1    g1299(.A(new_n1363_), .ZN(new_n1364_));
  NAND2_X1  g1300(.A1(new_n1311_), .A2(new_n1306_), .ZN(new_n1365_));
  NOR2_X1   g1301(.A1(new_n1298_), .A2(new_n1299_), .ZN(new_n1366_));
  NOR2_X1   g1302(.A1(new_n1303_), .A2(new_n1183_), .ZN(new_n1367_));
  NOR2_X1   g1303(.A1(new_n1366_), .A2(new_n1367_), .ZN(new_n1368_));
  INV_X1    g1304(.A(new_n1368_), .ZN(new_n1369_));
  NAND2_X1  g1305(.A1(new_n1301_), .A2(new_n1296_), .ZN(new_n1370_));
  NOR2_X1   g1306(.A1(new_n1288_), .A2(new_n1289_), .ZN(new_n1371_));
  NOR2_X1   g1307(.A1(new_n1293_), .A2(new_n1188_), .ZN(new_n1372_));
  NOR2_X1   g1308(.A1(new_n1371_), .A2(new_n1372_), .ZN(new_n1373_));
  INV_X1    g1309(.A(new_n1373_), .ZN(new_n1374_));
  NAND2_X1  g1310(.A1(new_n1291_), .A2(new_n1286_), .ZN(new_n1375_));
  NOR2_X1   g1311(.A1(new_n1278_), .A2(new_n1279_), .ZN(new_n1376_));
  NOR2_X1   g1312(.A1(new_n1283_), .A2(new_n1193_), .ZN(new_n1377_));
  NOR2_X1   g1313(.A1(new_n1376_), .A2(new_n1377_), .ZN(new_n1378_));
  INV_X1    g1314(.A(new_n1378_), .ZN(new_n1379_));
  NAND2_X1  g1315(.A1(new_n1281_), .A2(new_n1276_), .ZN(new_n1380_));
  NOR2_X1   g1316(.A1(new_n1268_), .A2(new_n1269_), .ZN(new_n1381_));
  NOR2_X1   g1317(.A1(new_n1273_), .A2(new_n1198_), .ZN(new_n1382_));
  NOR2_X1   g1318(.A1(new_n1381_), .A2(new_n1382_), .ZN(new_n1383_));
  INV_X1    g1319(.A(new_n1383_), .ZN(new_n1384_));
  NAND2_X1  g1320(.A1(new_n1271_), .A2(new_n1266_), .ZN(new_n1385_));
  NOR2_X1   g1321(.A1(new_n1258_), .A2(new_n1259_), .ZN(new_n1386_));
  NOR2_X1   g1322(.A1(new_n1263_), .A2(new_n1203_), .ZN(new_n1387_));
  NOR2_X1   g1323(.A1(new_n1386_), .A2(new_n1387_), .ZN(new_n1388_));
  INV_X1    g1324(.A(new_n1388_), .ZN(new_n1389_));
  NAND2_X1  g1325(.A1(new_n1261_), .A2(new_n1256_), .ZN(new_n1390_));
  NOR2_X1   g1326(.A1(new_n1248_), .A2(new_n1249_), .ZN(new_n1391_));
  NOR2_X1   g1327(.A1(new_n1253_), .A2(new_n1208_), .ZN(new_n1392_));
  NOR2_X1   g1328(.A1(new_n1391_), .A2(new_n1392_), .ZN(new_n1393_));
  INV_X1    g1329(.A(new_n1393_), .ZN(new_n1394_));
  NAND2_X1  g1330(.A1(new_n1251_), .A2(new_n1246_), .ZN(new_n1395_));
  NOR2_X1   g1331(.A1(new_n1238_), .A2(new_n1239_), .ZN(new_n1396_));
  NOR2_X1   g1332(.A1(new_n1243_), .A2(new_n1211_), .ZN(new_n1397_));
  NOR2_X1   g1333(.A1(new_n1396_), .A2(new_n1397_), .ZN(new_n1398_));
  INV_X1    g1334(.A(new_n1398_), .ZN(new_n1399_));
  NAND2_X1  g1335(.A1(new_n1241_), .A2(new_n1236_), .ZN(new_n1400_));
  AOI22_X1  g1336(.A1(new_n1215_), .A2(new_n1213_), .B1(new_n1231_), .B2(new_n1232_), .ZN(new_n1401_));
  INV_X1    g1337(.A(new_n1401_), .ZN(new_n1402_));
  AOI21_X1  g1338(.A(new_n1037_), .B1(new_n1221_), .B2(new_n1222_), .ZN(new_n1403_));
  INV_X1    g1339(.A(new_n1403_), .ZN(new_n1404_));
  OAI21_X1  g1340(.A(new_n1224_), .B1(new_n1229_), .B2(new_n1230_), .ZN(new_n1405_));
  AND4_X1   g1341(.A1(G239gat), .A2(G256gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1406_));
  AOI22_X1  g1342(.A1(G239gat), .A2(G290gat), .B1(G256gat), .B2(G273gat), .ZN(new_n1407_));
  OAI21_X1  g1343(.A(new_n1216_), .B1(new_n1406_), .B2(new_n1407_), .ZN(new_n1408_));
  NAND2_X1  g1344(.A1(G256gat), .A2(G273gat), .ZN(new_n1409_));
  NAND2_X1  g1345(.A1(G239gat), .A2(G290gat), .ZN(new_n1410_));
  NAND2_X1  g1346(.A1(new_n1409_), .A2(new_n1410_), .ZN(new_n1411_));
  NAND4_X1  g1347(.A1(G239gat), .A2(G256gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1412_));
  NAND3_X1  g1348(.A1(new_n1411_), .A2(new_n1222_), .A3(new_n1412_), .ZN(new_n1413_));
  NAND2_X1  g1349(.A1(G222gat), .A2(G307gat), .ZN(new_n1414_));
  AND3_X1   g1350(.A1(new_n1408_), .A2(new_n1413_), .A3(new_n1414_), .ZN(new_n1415_));
  AOI21_X1  g1351(.A(new_n1414_), .B1(new_n1408_), .B2(new_n1413_), .ZN(new_n1416_));
  OAI211_X1 g1352(.A(new_n1404_), .B(new_n1405_), .C1(new_n1415_), .C2(new_n1416_), .ZN(new_n1417_));
  INV_X1    g1353(.A(new_n1414_), .ZN(new_n1418_));
  AND3_X1   g1354(.A1(new_n1411_), .A2(new_n1222_), .A3(new_n1412_), .ZN(new_n1419_));
  AOI21_X1  g1355(.A(new_n1222_), .B1(new_n1411_), .B2(new_n1412_), .ZN(new_n1420_));
  OAI21_X1  g1356(.A(new_n1418_), .B1(new_n1419_), .B2(new_n1420_), .ZN(new_n1421_));
  NAND3_X1  g1357(.A1(new_n1408_), .A2(new_n1413_), .A3(new_n1414_), .ZN(new_n1422_));
  AOI21_X1  g1358(.A(new_n1228_), .B1(new_n1218_), .B2(new_n1223_), .ZN(new_n1423_));
  OAI211_X1 g1359(.A(new_n1421_), .B(new_n1422_), .C1(new_n1423_), .C2(new_n1403_), .ZN(new_n1424_));
  NOR2_X1   g1360(.A1(new_n873_), .A2(new_n130_), .ZN(new_n1425_));
  INV_X1    g1361(.A(new_n1425_), .ZN(new_n1426_));
  NAND3_X1  g1362(.A1(new_n1417_), .A2(new_n1424_), .A3(new_n1426_), .ZN(new_n1427_));
  INV_X1    g1363(.A(new_n1427_), .ZN(new_n1428_));
  AOI21_X1  g1364(.A(new_n1426_), .B1(new_n1417_), .B2(new_n1424_), .ZN(new_n1429_));
  OAI211_X1 g1365(.A(new_n1400_), .B(new_n1402_), .C1(new_n1428_), .C2(new_n1429_), .ZN(new_n1430_));
  NAND2_X1  g1366(.A1(new_n1417_), .A2(new_n1424_), .ZN(new_n1431_));
  NAND2_X1  g1367(.A1(new_n1431_), .A2(new_n1425_), .ZN(new_n1432_));
  AOI21_X1  g1368(.A(new_n1235_), .B1(new_n1227_), .B2(new_n1234_), .ZN(new_n1433_));
  OAI211_X1 g1369(.A(new_n1432_), .B(new_n1427_), .C1(new_n1401_), .C2(new_n1433_), .ZN(new_n1434_));
  NOR2_X1   g1370(.A1(new_n719_), .A2(new_n178_), .ZN(new_n1435_));
  INV_X1    g1371(.A(new_n1435_), .ZN(new_n1436_));
  AND3_X1   g1372(.A1(new_n1430_), .A2(new_n1434_), .A3(new_n1436_), .ZN(new_n1437_));
  AOI21_X1  g1373(.A(new_n1436_), .B1(new_n1430_), .B2(new_n1434_), .ZN(new_n1438_));
  OAI211_X1 g1374(.A(new_n1395_), .B(new_n1399_), .C1(new_n1437_), .C2(new_n1438_), .ZN(new_n1439_));
  NAND2_X1  g1375(.A1(new_n1430_), .A2(new_n1434_), .ZN(new_n1440_));
  NAND2_X1  g1376(.A1(new_n1440_), .A2(new_n1435_), .ZN(new_n1441_));
  NAND3_X1  g1377(.A1(new_n1430_), .A2(new_n1434_), .A3(new_n1436_), .ZN(new_n1442_));
  AOI21_X1  g1378(.A(new_n1245_), .B1(new_n1240_), .B2(new_n1244_), .ZN(new_n1443_));
  OAI211_X1 g1379(.A(new_n1441_), .B(new_n1442_), .C1(new_n1398_), .C2(new_n1443_), .ZN(new_n1444_));
  NOR2_X1   g1380(.A1(new_n876_), .A2(new_n190_), .ZN(new_n1445_));
  INV_X1    g1381(.A(new_n1445_), .ZN(new_n1446_));
  AND3_X1   g1382(.A1(new_n1439_), .A2(new_n1444_), .A3(new_n1446_), .ZN(new_n1447_));
  AOI21_X1  g1383(.A(new_n1446_), .B1(new_n1439_), .B2(new_n1444_), .ZN(new_n1448_));
  OAI211_X1 g1384(.A(new_n1390_), .B(new_n1394_), .C1(new_n1447_), .C2(new_n1448_), .ZN(new_n1449_));
  NAND2_X1  g1385(.A1(new_n1439_), .A2(new_n1444_), .ZN(new_n1450_));
  NAND2_X1  g1386(.A1(new_n1450_), .A2(new_n1445_), .ZN(new_n1451_));
  NAND3_X1  g1387(.A1(new_n1439_), .A2(new_n1444_), .A3(new_n1446_), .ZN(new_n1452_));
  AOI21_X1  g1388(.A(new_n1255_), .B1(new_n1250_), .B2(new_n1254_), .ZN(new_n1453_));
  OAI211_X1 g1389(.A(new_n1451_), .B(new_n1452_), .C1(new_n1393_), .C2(new_n1453_), .ZN(new_n1454_));
  NOR2_X1   g1390(.A1(new_n889_), .A2(new_n253_), .ZN(new_n1455_));
  INV_X1    g1391(.A(new_n1455_), .ZN(new_n1456_));
  AND3_X1   g1392(.A1(new_n1449_), .A2(new_n1454_), .A3(new_n1456_), .ZN(new_n1457_));
  AOI21_X1  g1393(.A(new_n1456_), .B1(new_n1449_), .B2(new_n1454_), .ZN(new_n1458_));
  OAI211_X1 g1394(.A(new_n1385_), .B(new_n1389_), .C1(new_n1457_), .C2(new_n1458_), .ZN(new_n1459_));
  NAND2_X1  g1395(.A1(new_n1449_), .A2(new_n1454_), .ZN(new_n1460_));
  NAND2_X1  g1396(.A1(new_n1460_), .A2(new_n1455_), .ZN(new_n1461_));
  NAND3_X1  g1397(.A1(new_n1449_), .A2(new_n1454_), .A3(new_n1456_), .ZN(new_n1462_));
  AOI21_X1  g1398(.A(new_n1265_), .B1(new_n1260_), .B2(new_n1264_), .ZN(new_n1463_));
  OAI211_X1 g1399(.A(new_n1461_), .B(new_n1462_), .C1(new_n1388_), .C2(new_n1463_), .ZN(new_n1464_));
  NOR2_X1   g1400(.A1(new_n733_), .A2(new_n336_), .ZN(new_n1465_));
  INV_X1    g1401(.A(new_n1465_), .ZN(new_n1466_));
  AND3_X1   g1402(.A1(new_n1459_), .A2(new_n1464_), .A3(new_n1466_), .ZN(new_n1467_));
  AOI21_X1  g1403(.A(new_n1466_), .B1(new_n1459_), .B2(new_n1464_), .ZN(new_n1468_));
  OAI211_X1 g1404(.A(new_n1380_), .B(new_n1384_), .C1(new_n1467_), .C2(new_n1468_), .ZN(new_n1469_));
  NAND2_X1  g1405(.A1(new_n1459_), .A2(new_n1464_), .ZN(new_n1470_));
  NAND2_X1  g1406(.A1(new_n1470_), .A2(new_n1465_), .ZN(new_n1471_));
  NAND3_X1  g1407(.A1(new_n1459_), .A2(new_n1464_), .A3(new_n1466_), .ZN(new_n1472_));
  AOI21_X1  g1408(.A(new_n1275_), .B1(new_n1270_), .B2(new_n1274_), .ZN(new_n1473_));
  OAI211_X1 g1409(.A(new_n1471_), .B(new_n1472_), .C1(new_n1383_), .C2(new_n1473_), .ZN(new_n1474_));
  NOR2_X1   g1410(.A1(new_n276_), .A2(new_n432_), .ZN(new_n1475_));
  INV_X1    g1411(.A(new_n1475_), .ZN(new_n1476_));
  AND3_X1   g1412(.A1(new_n1469_), .A2(new_n1474_), .A3(new_n1476_), .ZN(new_n1477_));
  AOI21_X1  g1413(.A(new_n1476_), .B1(new_n1469_), .B2(new_n1474_), .ZN(new_n1478_));
  OAI211_X1 g1414(.A(new_n1375_), .B(new_n1379_), .C1(new_n1477_), .C2(new_n1478_), .ZN(new_n1479_));
  NAND2_X1  g1415(.A1(new_n1469_), .A2(new_n1474_), .ZN(new_n1480_));
  NAND2_X1  g1416(.A1(new_n1480_), .A2(new_n1475_), .ZN(new_n1481_));
  NAND3_X1  g1417(.A1(new_n1469_), .A2(new_n1474_), .A3(new_n1476_), .ZN(new_n1482_));
  AOI21_X1  g1418(.A(new_n1285_), .B1(new_n1280_), .B2(new_n1284_), .ZN(new_n1483_));
  OAI211_X1 g1419(.A(new_n1481_), .B(new_n1482_), .C1(new_n1378_), .C2(new_n1483_), .ZN(new_n1484_));
  NOR2_X1   g1420(.A1(new_n205_), .A2(new_n544_), .ZN(new_n1485_));
  INV_X1    g1421(.A(new_n1485_), .ZN(new_n1486_));
  AND3_X1   g1422(.A1(new_n1479_), .A2(new_n1484_), .A3(new_n1486_), .ZN(new_n1487_));
  AOI21_X1  g1423(.A(new_n1486_), .B1(new_n1479_), .B2(new_n1484_), .ZN(new_n1488_));
  OAI211_X1 g1424(.A(new_n1370_), .B(new_n1374_), .C1(new_n1487_), .C2(new_n1488_), .ZN(new_n1489_));
  NAND2_X1  g1425(.A1(new_n1479_), .A2(new_n1484_), .ZN(new_n1490_));
  NAND2_X1  g1426(.A1(new_n1490_), .A2(new_n1485_), .ZN(new_n1491_));
  NAND3_X1  g1427(.A1(new_n1479_), .A2(new_n1484_), .A3(new_n1486_), .ZN(new_n1492_));
  AOI21_X1  g1428(.A(new_n1295_), .B1(new_n1290_), .B2(new_n1294_), .ZN(new_n1493_));
  OAI211_X1 g1429(.A(new_n1491_), .B(new_n1492_), .C1(new_n1373_), .C2(new_n1493_), .ZN(new_n1494_));
  NOR2_X1   g1430(.A1(new_n146_), .A2(new_n673_), .ZN(new_n1495_));
  INV_X1    g1431(.A(new_n1495_), .ZN(new_n1496_));
  AND3_X1   g1432(.A1(new_n1489_), .A2(new_n1494_), .A3(new_n1496_), .ZN(new_n1497_));
  AOI21_X1  g1433(.A(new_n1496_), .B1(new_n1489_), .B2(new_n1494_), .ZN(new_n1498_));
  OAI211_X1 g1434(.A(new_n1365_), .B(new_n1369_), .C1(new_n1497_), .C2(new_n1498_), .ZN(new_n1499_));
  NAND2_X1  g1435(.A1(new_n1489_), .A2(new_n1494_), .ZN(new_n1500_));
  NAND2_X1  g1436(.A1(new_n1500_), .A2(new_n1495_), .ZN(new_n1501_));
  NAND3_X1  g1437(.A1(new_n1489_), .A2(new_n1494_), .A3(new_n1496_), .ZN(new_n1502_));
  AOI21_X1  g1438(.A(new_n1305_), .B1(new_n1300_), .B2(new_n1304_), .ZN(new_n1503_));
  OAI211_X1 g1439(.A(new_n1501_), .B(new_n1502_), .C1(new_n1368_), .C2(new_n1503_), .ZN(new_n1504_));
  NOR2_X1   g1440(.A1(new_n113_), .A2(new_n816_), .ZN(new_n1505_));
  INV_X1    g1441(.A(new_n1505_), .ZN(new_n1506_));
  AND3_X1   g1442(.A1(new_n1499_), .A2(new_n1504_), .A3(new_n1506_), .ZN(new_n1507_));
  AOI21_X1  g1443(.A(new_n1506_), .B1(new_n1499_), .B2(new_n1504_), .ZN(new_n1508_));
  OAI211_X1 g1444(.A(new_n1360_), .B(new_n1364_), .C1(new_n1507_), .C2(new_n1508_), .ZN(new_n1509_));
  NAND2_X1  g1445(.A1(new_n1499_), .A2(new_n1504_), .ZN(new_n1510_));
  NAND2_X1  g1446(.A1(new_n1510_), .A2(new_n1505_), .ZN(new_n1511_));
  NAND3_X1  g1447(.A1(new_n1499_), .A2(new_n1504_), .A3(new_n1506_), .ZN(new_n1512_));
  AOI21_X1  g1448(.A(new_n1315_), .B1(new_n1310_), .B2(new_n1314_), .ZN(new_n1513_));
  OAI211_X1 g1449(.A(new_n1511_), .B(new_n1512_), .C1(new_n1363_), .C2(new_n1513_), .ZN(new_n1514_));
  NOR2_X1   g1450(.A1(new_n86_), .A2(new_n980_), .ZN(new_n1515_));
  INV_X1    g1451(.A(new_n1515_), .ZN(new_n1516_));
  AND3_X1   g1452(.A1(new_n1509_), .A2(new_n1514_), .A3(new_n1516_), .ZN(new_n1517_));
  AOI21_X1  g1453(.A(new_n1516_), .B1(new_n1509_), .B2(new_n1514_), .ZN(new_n1518_));
  OAI211_X1 g1454(.A(new_n1355_), .B(new_n1359_), .C1(new_n1517_), .C2(new_n1518_), .ZN(new_n1519_));
  NAND2_X1  g1455(.A1(new_n1509_), .A2(new_n1514_), .ZN(new_n1520_));
  NAND2_X1  g1456(.A1(new_n1520_), .A2(new_n1515_), .ZN(new_n1521_));
  NAND3_X1  g1457(.A1(new_n1509_), .A2(new_n1514_), .A3(new_n1516_), .ZN(new_n1522_));
  AOI21_X1  g1458(.A(new_n1325_), .B1(new_n1320_), .B2(new_n1324_), .ZN(new_n1523_));
  OAI211_X1 g1459(.A(new_n1521_), .B(new_n1522_), .C1(new_n1358_), .C2(new_n1523_), .ZN(new_n1524_));
  NOR2_X1   g1460(.A1(new_n76_), .A2(new_n1155_), .ZN(new_n1525_));
  INV_X1    g1461(.A(new_n1525_), .ZN(new_n1526_));
  NAND3_X1  g1462(.A1(new_n1519_), .A2(new_n1524_), .A3(new_n1526_), .ZN(new_n1527_));
  INV_X1    g1463(.A(new_n1527_), .ZN(new_n1528_));
  AOI21_X1  g1464(.A(new_n1526_), .B1(new_n1519_), .B2(new_n1524_), .ZN(new_n1529_));
  OAI211_X1 g1465(.A(new_n1350_), .B(new_n1354_), .C1(new_n1528_), .C2(new_n1529_), .ZN(new_n1530_));
  NAND2_X1  g1466(.A1(new_n1519_), .A2(new_n1524_), .ZN(new_n1531_));
  NAND2_X1  g1467(.A1(new_n1531_), .A2(new_n1525_), .ZN(new_n1532_));
  AOI21_X1  g1468(.A(new_n1335_), .B1(new_n1330_), .B2(new_n1334_), .ZN(new_n1533_));
  OAI211_X1 g1469(.A(new_n1532_), .B(new_n1527_), .C1(new_n1353_), .C2(new_n1533_), .ZN(new_n1534_));
  NAND2_X1  g1470(.A1(new_n1530_), .A2(new_n1534_), .ZN(new_n1535_));
  NOR2_X1   g1471(.A1(new_n68_), .A2(new_n1345_), .ZN(new_n1536_));
  NAND2_X1  g1472(.A1(new_n1535_), .A2(new_n1536_), .ZN(new_n1537_));
  INV_X1    g1473(.A(new_n1536_), .ZN(new_n1538_));
  NAND3_X1  g1474(.A1(new_n1530_), .A2(new_n1534_), .A3(new_n1538_), .ZN(new_n1539_));
  NAND2_X1  g1475(.A1(new_n1537_), .A2(new_n1539_), .ZN(new_n1540_));
  NOR2_X1   g1476(.A1(new_n1342_), .A2(new_n1162_), .ZN(new_n1541_));
  NOR2_X1   g1477(.A1(new_n1338_), .A2(new_n1339_), .ZN(new_n1542_));
  NOR2_X1   g1478(.A1(new_n1541_), .A2(new_n1542_), .ZN(new_n1543_));
  INV_X1    g1479(.A(new_n1543_), .ZN(new_n1544_));
  NAND2_X1  g1480(.A1(new_n1344_), .A2(new_n1347_), .ZN(new_n1545_));
  NAND3_X1  g1481(.A1(new_n1540_), .A2(new_n1544_), .A3(new_n1545_), .ZN(new_n1546_));
  AOI21_X1  g1482(.A(new_n1346_), .B1(new_n1340_), .B2(new_n1343_), .ZN(new_n1547_));
  OAI211_X1 g1483(.A(new_n1537_), .B(new_n1539_), .C1(new_n1547_), .C2(new_n1543_), .ZN(new_n1548_));
  NAND2_X1  g1484(.A1(new_n1546_), .A2(new_n1548_), .ZN(new_n1549_));
  NAND2_X1  g1485(.A1(G1gat), .A2(G528gat), .ZN(new_n1550_));
  XNOR2_X1  g1486(.A(new_n1549_), .B(new_n1550_), .ZN(G6123gat));
  AOI22_X1  g1487(.A1(new_n1545_), .A2(new_n1544_), .B1(new_n1537_), .B2(new_n1539_), .ZN(new_n1552_));
  AOI21_X1  g1488(.A(new_n1552_), .B1(new_n1549_), .B2(new_n1550_), .ZN(new_n1553_));
  NAND2_X1  g1489(.A1(new_n1535_), .A2(new_n1538_), .ZN(new_n1554_));
  NOR2_X1   g1490(.A1(new_n1528_), .A2(new_n1529_), .ZN(new_n1555_));
  NOR2_X1   g1491(.A1(new_n1533_), .A2(new_n1353_), .ZN(new_n1556_));
  NOR2_X1   g1492(.A1(new_n1555_), .A2(new_n1556_), .ZN(new_n1557_));
  INV_X1    g1493(.A(new_n1557_), .ZN(new_n1558_));
  NAND2_X1  g1494(.A1(new_n1531_), .A2(new_n1526_), .ZN(new_n1559_));
  NOR2_X1   g1495(.A1(new_n1517_), .A2(new_n1518_), .ZN(new_n1560_));
  NOR2_X1   g1496(.A1(new_n1523_), .A2(new_n1358_), .ZN(new_n1561_));
  NOR2_X1   g1497(.A1(new_n1560_), .A2(new_n1561_), .ZN(new_n1562_));
  INV_X1    g1498(.A(new_n1562_), .ZN(new_n1563_));
  NAND2_X1  g1499(.A1(new_n1520_), .A2(new_n1516_), .ZN(new_n1564_));
  NOR2_X1   g1500(.A1(new_n1507_), .A2(new_n1508_), .ZN(new_n1565_));
  NOR2_X1   g1501(.A1(new_n1513_), .A2(new_n1363_), .ZN(new_n1566_));
  NOR2_X1   g1502(.A1(new_n1565_), .A2(new_n1566_), .ZN(new_n1567_));
  INV_X1    g1503(.A(new_n1567_), .ZN(new_n1568_));
  NAND2_X1  g1504(.A1(new_n1510_), .A2(new_n1506_), .ZN(new_n1569_));
  NOR2_X1   g1505(.A1(new_n1497_), .A2(new_n1498_), .ZN(new_n1570_));
  NOR2_X1   g1506(.A1(new_n1503_), .A2(new_n1368_), .ZN(new_n1571_));
  NOR2_X1   g1507(.A1(new_n1570_), .A2(new_n1571_), .ZN(new_n1572_));
  INV_X1    g1508(.A(new_n1572_), .ZN(new_n1573_));
  NAND2_X1  g1509(.A1(new_n1500_), .A2(new_n1496_), .ZN(new_n1574_));
  NOR2_X1   g1510(.A1(new_n1487_), .A2(new_n1488_), .ZN(new_n1575_));
  NOR2_X1   g1511(.A1(new_n1493_), .A2(new_n1373_), .ZN(new_n1576_));
  NOR2_X1   g1512(.A1(new_n1575_), .A2(new_n1576_), .ZN(new_n1577_));
  INV_X1    g1513(.A(new_n1577_), .ZN(new_n1578_));
  NAND2_X1  g1514(.A1(new_n1490_), .A2(new_n1486_), .ZN(new_n1579_));
  NOR2_X1   g1515(.A1(new_n1477_), .A2(new_n1478_), .ZN(new_n1580_));
  NOR2_X1   g1516(.A1(new_n1483_), .A2(new_n1378_), .ZN(new_n1581_));
  NOR2_X1   g1517(.A1(new_n1580_), .A2(new_n1581_), .ZN(new_n1582_));
  INV_X1    g1518(.A(new_n1582_), .ZN(new_n1583_));
  NAND2_X1  g1519(.A1(new_n1480_), .A2(new_n1476_), .ZN(new_n1584_));
  NOR2_X1   g1520(.A1(new_n1467_), .A2(new_n1468_), .ZN(new_n1585_));
  NOR2_X1   g1521(.A1(new_n1473_), .A2(new_n1383_), .ZN(new_n1586_));
  NOR2_X1   g1522(.A1(new_n1585_), .A2(new_n1586_), .ZN(new_n1587_));
  INV_X1    g1523(.A(new_n1587_), .ZN(new_n1588_));
  NAND2_X1  g1524(.A1(new_n1470_), .A2(new_n1466_), .ZN(new_n1589_));
  NOR2_X1   g1525(.A1(new_n1457_), .A2(new_n1458_), .ZN(new_n1590_));
  NOR2_X1   g1526(.A1(new_n1463_), .A2(new_n1388_), .ZN(new_n1591_));
  NOR2_X1   g1527(.A1(new_n1590_), .A2(new_n1591_), .ZN(new_n1592_));
  INV_X1    g1528(.A(new_n1592_), .ZN(new_n1593_));
  NAND2_X1  g1529(.A1(new_n1460_), .A2(new_n1456_), .ZN(new_n1594_));
  NOR2_X1   g1530(.A1(new_n1447_), .A2(new_n1448_), .ZN(new_n1595_));
  NOR2_X1   g1531(.A1(new_n1453_), .A2(new_n1393_), .ZN(new_n1596_));
  NOR2_X1   g1532(.A1(new_n1595_), .A2(new_n1596_), .ZN(new_n1597_));
  INV_X1    g1533(.A(new_n1597_), .ZN(new_n1598_));
  NAND2_X1  g1534(.A1(new_n1450_), .A2(new_n1446_), .ZN(new_n1599_));
  NOR2_X1   g1535(.A1(new_n1437_), .A2(new_n1438_), .ZN(new_n1600_));
  NOR2_X1   g1536(.A1(new_n1443_), .A2(new_n1398_), .ZN(new_n1601_));
  NOR2_X1   g1537(.A1(new_n1600_), .A2(new_n1601_), .ZN(new_n1602_));
  INV_X1    g1538(.A(new_n1602_), .ZN(new_n1603_));
  NAND2_X1  g1539(.A1(new_n1440_), .A2(new_n1436_), .ZN(new_n1604_));
  NAND2_X1  g1540(.A1(new_n1400_), .A2(new_n1402_), .ZN(new_n1605_));
  OAI21_X1  g1541(.A(new_n1605_), .B1(new_n1429_), .B2(new_n1428_), .ZN(new_n1606_));
  NOR2_X1   g1542(.A1(new_n873_), .A2(new_n178_), .ZN(new_n1607_));
  INV_X1    g1543(.A(new_n1607_), .ZN(new_n1608_));
  AOI22_X1  g1544(.A1(new_n1404_), .A2(new_n1405_), .B1(new_n1421_), .B2(new_n1422_), .ZN(new_n1609_));
  AOI21_X1  g1545(.A(new_n1609_), .B1(new_n1431_), .B2(new_n1426_), .ZN(new_n1610_));
  NOR2_X1   g1546(.A1(new_n1041_), .A2(new_n130_), .ZN(new_n1611_));
  AOI21_X1  g1547(.A(new_n1418_), .B1(new_n1408_), .B2(new_n1413_), .ZN(new_n1612_));
  OAI211_X1 g1548(.A(G256gat), .B(G290gat), .C1(new_n1220_), .C2(new_n66_), .ZN(new_n1613_));
  NAND2_X1  g1549(.A1(G239gat), .A2(G307gat), .ZN(new_n1614_));
  INV_X1    g1550(.A(new_n1614_), .ZN(new_n1615_));
  XNOR2_X1  g1551(.A(new_n1613_), .B(new_n1615_), .ZN(new_n1616_));
  AOI21_X1  g1552(.A(new_n1216_), .B1(new_n1412_), .B2(new_n1411_), .ZN(new_n1617_));
  NOR3_X1   g1553(.A1(new_n1612_), .A2(new_n1616_), .A3(new_n1617_), .ZN(new_n1618_));
  XNOR2_X1  g1554(.A(new_n1613_), .B(new_n1614_), .ZN(new_n1619_));
  OAI21_X1  g1555(.A(new_n1414_), .B1(new_n1419_), .B2(new_n1420_), .ZN(new_n1620_));
  INV_X1    g1556(.A(new_n1617_), .ZN(new_n1621_));
  AOI21_X1  g1557(.A(new_n1619_), .B1(new_n1620_), .B2(new_n1621_), .ZN(new_n1622_));
  OAI21_X1  g1558(.A(new_n1611_), .B1(new_n1618_), .B2(new_n1622_), .ZN(new_n1623_));
  OAI21_X1  g1559(.A(new_n1616_), .B1(new_n1612_), .B2(new_n1617_), .ZN(new_n1624_));
  NAND3_X1  g1560(.A1(new_n1620_), .A2(new_n1621_), .A3(new_n1619_), .ZN(new_n1625_));
  INV_X1    g1561(.A(new_n1611_), .ZN(new_n1626_));
  NAND3_X1  g1562(.A1(new_n1624_), .A2(new_n1625_), .A3(new_n1626_), .ZN(new_n1627_));
  NAND2_X1  g1563(.A1(new_n1623_), .A2(new_n1627_), .ZN(new_n1628_));
  NAND2_X1  g1564(.A1(new_n1610_), .A2(new_n1628_), .ZN(new_n1629_));
  AOI21_X1  g1565(.A(new_n1425_), .B1(new_n1417_), .B2(new_n1424_), .ZN(new_n1630_));
  OAI211_X1 g1566(.A(new_n1623_), .B(new_n1627_), .C1(new_n1630_), .C2(new_n1609_), .ZN(new_n1631_));
  AOI21_X1  g1567(.A(new_n1608_), .B1(new_n1629_), .B2(new_n1631_), .ZN(new_n1632_));
  AND3_X1   g1568(.A1(new_n1629_), .A2(new_n1631_), .A3(new_n1608_), .ZN(new_n1633_));
  OAI211_X1 g1569(.A(new_n1604_), .B(new_n1606_), .C1(new_n1632_), .C2(new_n1633_), .ZN(new_n1634_));
  NAND2_X1  g1570(.A1(new_n1629_), .A2(new_n1631_), .ZN(new_n1635_));
  NAND2_X1  g1571(.A1(new_n1635_), .A2(new_n1607_), .ZN(new_n1636_));
  NAND3_X1  g1572(.A1(new_n1629_), .A2(new_n1631_), .A3(new_n1608_), .ZN(new_n1637_));
  AOI21_X1  g1573(.A(new_n1435_), .B1(new_n1430_), .B2(new_n1434_), .ZN(new_n1638_));
  INV_X1    g1574(.A(new_n1606_), .ZN(new_n1639_));
  OAI211_X1 g1575(.A(new_n1636_), .B(new_n1637_), .C1(new_n1638_), .C2(new_n1639_), .ZN(new_n1640_));
  NOR2_X1   g1576(.A1(new_n719_), .A2(new_n190_), .ZN(new_n1641_));
  INV_X1    g1577(.A(new_n1641_), .ZN(new_n1642_));
  NAND3_X1  g1578(.A1(new_n1634_), .A2(new_n1640_), .A3(new_n1642_), .ZN(new_n1643_));
  INV_X1    g1579(.A(new_n1643_), .ZN(new_n1644_));
  AOI21_X1  g1580(.A(new_n1642_), .B1(new_n1634_), .B2(new_n1640_), .ZN(new_n1645_));
  OAI211_X1 g1581(.A(new_n1599_), .B(new_n1603_), .C1(new_n1644_), .C2(new_n1645_), .ZN(new_n1646_));
  NAND2_X1  g1582(.A1(new_n1634_), .A2(new_n1640_), .ZN(new_n1647_));
  NAND2_X1  g1583(.A1(new_n1647_), .A2(new_n1641_), .ZN(new_n1648_));
  AOI21_X1  g1584(.A(new_n1445_), .B1(new_n1439_), .B2(new_n1444_), .ZN(new_n1649_));
  OAI211_X1 g1585(.A(new_n1648_), .B(new_n1643_), .C1(new_n1649_), .C2(new_n1602_), .ZN(new_n1650_));
  NOR2_X1   g1586(.A1(new_n876_), .A2(new_n253_), .ZN(new_n1651_));
  INV_X1    g1587(.A(new_n1651_), .ZN(new_n1652_));
  AND3_X1   g1588(.A1(new_n1646_), .A2(new_n1650_), .A3(new_n1652_), .ZN(new_n1653_));
  AOI21_X1  g1589(.A(new_n1652_), .B1(new_n1646_), .B2(new_n1650_), .ZN(new_n1654_));
  OAI211_X1 g1590(.A(new_n1594_), .B(new_n1598_), .C1(new_n1653_), .C2(new_n1654_), .ZN(new_n1655_));
  NAND2_X1  g1591(.A1(new_n1646_), .A2(new_n1650_), .ZN(new_n1656_));
  NAND2_X1  g1592(.A1(new_n1656_), .A2(new_n1651_), .ZN(new_n1657_));
  NAND3_X1  g1593(.A1(new_n1646_), .A2(new_n1650_), .A3(new_n1652_), .ZN(new_n1658_));
  AOI21_X1  g1594(.A(new_n1455_), .B1(new_n1449_), .B2(new_n1454_), .ZN(new_n1659_));
  OAI211_X1 g1595(.A(new_n1657_), .B(new_n1658_), .C1(new_n1659_), .C2(new_n1597_), .ZN(new_n1660_));
  NOR2_X1   g1596(.A1(new_n889_), .A2(new_n336_), .ZN(new_n1661_));
  INV_X1    g1597(.A(new_n1661_), .ZN(new_n1662_));
  AND3_X1   g1598(.A1(new_n1655_), .A2(new_n1660_), .A3(new_n1662_), .ZN(new_n1663_));
  AOI21_X1  g1599(.A(new_n1662_), .B1(new_n1655_), .B2(new_n1660_), .ZN(new_n1664_));
  OAI211_X1 g1600(.A(new_n1589_), .B(new_n1593_), .C1(new_n1663_), .C2(new_n1664_), .ZN(new_n1665_));
  NAND2_X1  g1601(.A1(new_n1655_), .A2(new_n1660_), .ZN(new_n1666_));
  NAND2_X1  g1602(.A1(new_n1666_), .A2(new_n1661_), .ZN(new_n1667_));
  NAND3_X1  g1603(.A1(new_n1655_), .A2(new_n1660_), .A3(new_n1662_), .ZN(new_n1668_));
  AOI21_X1  g1604(.A(new_n1465_), .B1(new_n1459_), .B2(new_n1464_), .ZN(new_n1669_));
  OAI211_X1 g1605(.A(new_n1667_), .B(new_n1668_), .C1(new_n1669_), .C2(new_n1592_), .ZN(new_n1670_));
  NOR2_X1   g1606(.A1(new_n733_), .A2(new_n432_), .ZN(new_n1671_));
  INV_X1    g1607(.A(new_n1671_), .ZN(new_n1672_));
  AND3_X1   g1608(.A1(new_n1665_), .A2(new_n1670_), .A3(new_n1672_), .ZN(new_n1673_));
  AOI21_X1  g1609(.A(new_n1672_), .B1(new_n1665_), .B2(new_n1670_), .ZN(new_n1674_));
  OAI211_X1 g1610(.A(new_n1584_), .B(new_n1588_), .C1(new_n1673_), .C2(new_n1674_), .ZN(new_n1675_));
  NAND2_X1  g1611(.A1(new_n1665_), .A2(new_n1670_), .ZN(new_n1676_));
  NAND2_X1  g1612(.A1(new_n1676_), .A2(new_n1671_), .ZN(new_n1677_));
  NAND3_X1  g1613(.A1(new_n1665_), .A2(new_n1670_), .A3(new_n1672_), .ZN(new_n1678_));
  AOI21_X1  g1614(.A(new_n1475_), .B1(new_n1469_), .B2(new_n1474_), .ZN(new_n1679_));
  OAI211_X1 g1615(.A(new_n1677_), .B(new_n1678_), .C1(new_n1679_), .C2(new_n1587_), .ZN(new_n1680_));
  NOR2_X1   g1616(.A1(new_n276_), .A2(new_n544_), .ZN(new_n1681_));
  INV_X1    g1617(.A(new_n1681_), .ZN(new_n1682_));
  AND3_X1   g1618(.A1(new_n1675_), .A2(new_n1680_), .A3(new_n1682_), .ZN(new_n1683_));
  AOI21_X1  g1619(.A(new_n1682_), .B1(new_n1675_), .B2(new_n1680_), .ZN(new_n1684_));
  OAI211_X1 g1620(.A(new_n1579_), .B(new_n1583_), .C1(new_n1683_), .C2(new_n1684_), .ZN(new_n1685_));
  NAND2_X1  g1621(.A1(new_n1675_), .A2(new_n1680_), .ZN(new_n1686_));
  NAND2_X1  g1622(.A1(new_n1686_), .A2(new_n1681_), .ZN(new_n1687_));
  NAND3_X1  g1623(.A1(new_n1675_), .A2(new_n1680_), .A3(new_n1682_), .ZN(new_n1688_));
  AOI21_X1  g1624(.A(new_n1485_), .B1(new_n1479_), .B2(new_n1484_), .ZN(new_n1689_));
  OAI211_X1 g1625(.A(new_n1687_), .B(new_n1688_), .C1(new_n1689_), .C2(new_n1582_), .ZN(new_n1690_));
  NOR2_X1   g1626(.A1(new_n205_), .A2(new_n673_), .ZN(new_n1691_));
  INV_X1    g1627(.A(new_n1691_), .ZN(new_n1692_));
  AND3_X1   g1628(.A1(new_n1685_), .A2(new_n1690_), .A3(new_n1692_), .ZN(new_n1693_));
  AOI21_X1  g1629(.A(new_n1692_), .B1(new_n1685_), .B2(new_n1690_), .ZN(new_n1694_));
  OAI211_X1 g1630(.A(new_n1574_), .B(new_n1578_), .C1(new_n1693_), .C2(new_n1694_), .ZN(new_n1695_));
  NAND2_X1  g1631(.A1(new_n1685_), .A2(new_n1690_), .ZN(new_n1696_));
  NAND2_X1  g1632(.A1(new_n1696_), .A2(new_n1691_), .ZN(new_n1697_));
  NAND3_X1  g1633(.A1(new_n1685_), .A2(new_n1690_), .A3(new_n1692_), .ZN(new_n1698_));
  AOI21_X1  g1634(.A(new_n1495_), .B1(new_n1489_), .B2(new_n1494_), .ZN(new_n1699_));
  OAI211_X1 g1635(.A(new_n1697_), .B(new_n1698_), .C1(new_n1699_), .C2(new_n1577_), .ZN(new_n1700_));
  NOR2_X1   g1636(.A1(new_n146_), .A2(new_n816_), .ZN(new_n1701_));
  INV_X1    g1637(.A(new_n1701_), .ZN(new_n1702_));
  AND3_X1   g1638(.A1(new_n1695_), .A2(new_n1700_), .A3(new_n1702_), .ZN(new_n1703_));
  AOI21_X1  g1639(.A(new_n1702_), .B1(new_n1695_), .B2(new_n1700_), .ZN(new_n1704_));
  OAI211_X1 g1640(.A(new_n1569_), .B(new_n1573_), .C1(new_n1703_), .C2(new_n1704_), .ZN(new_n1705_));
  NAND2_X1  g1641(.A1(new_n1695_), .A2(new_n1700_), .ZN(new_n1706_));
  NAND2_X1  g1642(.A1(new_n1706_), .A2(new_n1701_), .ZN(new_n1707_));
  NAND3_X1  g1643(.A1(new_n1695_), .A2(new_n1700_), .A3(new_n1702_), .ZN(new_n1708_));
  AOI21_X1  g1644(.A(new_n1505_), .B1(new_n1499_), .B2(new_n1504_), .ZN(new_n1709_));
  OAI211_X1 g1645(.A(new_n1707_), .B(new_n1708_), .C1(new_n1709_), .C2(new_n1572_), .ZN(new_n1710_));
  NOR2_X1   g1646(.A1(new_n113_), .A2(new_n980_), .ZN(new_n1711_));
  INV_X1    g1647(.A(new_n1711_), .ZN(new_n1712_));
  AND3_X1   g1648(.A1(new_n1705_), .A2(new_n1710_), .A3(new_n1712_), .ZN(new_n1713_));
  AOI21_X1  g1649(.A(new_n1712_), .B1(new_n1705_), .B2(new_n1710_), .ZN(new_n1714_));
  OAI211_X1 g1650(.A(new_n1564_), .B(new_n1568_), .C1(new_n1713_), .C2(new_n1714_), .ZN(new_n1715_));
  NAND2_X1  g1651(.A1(new_n1705_), .A2(new_n1710_), .ZN(new_n1716_));
  NAND2_X1  g1652(.A1(new_n1716_), .A2(new_n1711_), .ZN(new_n1717_));
  NAND3_X1  g1653(.A1(new_n1705_), .A2(new_n1710_), .A3(new_n1712_), .ZN(new_n1718_));
  AOI21_X1  g1654(.A(new_n1515_), .B1(new_n1509_), .B2(new_n1514_), .ZN(new_n1719_));
  OAI211_X1 g1655(.A(new_n1717_), .B(new_n1718_), .C1(new_n1719_), .C2(new_n1567_), .ZN(new_n1720_));
  NOR2_X1   g1656(.A1(new_n86_), .A2(new_n1155_), .ZN(new_n1721_));
  INV_X1    g1657(.A(new_n1721_), .ZN(new_n1722_));
  AND3_X1   g1658(.A1(new_n1715_), .A2(new_n1720_), .A3(new_n1722_), .ZN(new_n1723_));
  AOI21_X1  g1659(.A(new_n1722_), .B1(new_n1715_), .B2(new_n1720_), .ZN(new_n1724_));
  OAI211_X1 g1660(.A(new_n1559_), .B(new_n1563_), .C1(new_n1723_), .C2(new_n1724_), .ZN(new_n1725_));
  NAND2_X1  g1661(.A1(new_n1715_), .A2(new_n1720_), .ZN(new_n1726_));
  NAND2_X1  g1662(.A1(new_n1726_), .A2(new_n1721_), .ZN(new_n1727_));
  NAND3_X1  g1663(.A1(new_n1715_), .A2(new_n1720_), .A3(new_n1722_), .ZN(new_n1728_));
  AOI21_X1  g1664(.A(new_n1525_), .B1(new_n1519_), .B2(new_n1524_), .ZN(new_n1729_));
  OAI211_X1 g1665(.A(new_n1727_), .B(new_n1728_), .C1(new_n1729_), .C2(new_n1562_), .ZN(new_n1730_));
  NOR2_X1   g1666(.A1(new_n76_), .A2(new_n1345_), .ZN(new_n1731_));
  INV_X1    g1667(.A(new_n1731_), .ZN(new_n1732_));
  NAND3_X1  g1668(.A1(new_n1725_), .A2(new_n1730_), .A3(new_n1732_), .ZN(new_n1733_));
  INV_X1    g1669(.A(new_n1733_), .ZN(new_n1734_));
  AOI21_X1  g1670(.A(new_n1732_), .B1(new_n1725_), .B2(new_n1730_), .ZN(new_n1735_));
  OAI211_X1 g1671(.A(new_n1554_), .B(new_n1558_), .C1(new_n1734_), .C2(new_n1735_), .ZN(new_n1736_));
  NAND2_X1  g1672(.A1(new_n1725_), .A2(new_n1730_), .ZN(new_n1737_));
  NAND2_X1  g1673(.A1(new_n1737_), .A2(new_n1731_), .ZN(new_n1738_));
  AOI21_X1  g1674(.A(new_n1536_), .B1(new_n1530_), .B2(new_n1534_), .ZN(new_n1739_));
  OAI211_X1 g1675(.A(new_n1738_), .B(new_n1733_), .C1(new_n1739_), .C2(new_n1557_), .ZN(new_n1740_));
  INV_X1    g1676(.A(G528gat), .ZN(new_n1741_));
  NOR2_X1   g1677(.A1(new_n68_), .A2(new_n1741_), .ZN(new_n1742_));
  INV_X1    g1678(.A(new_n1742_), .ZN(new_n1743_));
  AND3_X1   g1679(.A1(new_n1736_), .A2(new_n1740_), .A3(new_n1743_), .ZN(new_n1744_));
  AOI21_X1  g1680(.A(new_n1743_), .B1(new_n1736_), .B2(new_n1740_), .ZN(new_n1745_));
  NOR2_X1   g1681(.A1(new_n1744_), .A2(new_n1745_), .ZN(new_n1746_));
  XOR2_X1   g1682(.A(new_n1553_), .B(new_n1746_), .Z(G6150gat));
  NAND2_X1  g1683(.A1(new_n1736_), .A2(new_n1740_), .ZN(new_n1748_));
  NAND2_X1  g1684(.A1(new_n1748_), .A2(new_n1743_), .ZN(new_n1749_));
  NOR2_X1   g1685(.A1(new_n1734_), .A2(new_n1735_), .ZN(new_n1750_));
  NOR2_X1   g1686(.A1(new_n1739_), .A2(new_n1557_), .ZN(new_n1751_));
  NOR2_X1   g1687(.A1(new_n1750_), .A2(new_n1751_), .ZN(new_n1752_));
  INV_X1    g1688(.A(new_n1752_), .ZN(new_n1753_));
  NAND2_X1  g1689(.A1(new_n1737_), .A2(new_n1732_), .ZN(new_n1754_));
  NOR2_X1   g1690(.A1(new_n1723_), .A2(new_n1724_), .ZN(new_n1755_));
  NOR2_X1   g1691(.A1(new_n1729_), .A2(new_n1562_), .ZN(new_n1756_));
  NOR2_X1   g1692(.A1(new_n1755_), .A2(new_n1756_), .ZN(new_n1757_));
  INV_X1    g1693(.A(new_n1757_), .ZN(new_n1758_));
  NAND2_X1  g1694(.A1(new_n1726_), .A2(new_n1722_), .ZN(new_n1759_));
  NOR2_X1   g1695(.A1(new_n1713_), .A2(new_n1714_), .ZN(new_n1760_));
  NOR2_X1   g1696(.A1(new_n1719_), .A2(new_n1567_), .ZN(new_n1761_));
  NOR2_X1   g1697(.A1(new_n1760_), .A2(new_n1761_), .ZN(new_n1762_));
  INV_X1    g1698(.A(new_n1762_), .ZN(new_n1763_));
  NAND2_X1  g1699(.A1(new_n1716_), .A2(new_n1712_), .ZN(new_n1764_));
  NOR2_X1   g1700(.A1(new_n1703_), .A2(new_n1704_), .ZN(new_n1765_));
  NOR2_X1   g1701(.A1(new_n1709_), .A2(new_n1572_), .ZN(new_n1766_));
  NOR2_X1   g1702(.A1(new_n1765_), .A2(new_n1766_), .ZN(new_n1767_));
  INV_X1    g1703(.A(new_n1767_), .ZN(new_n1768_));
  NAND2_X1  g1704(.A1(new_n1706_), .A2(new_n1702_), .ZN(new_n1769_));
  NOR2_X1   g1705(.A1(new_n1693_), .A2(new_n1694_), .ZN(new_n1770_));
  NOR2_X1   g1706(.A1(new_n1699_), .A2(new_n1577_), .ZN(new_n1771_));
  NOR2_X1   g1707(.A1(new_n1770_), .A2(new_n1771_), .ZN(new_n1772_));
  INV_X1    g1708(.A(new_n1772_), .ZN(new_n1773_));
  NAND2_X1  g1709(.A1(new_n1696_), .A2(new_n1692_), .ZN(new_n1774_));
  NOR2_X1   g1710(.A1(new_n1683_), .A2(new_n1684_), .ZN(new_n1775_));
  NOR2_X1   g1711(.A1(new_n1689_), .A2(new_n1582_), .ZN(new_n1776_));
  NOR2_X1   g1712(.A1(new_n1775_), .A2(new_n1776_), .ZN(new_n1777_));
  INV_X1    g1713(.A(new_n1777_), .ZN(new_n1778_));
  NAND2_X1  g1714(.A1(new_n1686_), .A2(new_n1682_), .ZN(new_n1779_));
  NOR2_X1   g1715(.A1(new_n1673_), .A2(new_n1674_), .ZN(new_n1780_));
  NOR2_X1   g1716(.A1(new_n1679_), .A2(new_n1587_), .ZN(new_n1781_));
  NOR2_X1   g1717(.A1(new_n1780_), .A2(new_n1781_), .ZN(new_n1782_));
  INV_X1    g1718(.A(new_n1782_), .ZN(new_n1783_));
  NAND2_X1  g1719(.A1(new_n1676_), .A2(new_n1672_), .ZN(new_n1784_));
  NOR2_X1   g1720(.A1(new_n1663_), .A2(new_n1664_), .ZN(new_n1785_));
  NOR2_X1   g1721(.A1(new_n1669_), .A2(new_n1592_), .ZN(new_n1786_));
  NOR2_X1   g1722(.A1(new_n1785_), .A2(new_n1786_), .ZN(new_n1787_));
  INV_X1    g1723(.A(new_n1787_), .ZN(new_n1788_));
  NAND2_X1  g1724(.A1(new_n1666_), .A2(new_n1662_), .ZN(new_n1789_));
  NOR2_X1   g1725(.A1(new_n1653_), .A2(new_n1654_), .ZN(new_n1790_));
  NOR2_X1   g1726(.A1(new_n1659_), .A2(new_n1597_), .ZN(new_n1791_));
  NOR2_X1   g1727(.A1(new_n1790_), .A2(new_n1791_), .ZN(new_n1792_));
  INV_X1    g1728(.A(new_n1792_), .ZN(new_n1793_));
  NAND2_X1  g1729(.A1(new_n1656_), .A2(new_n1652_), .ZN(new_n1794_));
  NOR2_X1   g1730(.A1(new_n1644_), .A2(new_n1645_), .ZN(new_n1795_));
  NOR2_X1   g1731(.A1(new_n1649_), .A2(new_n1602_), .ZN(new_n1796_));
  NOR2_X1   g1732(.A1(new_n1795_), .A2(new_n1796_), .ZN(new_n1797_));
  INV_X1    g1733(.A(new_n1797_), .ZN(new_n1798_));
  NOR2_X1   g1734(.A1(new_n719_), .A2(new_n253_), .ZN(new_n1799_));
  INV_X1    g1735(.A(new_n1799_), .ZN(new_n1800_));
  AOI22_X1  g1736(.A1(new_n1604_), .A2(new_n1606_), .B1(new_n1636_), .B2(new_n1637_), .ZN(new_n1801_));
  AOI21_X1  g1737(.A(new_n1801_), .B1(new_n1647_), .B2(new_n1642_), .ZN(new_n1802_));
  NAND2_X1  g1738(.A1(new_n1635_), .A2(new_n1608_), .ZN(new_n1803_));
  NOR2_X1   g1739(.A1(new_n1041_), .A2(new_n178_), .ZN(new_n1804_));
  INV_X1    g1740(.A(G256gat), .ZN(new_n1805_));
  OAI21_X1  g1741(.A(new_n1412_), .B1(new_n1805_), .B2(new_n70_), .ZN(new_n1806_));
  NAND2_X1  g1742(.A1(G256gat), .A2(G307gat), .ZN(new_n1807_));
  OAI211_X1 g1743(.A(new_n1806_), .B(new_n1807_), .C1(new_n1613_), .C2(new_n1615_), .ZN(new_n1808_));
  OAI211_X1 g1744(.A(G256gat), .B(G307gat), .C1(new_n1220_), .C2(new_n70_), .ZN(new_n1809_));
  NAND2_X1  g1745(.A1(G239gat), .A2(G324gat), .ZN(new_n1810_));
  AND3_X1   g1746(.A1(new_n1808_), .A2(new_n1809_), .A3(new_n1810_), .ZN(new_n1811_));
  AOI21_X1  g1747(.A(new_n1810_), .B1(new_n1808_), .B2(new_n1809_), .ZN(new_n1812_));
  NOR2_X1   g1748(.A1(new_n1811_), .A2(new_n1812_), .ZN(new_n1813_));
  INV_X1    g1749(.A(new_n1813_), .ZN(new_n1814_));
  OAI21_X1  g1750(.A(new_n1626_), .B1(new_n1618_), .B2(new_n1622_), .ZN(new_n1815_));
  AOI21_X1  g1751(.A(new_n1616_), .B1(new_n1620_), .B2(new_n1621_), .ZN(new_n1816_));
  INV_X1    g1752(.A(new_n1816_), .ZN(new_n1817_));
  AOI21_X1  g1753(.A(new_n1814_), .B1(new_n1815_), .B2(new_n1817_), .ZN(new_n1818_));
  AOI21_X1  g1754(.A(new_n1611_), .B1(new_n1624_), .B2(new_n1625_), .ZN(new_n1819_));
  NOR3_X1   g1755(.A1(new_n1819_), .A2(new_n1816_), .A3(new_n1813_), .ZN(new_n1820_));
  OAI21_X1  g1756(.A(new_n1804_), .B1(new_n1818_), .B2(new_n1820_), .ZN(new_n1821_));
  NAND3_X1  g1757(.A1(new_n1815_), .A2(new_n1817_), .A3(new_n1814_), .ZN(new_n1822_));
  OAI21_X1  g1758(.A(new_n1813_), .B1(new_n1819_), .B2(new_n1816_), .ZN(new_n1823_));
  INV_X1    g1759(.A(new_n1804_), .ZN(new_n1824_));
  NAND3_X1  g1760(.A1(new_n1822_), .A2(new_n1823_), .A3(new_n1824_), .ZN(new_n1825_));
  NAND2_X1  g1761(.A1(new_n1821_), .A2(new_n1825_), .ZN(new_n1826_));
  AOI21_X1  g1762(.A(new_n1610_), .B1(new_n1623_), .B2(new_n1627_), .ZN(new_n1827_));
  INV_X1    g1763(.A(new_n1827_), .ZN(new_n1828_));
  NAND3_X1  g1764(.A1(new_n1803_), .A2(new_n1826_), .A3(new_n1828_), .ZN(new_n1829_));
  AOI21_X1  g1765(.A(new_n1607_), .B1(new_n1629_), .B2(new_n1631_), .ZN(new_n1830_));
  OAI211_X1 g1766(.A(new_n1821_), .B(new_n1825_), .C1(new_n1830_), .C2(new_n1827_), .ZN(new_n1831_));
  NAND2_X1  g1767(.A1(new_n1829_), .A2(new_n1831_), .ZN(new_n1832_));
  NOR2_X1   g1768(.A1(new_n873_), .A2(new_n190_), .ZN(new_n1833_));
  NAND2_X1  g1769(.A1(new_n1832_), .A2(new_n1833_), .ZN(new_n1834_));
  INV_X1    g1770(.A(new_n1833_), .ZN(new_n1835_));
  NAND3_X1  g1771(.A1(new_n1829_), .A2(new_n1831_), .A3(new_n1835_), .ZN(new_n1836_));
  NAND2_X1  g1772(.A1(new_n1834_), .A2(new_n1836_), .ZN(new_n1837_));
  NAND2_X1  g1773(.A1(new_n1802_), .A2(new_n1837_), .ZN(new_n1838_));
  AOI21_X1  g1774(.A(new_n1641_), .B1(new_n1634_), .B2(new_n1640_), .ZN(new_n1839_));
  OAI211_X1 g1775(.A(new_n1834_), .B(new_n1836_), .C1(new_n1839_), .C2(new_n1801_), .ZN(new_n1840_));
  AOI21_X1  g1776(.A(new_n1800_), .B1(new_n1838_), .B2(new_n1840_), .ZN(new_n1841_));
  AND3_X1   g1777(.A1(new_n1838_), .A2(new_n1840_), .A3(new_n1800_), .ZN(new_n1842_));
  OAI211_X1 g1778(.A(new_n1794_), .B(new_n1798_), .C1(new_n1841_), .C2(new_n1842_), .ZN(new_n1843_));
  NAND2_X1  g1779(.A1(new_n1838_), .A2(new_n1840_), .ZN(new_n1844_));
  NAND2_X1  g1780(.A1(new_n1844_), .A2(new_n1799_), .ZN(new_n1845_));
  NAND3_X1  g1781(.A1(new_n1838_), .A2(new_n1840_), .A3(new_n1800_), .ZN(new_n1846_));
  AOI21_X1  g1782(.A(new_n1651_), .B1(new_n1646_), .B2(new_n1650_), .ZN(new_n1847_));
  OAI211_X1 g1783(.A(new_n1845_), .B(new_n1846_), .C1(new_n1847_), .C2(new_n1797_), .ZN(new_n1848_));
  NOR2_X1   g1784(.A1(new_n876_), .A2(new_n336_), .ZN(new_n1849_));
  INV_X1    g1785(.A(new_n1849_), .ZN(new_n1850_));
  NAND3_X1  g1786(.A1(new_n1843_), .A2(new_n1848_), .A3(new_n1850_), .ZN(new_n1851_));
  INV_X1    g1787(.A(new_n1851_), .ZN(new_n1852_));
  AOI21_X1  g1788(.A(new_n1850_), .B1(new_n1843_), .B2(new_n1848_), .ZN(new_n1853_));
  OAI211_X1 g1789(.A(new_n1789_), .B(new_n1793_), .C1(new_n1852_), .C2(new_n1853_), .ZN(new_n1854_));
  NAND2_X1  g1790(.A1(new_n1843_), .A2(new_n1848_), .ZN(new_n1855_));
  NAND2_X1  g1791(.A1(new_n1855_), .A2(new_n1849_), .ZN(new_n1856_));
  AOI21_X1  g1792(.A(new_n1661_), .B1(new_n1655_), .B2(new_n1660_), .ZN(new_n1857_));
  OAI211_X1 g1793(.A(new_n1856_), .B(new_n1851_), .C1(new_n1857_), .C2(new_n1792_), .ZN(new_n1858_));
  NOR2_X1   g1794(.A1(new_n889_), .A2(new_n432_), .ZN(new_n1859_));
  INV_X1    g1795(.A(new_n1859_), .ZN(new_n1860_));
  AND3_X1   g1796(.A1(new_n1854_), .A2(new_n1858_), .A3(new_n1860_), .ZN(new_n1861_));
  AOI21_X1  g1797(.A(new_n1860_), .B1(new_n1854_), .B2(new_n1858_), .ZN(new_n1862_));
  OAI211_X1 g1798(.A(new_n1784_), .B(new_n1788_), .C1(new_n1861_), .C2(new_n1862_), .ZN(new_n1863_));
  NAND2_X1  g1799(.A1(new_n1854_), .A2(new_n1858_), .ZN(new_n1864_));
  NAND2_X1  g1800(.A1(new_n1864_), .A2(new_n1859_), .ZN(new_n1865_));
  NAND3_X1  g1801(.A1(new_n1854_), .A2(new_n1858_), .A3(new_n1860_), .ZN(new_n1866_));
  AOI21_X1  g1802(.A(new_n1671_), .B1(new_n1665_), .B2(new_n1670_), .ZN(new_n1867_));
  OAI211_X1 g1803(.A(new_n1865_), .B(new_n1866_), .C1(new_n1867_), .C2(new_n1787_), .ZN(new_n1868_));
  NOR2_X1   g1804(.A1(new_n733_), .A2(new_n544_), .ZN(new_n1869_));
  INV_X1    g1805(.A(new_n1869_), .ZN(new_n1870_));
  AND3_X1   g1806(.A1(new_n1863_), .A2(new_n1868_), .A3(new_n1870_), .ZN(new_n1871_));
  AOI21_X1  g1807(.A(new_n1870_), .B1(new_n1863_), .B2(new_n1868_), .ZN(new_n1872_));
  OAI211_X1 g1808(.A(new_n1779_), .B(new_n1783_), .C1(new_n1871_), .C2(new_n1872_), .ZN(new_n1873_));
  NAND2_X1  g1809(.A1(new_n1863_), .A2(new_n1868_), .ZN(new_n1874_));
  NAND2_X1  g1810(.A1(new_n1874_), .A2(new_n1869_), .ZN(new_n1875_));
  NAND3_X1  g1811(.A1(new_n1863_), .A2(new_n1868_), .A3(new_n1870_), .ZN(new_n1876_));
  AOI21_X1  g1812(.A(new_n1681_), .B1(new_n1675_), .B2(new_n1680_), .ZN(new_n1877_));
  OAI211_X1 g1813(.A(new_n1875_), .B(new_n1876_), .C1(new_n1877_), .C2(new_n1782_), .ZN(new_n1878_));
  NOR2_X1   g1814(.A1(new_n276_), .A2(new_n673_), .ZN(new_n1879_));
  INV_X1    g1815(.A(new_n1879_), .ZN(new_n1880_));
  AND3_X1   g1816(.A1(new_n1873_), .A2(new_n1878_), .A3(new_n1880_), .ZN(new_n1881_));
  AOI21_X1  g1817(.A(new_n1880_), .B1(new_n1873_), .B2(new_n1878_), .ZN(new_n1882_));
  OAI211_X1 g1818(.A(new_n1774_), .B(new_n1778_), .C1(new_n1881_), .C2(new_n1882_), .ZN(new_n1883_));
  NAND2_X1  g1819(.A1(new_n1873_), .A2(new_n1878_), .ZN(new_n1884_));
  NAND2_X1  g1820(.A1(new_n1884_), .A2(new_n1879_), .ZN(new_n1885_));
  NAND3_X1  g1821(.A1(new_n1873_), .A2(new_n1878_), .A3(new_n1880_), .ZN(new_n1886_));
  AOI21_X1  g1822(.A(new_n1691_), .B1(new_n1685_), .B2(new_n1690_), .ZN(new_n1887_));
  OAI211_X1 g1823(.A(new_n1885_), .B(new_n1886_), .C1(new_n1887_), .C2(new_n1777_), .ZN(new_n1888_));
  NOR2_X1   g1824(.A1(new_n205_), .A2(new_n816_), .ZN(new_n1889_));
  INV_X1    g1825(.A(new_n1889_), .ZN(new_n1890_));
  AND3_X1   g1826(.A1(new_n1883_), .A2(new_n1888_), .A3(new_n1890_), .ZN(new_n1891_));
  AOI21_X1  g1827(.A(new_n1890_), .B1(new_n1883_), .B2(new_n1888_), .ZN(new_n1892_));
  OAI211_X1 g1828(.A(new_n1769_), .B(new_n1773_), .C1(new_n1891_), .C2(new_n1892_), .ZN(new_n1893_));
  NAND2_X1  g1829(.A1(new_n1883_), .A2(new_n1888_), .ZN(new_n1894_));
  NAND2_X1  g1830(.A1(new_n1894_), .A2(new_n1889_), .ZN(new_n1895_));
  NAND3_X1  g1831(.A1(new_n1883_), .A2(new_n1888_), .A3(new_n1890_), .ZN(new_n1896_));
  AOI21_X1  g1832(.A(new_n1701_), .B1(new_n1695_), .B2(new_n1700_), .ZN(new_n1897_));
  OAI211_X1 g1833(.A(new_n1895_), .B(new_n1896_), .C1(new_n1897_), .C2(new_n1772_), .ZN(new_n1898_));
  NOR2_X1   g1834(.A1(new_n146_), .A2(new_n980_), .ZN(new_n1899_));
  INV_X1    g1835(.A(new_n1899_), .ZN(new_n1900_));
  AND3_X1   g1836(.A1(new_n1893_), .A2(new_n1898_), .A3(new_n1900_), .ZN(new_n1901_));
  AOI21_X1  g1837(.A(new_n1900_), .B1(new_n1893_), .B2(new_n1898_), .ZN(new_n1902_));
  OAI211_X1 g1838(.A(new_n1764_), .B(new_n1768_), .C1(new_n1901_), .C2(new_n1902_), .ZN(new_n1903_));
  NAND2_X1  g1839(.A1(new_n1893_), .A2(new_n1898_), .ZN(new_n1904_));
  NAND2_X1  g1840(.A1(new_n1904_), .A2(new_n1899_), .ZN(new_n1905_));
  NAND3_X1  g1841(.A1(new_n1893_), .A2(new_n1898_), .A3(new_n1900_), .ZN(new_n1906_));
  AOI21_X1  g1842(.A(new_n1711_), .B1(new_n1705_), .B2(new_n1710_), .ZN(new_n1907_));
  OAI211_X1 g1843(.A(new_n1905_), .B(new_n1906_), .C1(new_n1907_), .C2(new_n1767_), .ZN(new_n1908_));
  NOR2_X1   g1844(.A1(new_n113_), .A2(new_n1155_), .ZN(new_n1909_));
  INV_X1    g1845(.A(new_n1909_), .ZN(new_n1910_));
  AND3_X1   g1846(.A1(new_n1903_), .A2(new_n1908_), .A3(new_n1910_), .ZN(new_n1911_));
  AOI21_X1  g1847(.A(new_n1910_), .B1(new_n1903_), .B2(new_n1908_), .ZN(new_n1912_));
  OAI211_X1 g1848(.A(new_n1759_), .B(new_n1763_), .C1(new_n1911_), .C2(new_n1912_), .ZN(new_n1913_));
  NAND2_X1  g1849(.A1(new_n1903_), .A2(new_n1908_), .ZN(new_n1914_));
  NAND2_X1  g1850(.A1(new_n1914_), .A2(new_n1909_), .ZN(new_n1915_));
  NAND3_X1  g1851(.A1(new_n1903_), .A2(new_n1908_), .A3(new_n1910_), .ZN(new_n1916_));
  AOI21_X1  g1852(.A(new_n1721_), .B1(new_n1715_), .B2(new_n1720_), .ZN(new_n1917_));
  OAI211_X1 g1853(.A(new_n1915_), .B(new_n1916_), .C1(new_n1917_), .C2(new_n1762_), .ZN(new_n1918_));
  NOR2_X1   g1854(.A1(new_n86_), .A2(new_n1345_), .ZN(new_n1919_));
  INV_X1    g1855(.A(new_n1919_), .ZN(new_n1920_));
  AND3_X1   g1856(.A1(new_n1913_), .A2(new_n1918_), .A3(new_n1920_), .ZN(new_n1921_));
  AOI21_X1  g1857(.A(new_n1920_), .B1(new_n1913_), .B2(new_n1918_), .ZN(new_n1922_));
  OAI211_X1 g1858(.A(new_n1754_), .B(new_n1758_), .C1(new_n1921_), .C2(new_n1922_), .ZN(new_n1923_));
  NAND2_X1  g1859(.A1(new_n1913_), .A2(new_n1918_), .ZN(new_n1924_));
  NAND2_X1  g1860(.A1(new_n1924_), .A2(new_n1919_), .ZN(new_n1925_));
  NAND3_X1  g1861(.A1(new_n1913_), .A2(new_n1918_), .A3(new_n1920_), .ZN(new_n1926_));
  AOI21_X1  g1862(.A(new_n1731_), .B1(new_n1725_), .B2(new_n1730_), .ZN(new_n1927_));
  OAI211_X1 g1863(.A(new_n1925_), .B(new_n1926_), .C1(new_n1927_), .C2(new_n1757_), .ZN(new_n1928_));
  NOR2_X1   g1864(.A1(new_n76_), .A2(new_n1741_), .ZN(new_n1929_));
  INV_X1    g1865(.A(new_n1929_), .ZN(new_n1930_));
  NAND3_X1  g1866(.A1(new_n1923_), .A2(new_n1928_), .A3(new_n1930_), .ZN(new_n1931_));
  INV_X1    g1867(.A(new_n1931_), .ZN(new_n1932_));
  AOI21_X1  g1868(.A(new_n1930_), .B1(new_n1923_), .B2(new_n1928_), .ZN(new_n1933_));
  OAI211_X1 g1869(.A(new_n1749_), .B(new_n1753_), .C1(new_n1932_), .C2(new_n1933_), .ZN(new_n1934_));
  NAND2_X1  g1870(.A1(new_n1923_), .A2(new_n1928_), .ZN(new_n1935_));
  NAND2_X1  g1871(.A1(new_n1935_), .A2(new_n1929_), .ZN(new_n1936_));
  AOI21_X1  g1872(.A(new_n1742_), .B1(new_n1736_), .B2(new_n1740_), .ZN(new_n1937_));
  OAI211_X1 g1873(.A(new_n1936_), .B(new_n1931_), .C1(new_n1937_), .C2(new_n1752_), .ZN(new_n1938_));
  NAND2_X1  g1874(.A1(new_n1934_), .A2(new_n1938_), .ZN(new_n1939_));
  NAND2_X1  g1875(.A1(new_n1553_), .A2(new_n1746_), .ZN(new_n1940_));
  XNOR2_X1  g1876(.A(new_n1939_), .B(new_n1940_), .ZN(G6160gat));
  AOI21_X1  g1877(.A(new_n1909_), .B1(new_n1903_), .B2(new_n1908_), .ZN(new_n1942_));
  AOI22_X1  g1878(.A1(new_n1768_), .A2(new_n1764_), .B1(new_n1905_), .B2(new_n1906_), .ZN(new_n1943_));
  NOR2_X1   g1879(.A1(new_n1942_), .A2(new_n1943_), .ZN(new_n1944_));
  NOR2_X1   g1880(.A1(new_n146_), .A2(new_n1155_), .ZN(new_n1945_));
  INV_X1    g1881(.A(new_n1945_), .ZN(new_n1946_));
  AOI21_X1  g1882(.A(new_n1869_), .B1(new_n1863_), .B2(new_n1868_), .ZN(new_n1947_));
  AOI22_X1  g1883(.A1(new_n1788_), .A2(new_n1784_), .B1(new_n1865_), .B2(new_n1866_), .ZN(new_n1948_));
  NOR2_X1   g1884(.A1(new_n1947_), .A2(new_n1948_), .ZN(new_n1949_));
  NOR2_X1   g1885(.A1(new_n889_), .A2(new_n544_), .ZN(new_n1950_));
  INV_X1    g1886(.A(new_n1950_), .ZN(new_n1951_));
  NOR2_X1   g1887(.A1(new_n1041_), .A2(new_n190_), .ZN(new_n1952_));
  INV_X1    g1888(.A(new_n1952_), .ZN(new_n1953_));
  NAND2_X1  g1889(.A1(new_n1808_), .A2(new_n1809_), .ZN(new_n1954_));
  NAND2_X1  g1890(.A1(new_n1954_), .A2(new_n1810_), .ZN(new_n1955_));
  OAI21_X1  g1891(.A(new_n1806_), .B1(new_n1613_), .B2(new_n1615_), .ZN(new_n1956_));
  NAND2_X1  g1892(.A1(new_n1956_), .A2(new_n1807_), .ZN(new_n1957_));
  NOR2_X1   g1893(.A1(new_n1805_), .A2(new_n130_), .ZN(new_n1958_));
  INV_X1    g1894(.A(new_n1958_), .ZN(new_n1959_));
  NAND3_X1  g1895(.A1(new_n1955_), .A2(new_n1957_), .A3(new_n1959_), .ZN(new_n1960_));
  AOI22_X1  g1896(.A1(new_n1808_), .A2(new_n1809_), .B1(G239gat), .B2(G324gat), .ZN(new_n1961_));
  INV_X1    g1897(.A(new_n1957_), .ZN(new_n1962_));
  OAI21_X1  g1898(.A(new_n1958_), .B1(new_n1961_), .B2(new_n1962_), .ZN(new_n1963_));
  NAND2_X1  g1899(.A1(G239gat), .A2(G341gat), .ZN(new_n1964_));
  AND3_X1   g1900(.A1(new_n1960_), .A2(new_n1963_), .A3(new_n1964_), .ZN(new_n1965_));
  AOI21_X1  g1901(.A(new_n1964_), .B1(new_n1960_), .B2(new_n1963_), .ZN(new_n1966_));
  NOR2_X1   g1902(.A1(new_n1965_), .A2(new_n1966_), .ZN(new_n1967_));
  INV_X1    g1903(.A(new_n1967_), .ZN(new_n1968_));
  OAI21_X1  g1904(.A(new_n1824_), .B1(new_n1818_), .B2(new_n1820_), .ZN(new_n1969_));
  AOI21_X1  g1905(.A(new_n1813_), .B1(new_n1815_), .B2(new_n1817_), .ZN(new_n1970_));
  INV_X1    g1906(.A(new_n1970_), .ZN(new_n1971_));
  NAND3_X1  g1907(.A1(new_n1968_), .A2(new_n1969_), .A3(new_n1971_), .ZN(new_n1972_));
  AOI21_X1  g1908(.A(new_n1804_), .B1(new_n1822_), .B2(new_n1823_), .ZN(new_n1973_));
  OAI21_X1  g1909(.A(new_n1967_), .B1(new_n1973_), .B2(new_n1970_), .ZN(new_n1974_));
  AOI21_X1  g1910(.A(new_n1953_), .B1(new_n1972_), .B2(new_n1974_), .ZN(new_n1975_));
  INV_X1    g1911(.A(new_n1975_), .ZN(new_n1976_));
  NAND3_X1  g1912(.A1(new_n1972_), .A2(new_n1974_), .A3(new_n1953_), .ZN(new_n1977_));
  NAND2_X1  g1913(.A1(new_n1976_), .A2(new_n1977_), .ZN(new_n1978_));
  NAND2_X1  g1914(.A1(new_n1832_), .A2(new_n1835_), .ZN(new_n1979_));
  OAI21_X1  g1915(.A(new_n1826_), .B1(new_n1827_), .B2(new_n1830_), .ZN(new_n1980_));
  NAND3_X1  g1916(.A1(new_n1978_), .A2(new_n1979_), .A3(new_n1980_), .ZN(new_n1981_));
  AND3_X1   g1917(.A1(new_n1972_), .A2(new_n1974_), .A3(new_n1953_), .ZN(new_n1982_));
  NOR2_X1   g1918(.A1(new_n1982_), .A2(new_n1975_), .ZN(new_n1983_));
  INV_X1    g1919(.A(new_n1980_), .ZN(new_n1984_));
  AOI21_X1  g1920(.A(new_n1833_), .B1(new_n1829_), .B2(new_n1831_), .ZN(new_n1985_));
  OAI21_X1  g1921(.A(new_n1983_), .B1(new_n1984_), .B2(new_n1985_), .ZN(new_n1986_));
  NAND2_X1  g1922(.A1(new_n1981_), .A2(new_n1986_), .ZN(new_n1987_));
  NOR2_X1   g1923(.A1(new_n873_), .A2(new_n253_), .ZN(new_n1988_));
  NAND2_X1  g1924(.A1(new_n1987_), .A2(new_n1988_), .ZN(new_n1989_));
  OAI211_X1 g1925(.A(new_n1981_), .B(new_n1986_), .C1(new_n873_), .C2(new_n253_), .ZN(new_n1990_));
  NAND2_X1  g1926(.A1(new_n1989_), .A2(new_n1990_), .ZN(new_n1991_));
  AOI21_X1  g1927(.A(new_n1799_), .B1(new_n1838_), .B2(new_n1840_), .ZN(new_n1992_));
  INV_X1    g1928(.A(new_n1992_), .ZN(new_n1993_));
  AOI21_X1  g1929(.A(new_n1802_), .B1(new_n1834_), .B2(new_n1836_), .ZN(new_n1994_));
  INV_X1    g1930(.A(new_n1994_), .ZN(new_n1995_));
  NAND3_X1  g1931(.A1(new_n1991_), .A2(new_n1993_), .A3(new_n1995_), .ZN(new_n1996_));
  OAI211_X1 g1932(.A(new_n1989_), .B(new_n1990_), .C1(new_n1992_), .C2(new_n1994_), .ZN(new_n1997_));
  NAND2_X1  g1933(.A1(new_n1996_), .A2(new_n1997_), .ZN(new_n1998_));
  NOR2_X1   g1934(.A1(new_n719_), .A2(new_n336_), .ZN(new_n1999_));
  NAND2_X1  g1935(.A1(new_n1998_), .A2(new_n1999_), .ZN(new_n2000_));
  INV_X1    g1936(.A(new_n1999_), .ZN(new_n2001_));
  NAND3_X1  g1937(.A1(new_n1996_), .A2(new_n1997_), .A3(new_n2001_), .ZN(new_n2002_));
  NAND2_X1  g1938(.A1(new_n2000_), .A2(new_n2002_), .ZN(new_n2003_));
  AOI21_X1  g1939(.A(new_n1849_), .B1(new_n1843_), .B2(new_n1848_), .ZN(new_n2004_));
  AOI22_X1  g1940(.A1(new_n1794_), .A2(new_n1798_), .B1(new_n1845_), .B2(new_n1846_), .ZN(new_n2005_));
  NOR2_X1   g1941(.A1(new_n2004_), .A2(new_n2005_), .ZN(new_n2006_));
  NAND2_X1  g1942(.A1(new_n2003_), .A2(new_n2006_), .ZN(new_n2007_));
  OAI211_X1 g1943(.A(new_n2000_), .B(new_n2002_), .C1(new_n2004_), .C2(new_n2005_), .ZN(new_n2008_));
  NAND2_X1  g1944(.A1(new_n2007_), .A2(new_n2008_), .ZN(new_n2009_));
  NOR2_X1   g1945(.A1(new_n876_), .A2(new_n432_), .ZN(new_n2010_));
  NAND2_X1  g1946(.A1(new_n2009_), .A2(new_n2010_), .ZN(new_n2011_));
  INV_X1    g1947(.A(new_n2010_), .ZN(new_n2012_));
  NAND3_X1  g1948(.A1(new_n2007_), .A2(new_n2008_), .A3(new_n2012_), .ZN(new_n2013_));
  NAND2_X1  g1949(.A1(new_n2011_), .A2(new_n2013_), .ZN(new_n2014_));
  AOI21_X1  g1950(.A(new_n1859_), .B1(new_n1854_), .B2(new_n1858_), .ZN(new_n2015_));
  AOI22_X1  g1951(.A1(new_n1793_), .A2(new_n1789_), .B1(new_n1856_), .B2(new_n1851_), .ZN(new_n2016_));
  NOR2_X1   g1952(.A1(new_n2015_), .A2(new_n2016_), .ZN(new_n2017_));
  NAND2_X1  g1953(.A1(new_n2014_), .A2(new_n2017_), .ZN(new_n2018_));
  OAI211_X1 g1954(.A(new_n2011_), .B(new_n2013_), .C1(new_n2016_), .C2(new_n2015_), .ZN(new_n2019_));
  AOI21_X1  g1955(.A(new_n1951_), .B1(new_n2018_), .B2(new_n2019_), .ZN(new_n2020_));
  NAND3_X1  g1956(.A1(new_n2018_), .A2(new_n2019_), .A3(new_n1951_), .ZN(new_n2021_));
  INV_X1    g1957(.A(new_n2021_), .ZN(new_n2022_));
  OAI21_X1  g1958(.A(new_n1949_), .B1(new_n2020_), .B2(new_n2022_), .ZN(new_n2023_));
  NAND2_X1  g1959(.A1(new_n2018_), .A2(new_n2019_), .ZN(new_n2024_));
  NAND2_X1  g1960(.A1(new_n2024_), .A2(new_n1950_), .ZN(new_n2025_));
  OAI211_X1 g1961(.A(new_n2025_), .B(new_n2021_), .C1(new_n1948_), .C2(new_n1947_), .ZN(new_n2026_));
  NAND2_X1  g1962(.A1(new_n2023_), .A2(new_n2026_), .ZN(new_n2027_));
  NOR2_X1   g1963(.A1(new_n733_), .A2(new_n673_), .ZN(new_n2028_));
  NAND2_X1  g1964(.A1(new_n2027_), .A2(new_n2028_), .ZN(new_n2029_));
  INV_X1    g1965(.A(new_n2028_), .ZN(new_n2030_));
  NAND3_X1  g1966(.A1(new_n2023_), .A2(new_n2026_), .A3(new_n2030_), .ZN(new_n2031_));
  NOR2_X1   g1967(.A1(new_n1871_), .A2(new_n1872_), .ZN(new_n2032_));
  NOR2_X1   g1968(.A1(new_n1877_), .A2(new_n1782_), .ZN(new_n2033_));
  NOR2_X1   g1969(.A1(new_n2032_), .A2(new_n2033_), .ZN(new_n2034_));
  AOI21_X1  g1970(.A(new_n1879_), .B1(new_n1873_), .B2(new_n1878_), .ZN(new_n2035_));
  OAI211_X1 g1971(.A(new_n2029_), .B(new_n2031_), .C1(new_n2034_), .C2(new_n2035_), .ZN(new_n2036_));
  NAND2_X1  g1972(.A1(new_n1884_), .A2(new_n1880_), .ZN(new_n2037_));
  INV_X1    g1973(.A(new_n2034_), .ZN(new_n2038_));
  AND3_X1   g1974(.A1(new_n2023_), .A2(new_n2026_), .A3(new_n2030_), .ZN(new_n2039_));
  AOI21_X1  g1975(.A(new_n2030_), .B1(new_n2023_), .B2(new_n2026_), .ZN(new_n2040_));
  OAI211_X1 g1976(.A(new_n2037_), .B(new_n2038_), .C1(new_n2039_), .C2(new_n2040_), .ZN(new_n2041_));
  NAND2_X1  g1977(.A1(new_n2036_), .A2(new_n2041_), .ZN(new_n2042_));
  NOR2_X1   g1978(.A1(new_n276_), .A2(new_n816_), .ZN(new_n2043_));
  NAND2_X1  g1979(.A1(new_n2042_), .A2(new_n2043_), .ZN(new_n2044_));
  INV_X1    g1980(.A(new_n2043_), .ZN(new_n2045_));
  NAND3_X1  g1981(.A1(new_n2036_), .A2(new_n2041_), .A3(new_n2045_), .ZN(new_n2046_));
  NOR2_X1   g1982(.A1(new_n1881_), .A2(new_n1882_), .ZN(new_n2047_));
  NOR2_X1   g1983(.A1(new_n1887_), .A2(new_n1777_), .ZN(new_n2048_));
  NOR2_X1   g1984(.A1(new_n2047_), .A2(new_n2048_), .ZN(new_n2049_));
  AOI21_X1  g1985(.A(new_n1889_), .B1(new_n1883_), .B2(new_n1888_), .ZN(new_n2050_));
  OAI211_X1 g1986(.A(new_n2044_), .B(new_n2046_), .C1(new_n2049_), .C2(new_n2050_), .ZN(new_n2051_));
  NAND2_X1  g1987(.A1(new_n1894_), .A2(new_n1890_), .ZN(new_n2052_));
  INV_X1    g1988(.A(new_n2049_), .ZN(new_n2053_));
  AND3_X1   g1989(.A1(new_n2036_), .A2(new_n2041_), .A3(new_n2045_), .ZN(new_n2054_));
  AOI21_X1  g1990(.A(new_n2045_), .B1(new_n2036_), .B2(new_n2041_), .ZN(new_n2055_));
  OAI211_X1 g1991(.A(new_n2052_), .B(new_n2053_), .C1(new_n2054_), .C2(new_n2055_), .ZN(new_n2056_));
  NAND2_X1  g1992(.A1(new_n2051_), .A2(new_n2056_), .ZN(new_n2057_));
  NOR2_X1   g1993(.A1(new_n205_), .A2(new_n980_), .ZN(new_n2058_));
  NAND2_X1  g1994(.A1(new_n2057_), .A2(new_n2058_), .ZN(new_n2059_));
  OAI211_X1 g1995(.A(new_n2051_), .B(new_n2056_), .C1(new_n205_), .C2(new_n980_), .ZN(new_n2060_));
  NAND2_X1  g1996(.A1(new_n2059_), .A2(new_n2060_), .ZN(new_n2061_));
  AOI21_X1  g1997(.A(new_n1899_), .B1(new_n1893_), .B2(new_n1898_), .ZN(new_n2062_));
  NOR2_X1   g1998(.A1(new_n1891_), .A2(new_n1892_), .ZN(new_n2063_));
  NOR2_X1   g1999(.A1(new_n1897_), .A2(new_n1772_), .ZN(new_n2064_));
  NOR2_X1   g2000(.A1(new_n2063_), .A2(new_n2064_), .ZN(new_n2065_));
  NOR2_X1   g2001(.A1(new_n2062_), .A2(new_n2065_), .ZN(new_n2066_));
  NAND2_X1  g2002(.A1(new_n2061_), .A2(new_n2066_), .ZN(new_n2067_));
  OAI211_X1 g2003(.A(new_n2059_), .B(new_n2060_), .C1(new_n2065_), .C2(new_n2062_), .ZN(new_n2068_));
  AOI21_X1  g2004(.A(new_n1946_), .B1(new_n2067_), .B2(new_n2068_), .ZN(new_n2069_));
  NAND3_X1  g2005(.A1(new_n2067_), .A2(new_n2068_), .A3(new_n1946_), .ZN(new_n2070_));
  INV_X1    g2006(.A(new_n2070_), .ZN(new_n2071_));
  OAI21_X1  g2007(.A(new_n1944_), .B1(new_n2069_), .B2(new_n2071_), .ZN(new_n2072_));
  NAND2_X1  g2008(.A1(new_n2067_), .A2(new_n2068_), .ZN(new_n2073_));
  NAND2_X1  g2009(.A1(new_n2073_), .A2(new_n1945_), .ZN(new_n2074_));
  OAI211_X1 g2010(.A(new_n2074_), .B(new_n2070_), .C1(new_n1943_), .C2(new_n1942_), .ZN(new_n2075_));
  NAND2_X1  g2011(.A1(new_n2072_), .A2(new_n2075_), .ZN(new_n2076_));
  NOR2_X1   g2012(.A1(new_n113_), .A2(new_n1345_), .ZN(new_n2077_));
  NAND2_X1  g2013(.A1(new_n2076_), .A2(new_n2077_), .ZN(new_n2078_));
  INV_X1    g2014(.A(new_n2077_), .ZN(new_n2079_));
  NAND3_X1  g2015(.A1(new_n2072_), .A2(new_n2075_), .A3(new_n2079_), .ZN(new_n2080_));
  NOR2_X1   g2016(.A1(new_n1911_), .A2(new_n1912_), .ZN(new_n2081_));
  NOR2_X1   g2017(.A1(new_n1917_), .A2(new_n1762_), .ZN(new_n2082_));
  NOR2_X1   g2018(.A1(new_n2081_), .A2(new_n2082_), .ZN(new_n2083_));
  AOI21_X1  g2019(.A(new_n1919_), .B1(new_n1913_), .B2(new_n1918_), .ZN(new_n2084_));
  OAI211_X1 g2020(.A(new_n2078_), .B(new_n2080_), .C1(new_n2083_), .C2(new_n2084_), .ZN(new_n2085_));
  INV_X1    g2021(.A(new_n2084_), .ZN(new_n2086_));
  INV_X1    g2022(.A(new_n2083_), .ZN(new_n2087_));
  AND3_X1   g2023(.A1(new_n2072_), .A2(new_n2075_), .A3(new_n2079_), .ZN(new_n2088_));
  AOI21_X1  g2024(.A(new_n2079_), .B1(new_n2072_), .B2(new_n2075_), .ZN(new_n2089_));
  OAI211_X1 g2025(.A(new_n2086_), .B(new_n2087_), .C1(new_n2088_), .C2(new_n2089_), .ZN(new_n2090_));
  NAND2_X1  g2026(.A1(new_n2085_), .A2(new_n2090_), .ZN(new_n2091_));
  NOR2_X1   g2027(.A1(new_n86_), .A2(new_n1741_), .ZN(new_n2092_));
  NAND2_X1  g2028(.A1(new_n2091_), .A2(new_n2092_), .ZN(new_n2093_));
  INV_X1    g2029(.A(new_n2092_), .ZN(new_n2094_));
  NAND3_X1  g2030(.A1(new_n2085_), .A2(new_n2090_), .A3(new_n2094_), .ZN(new_n2095_));
  NOR2_X1   g2031(.A1(new_n1921_), .A2(new_n1922_), .ZN(new_n2096_));
  NOR2_X1   g2032(.A1(new_n1927_), .A2(new_n1757_), .ZN(new_n2097_));
  NOR2_X1   g2033(.A1(new_n2096_), .A2(new_n2097_), .ZN(new_n2098_));
  AOI21_X1  g2034(.A(new_n1929_), .B1(new_n1923_), .B2(new_n1928_), .ZN(new_n2099_));
  OAI211_X1 g2035(.A(new_n2093_), .B(new_n2095_), .C1(new_n2098_), .C2(new_n2099_), .ZN(new_n2100_));
  INV_X1    g2036(.A(new_n2098_), .ZN(new_n2101_));
  NAND2_X1  g2037(.A1(new_n1935_), .A2(new_n1930_), .ZN(new_n2102_));
  AND3_X1   g2038(.A1(new_n2085_), .A2(new_n2090_), .A3(new_n2094_), .ZN(new_n2103_));
  AOI21_X1  g2039(.A(new_n2094_), .B1(new_n2085_), .B2(new_n2090_), .ZN(new_n2104_));
  OAI211_X1 g2040(.A(new_n2101_), .B(new_n2102_), .C1(new_n2103_), .C2(new_n2104_), .ZN(new_n2105_));
  NAND2_X1  g2041(.A1(new_n2100_), .A2(new_n2105_), .ZN(new_n2106_));
  NAND2_X1  g2042(.A1(new_n1939_), .A2(new_n1940_), .ZN(new_n2107_));
  NOR2_X1   g2043(.A1(new_n1932_), .A2(new_n1933_), .ZN(new_n2108_));
  NOR2_X1   g2044(.A1(new_n1937_), .A2(new_n1752_), .ZN(new_n2109_));
  NOR2_X1   g2045(.A1(new_n2108_), .A2(new_n2109_), .ZN(new_n2110_));
  INV_X1    g2046(.A(new_n2110_), .ZN(new_n2111_));
  AOI21_X1  g2047(.A(new_n2106_), .B1(new_n2107_), .B2(new_n2111_), .ZN(new_n2112_));
  AOI22_X1  g2048(.A1(new_n1934_), .A2(new_n1938_), .B1(new_n1746_), .B2(new_n1553_), .ZN(new_n2113_));
  OAI21_X1  g2049(.A(new_n2106_), .B1(new_n2113_), .B2(new_n2110_), .ZN(new_n2114_));
  AOI21_X1  g2050(.A(new_n2112_), .B1(new_n2106_), .B2(new_n2114_), .ZN(G6170gat));
  AOI21_X1  g2051(.A(new_n2077_), .B1(new_n2072_), .B2(new_n2075_), .ZN(new_n2116_));
  AOI21_X1  g2052(.A(new_n1944_), .B1(new_n2074_), .B2(new_n2070_), .ZN(new_n2117_));
  NOR2_X1   g2053(.A1(new_n2116_), .A2(new_n2117_), .ZN(new_n2118_));
  INV_X1    g2054(.A(new_n2118_), .ZN(new_n2119_));
  NOR2_X1   g2055(.A1(new_n876_), .A2(new_n544_), .ZN(new_n2120_));
  AOI21_X1  g2056(.A(new_n1988_), .B1(new_n1981_), .B2(new_n1986_), .ZN(new_n2121_));
  AOI21_X1  g2057(.A(new_n1983_), .B1(new_n1980_), .B2(new_n1979_), .ZN(new_n2122_));
  OR2_X1    g2058(.A1(new_n2121_), .A2(new_n2122_), .ZN(new_n2123_));
  INV_X1    g2059(.A(new_n1974_), .ZN(new_n2124_));
  NOR3_X1   g2060(.A1(new_n1973_), .A2(new_n1967_), .A3(new_n1970_), .ZN(new_n2125_));
  OAI21_X1  g2061(.A(new_n1953_), .B1(new_n2124_), .B2(new_n2125_), .ZN(new_n2126_));
  OAI21_X1  g2062(.A(new_n1968_), .B1(new_n1973_), .B2(new_n1970_), .ZN(new_n2127_));
  NAND2_X1  g2063(.A1(new_n2126_), .A2(new_n2127_), .ZN(new_n2128_));
  NAND2_X1  g2064(.A1(new_n1960_), .A2(new_n1963_), .ZN(new_n2129_));
  NAND2_X1  g2065(.A1(new_n2129_), .A2(new_n1964_), .ZN(new_n2130_));
  AOI21_X1  g2066(.A(new_n1958_), .B1(new_n1955_), .B2(new_n1957_), .ZN(new_n2131_));
  INV_X1    g2067(.A(new_n2131_), .ZN(new_n2132_));
  NAND2_X1  g2068(.A1(new_n2130_), .A2(new_n2132_), .ZN(new_n2133_));
  NOR2_X1   g2069(.A1(new_n1805_), .A2(new_n178_), .ZN(new_n2134_));
  NAND2_X1  g2070(.A1(new_n2133_), .A2(new_n2134_), .ZN(new_n2135_));
  INV_X1    g2071(.A(new_n2134_), .ZN(new_n2136_));
  NAND3_X1  g2072(.A1(new_n2130_), .A2(new_n2132_), .A3(new_n2136_), .ZN(new_n2137_));
  NAND2_X1  g2073(.A1(new_n2135_), .A2(new_n2137_), .ZN(new_n2138_));
  NOR2_X1   g2074(.A1(new_n1220_), .A2(new_n190_), .ZN(new_n2139_));
  NOR2_X1   g2075(.A1(new_n2138_), .A2(new_n2139_), .ZN(new_n2140_));
  INV_X1    g2076(.A(new_n2139_), .ZN(new_n2141_));
  AOI21_X1  g2077(.A(new_n2141_), .B1(new_n2135_), .B2(new_n2137_), .ZN(new_n2142_));
  NOR2_X1   g2078(.A1(new_n2140_), .A2(new_n2142_), .ZN(new_n2143_));
  NAND2_X1  g2079(.A1(new_n2128_), .A2(new_n2143_), .ZN(new_n2144_));
  OR2_X1    g2080(.A1(new_n2140_), .A2(new_n2142_), .ZN(new_n2145_));
  NAND3_X1  g2081(.A1(new_n2145_), .A2(new_n2127_), .A3(new_n2126_), .ZN(new_n2146_));
  NAND2_X1  g2082(.A1(new_n2144_), .A2(new_n2146_), .ZN(new_n2147_));
  NOR2_X1   g2083(.A1(new_n1041_), .A2(new_n253_), .ZN(new_n2148_));
  INV_X1    g2084(.A(new_n2148_), .ZN(new_n2149_));
  XNOR2_X1  g2085(.A(new_n2147_), .B(new_n2149_), .ZN(new_n2150_));
  NAND2_X1  g2086(.A1(new_n2123_), .A2(new_n2150_), .ZN(new_n2151_));
  XNOR2_X1  g2087(.A(new_n2147_), .B(new_n2148_), .ZN(new_n2152_));
  NOR2_X1   g2088(.A1(new_n2121_), .A2(new_n2122_), .ZN(new_n2153_));
  NAND2_X1  g2089(.A1(new_n2152_), .A2(new_n2153_), .ZN(new_n2154_));
  NAND2_X1  g2090(.A1(new_n2151_), .A2(new_n2154_), .ZN(new_n2155_));
  NAND3_X1  g2091(.A1(new_n2155_), .A2(G205gat), .A3(G392gat), .ZN(new_n2156_));
  NAND2_X1  g2092(.A1(G205gat), .A2(G392gat), .ZN(new_n2157_));
  NAND3_X1  g2093(.A1(new_n2151_), .A2(new_n2154_), .A3(new_n2157_), .ZN(new_n2158_));
  NAND2_X1  g2094(.A1(new_n2156_), .A2(new_n2158_), .ZN(new_n2159_));
  NAND2_X1  g2095(.A1(new_n1993_), .A2(new_n1995_), .ZN(new_n2160_));
  NAND2_X1  g2096(.A1(new_n2160_), .A2(new_n1991_), .ZN(new_n2161_));
  NAND2_X1  g2097(.A1(new_n1998_), .A2(new_n2001_), .ZN(new_n2162_));
  NAND3_X1  g2098(.A1(new_n2159_), .A2(new_n2161_), .A3(new_n2162_), .ZN(new_n2163_));
  INV_X1    g2099(.A(new_n2162_), .ZN(new_n2164_));
  INV_X1    g2100(.A(new_n2161_), .ZN(new_n2165_));
  OAI211_X1 g2101(.A(new_n2156_), .B(new_n2158_), .C1(new_n2164_), .C2(new_n2165_), .ZN(new_n2166_));
  NAND2_X1  g2102(.A1(new_n2163_), .A2(new_n2166_), .ZN(new_n2167_));
  NOR2_X1   g2103(.A1(new_n719_), .A2(new_n432_), .ZN(new_n2168_));
  NAND2_X1  g2104(.A1(new_n2167_), .A2(new_n2168_), .ZN(new_n2169_));
  OAI211_X1 g2105(.A(new_n2163_), .B(new_n2166_), .C1(new_n719_), .C2(new_n432_), .ZN(new_n2170_));
  NAND2_X1  g2106(.A1(new_n2169_), .A2(new_n2170_), .ZN(new_n2171_));
  AOI21_X1  g2107(.A(new_n2006_), .B1(new_n2000_), .B2(new_n2002_), .ZN(new_n2172_));
  AOI21_X1  g2108(.A(new_n2172_), .B1(new_n2009_), .B2(new_n2012_), .ZN(new_n2173_));
  AND2_X1   g2109(.A1(new_n2171_), .A2(new_n2173_), .ZN(new_n2174_));
  NOR2_X1   g2110(.A1(new_n2171_), .A2(new_n2173_), .ZN(new_n2175_));
  OAI21_X1  g2111(.A(new_n2120_), .B1(new_n2174_), .B2(new_n2175_), .ZN(new_n2176_));
  NAND2_X1  g2112(.A1(new_n2171_), .A2(new_n2173_), .ZN(new_n2177_));
  INV_X1    g2113(.A(new_n2120_), .ZN(new_n2178_));
  AOI21_X1  g2114(.A(new_n2173_), .B1(new_n2169_), .B2(new_n2170_), .ZN(new_n2179_));
  OAI211_X1 g2115(.A(new_n2177_), .B(new_n2178_), .C1(new_n2179_), .C2(new_n2173_), .ZN(new_n2180_));
  NAND2_X1  g2116(.A1(new_n2176_), .A2(new_n2180_), .ZN(new_n2181_));
  AOI21_X1  g2117(.A(new_n1950_), .B1(new_n2018_), .B2(new_n2019_), .ZN(new_n2182_));
  AOI21_X1  g2118(.A(new_n2017_), .B1(new_n2011_), .B2(new_n2013_), .ZN(new_n2183_));
  NOR2_X1   g2119(.A1(new_n2182_), .A2(new_n2183_), .ZN(new_n2184_));
  NAND2_X1  g2120(.A1(new_n2181_), .A2(new_n2184_), .ZN(new_n2185_));
  OAI211_X1 g2121(.A(new_n2176_), .B(new_n2180_), .C1(new_n2182_), .C2(new_n2183_), .ZN(new_n2186_));
  NAND2_X1  g2122(.A1(new_n2185_), .A2(new_n2186_), .ZN(new_n2187_));
  NOR2_X1   g2123(.A1(new_n889_), .A2(new_n673_), .ZN(new_n2188_));
  NAND2_X1  g2124(.A1(new_n2187_), .A2(new_n2188_), .ZN(new_n2189_));
  INV_X1    g2125(.A(new_n2188_), .ZN(new_n2190_));
  NAND3_X1  g2126(.A1(new_n2185_), .A2(new_n2186_), .A3(new_n2190_), .ZN(new_n2191_));
  AOI21_X1  g2127(.A(new_n1949_), .B1(new_n2025_), .B2(new_n2021_), .ZN(new_n2192_));
  AOI21_X1  g2128(.A(new_n2028_), .B1(new_n2023_), .B2(new_n2026_), .ZN(new_n2193_));
  OAI211_X1 g2129(.A(new_n2189_), .B(new_n2191_), .C1(new_n2192_), .C2(new_n2193_), .ZN(new_n2194_));
  NOR2_X1   g2130(.A1(new_n2193_), .A2(new_n2192_), .ZN(new_n2195_));
  INV_X1    g2131(.A(new_n2191_), .ZN(new_n2196_));
  AOI21_X1  g2132(.A(new_n2190_), .B1(new_n2185_), .B2(new_n2186_), .ZN(new_n2197_));
  OAI21_X1  g2133(.A(new_n2195_), .B1(new_n2196_), .B2(new_n2197_), .ZN(new_n2198_));
  NAND2_X1  g2134(.A1(new_n2194_), .A2(new_n2198_), .ZN(new_n2199_));
  NOR2_X1   g2135(.A1(new_n733_), .A2(new_n816_), .ZN(new_n2200_));
  NAND2_X1  g2136(.A1(new_n2199_), .A2(new_n2200_), .ZN(new_n2201_));
  OAI211_X1 g2137(.A(new_n2194_), .B(new_n2198_), .C1(new_n733_), .C2(new_n816_), .ZN(new_n2202_));
  NAND2_X1  g2138(.A1(new_n2201_), .A2(new_n2202_), .ZN(new_n2203_));
  AOI21_X1  g2139(.A(new_n2043_), .B1(new_n2036_), .B2(new_n2041_), .ZN(new_n2204_));
  AOI22_X1  g2140(.A1(new_n2029_), .A2(new_n2031_), .B1(new_n2037_), .B2(new_n2038_), .ZN(new_n2205_));
  NOR2_X1   g2141(.A1(new_n2204_), .A2(new_n2205_), .ZN(new_n2206_));
  NAND2_X1  g2142(.A1(new_n2203_), .A2(new_n2206_), .ZN(new_n2207_));
  OAI211_X1 g2143(.A(new_n2201_), .B(new_n2202_), .C1(new_n2205_), .C2(new_n2204_), .ZN(new_n2208_));
  NAND2_X1  g2144(.A1(new_n2207_), .A2(new_n2208_), .ZN(new_n2209_));
  NOR2_X1   g2145(.A1(new_n276_), .A2(new_n980_), .ZN(new_n2210_));
  NAND2_X1  g2146(.A1(new_n2209_), .A2(new_n2210_), .ZN(new_n2211_));
  INV_X1    g2147(.A(new_n2210_), .ZN(new_n2212_));
  NAND3_X1  g2148(.A1(new_n2207_), .A2(new_n2208_), .A3(new_n2212_), .ZN(new_n2213_));
  AOI22_X1  g2149(.A1(new_n2044_), .A2(new_n2046_), .B1(new_n2052_), .B2(new_n2053_), .ZN(new_n2214_));
  AOI21_X1  g2150(.A(new_n2058_), .B1(new_n2051_), .B2(new_n2056_), .ZN(new_n2215_));
  OAI211_X1 g2151(.A(new_n2211_), .B(new_n2213_), .C1(new_n2214_), .C2(new_n2215_), .ZN(new_n2216_));
  NOR2_X1   g2152(.A1(new_n2215_), .A2(new_n2214_), .ZN(new_n2217_));
  INV_X1    g2153(.A(new_n2213_), .ZN(new_n2218_));
  AOI21_X1  g2154(.A(new_n2212_), .B1(new_n2207_), .B2(new_n2208_), .ZN(new_n2219_));
  OAI21_X1  g2155(.A(new_n2217_), .B1(new_n2218_), .B2(new_n2219_), .ZN(new_n2220_));
  NAND2_X1  g2156(.A1(new_n2216_), .A2(new_n2220_), .ZN(new_n2221_));
  NOR2_X1   g2157(.A1(new_n205_), .A2(new_n1155_), .ZN(new_n2222_));
  NAND2_X1  g2158(.A1(new_n2221_), .A2(new_n2222_), .ZN(new_n2223_));
  INV_X1    g2159(.A(new_n2222_), .ZN(new_n2224_));
  NAND3_X1  g2160(.A1(new_n2216_), .A2(new_n2220_), .A3(new_n2224_), .ZN(new_n2225_));
  AOI21_X1  g2161(.A(new_n2066_), .B1(new_n2059_), .B2(new_n2060_), .ZN(new_n2226_));
  AOI21_X1  g2162(.A(new_n1945_), .B1(new_n2067_), .B2(new_n2068_), .ZN(new_n2227_));
  OAI211_X1 g2163(.A(new_n2223_), .B(new_n2225_), .C1(new_n2226_), .C2(new_n2227_), .ZN(new_n2228_));
  NOR2_X1   g2164(.A1(new_n2227_), .A2(new_n2226_), .ZN(new_n2229_));
  INV_X1    g2165(.A(new_n2225_), .ZN(new_n2230_));
  AOI21_X1  g2166(.A(new_n2224_), .B1(new_n2216_), .B2(new_n2220_), .ZN(new_n2231_));
  OAI21_X1  g2167(.A(new_n2229_), .B1(new_n2230_), .B2(new_n2231_), .ZN(new_n2232_));
  NAND2_X1  g2168(.A1(new_n2228_), .A2(new_n2232_), .ZN(new_n2233_));
  NOR2_X1   g2169(.A1(new_n146_), .A2(new_n1345_), .ZN(new_n2234_));
  NAND2_X1  g2170(.A1(new_n2233_), .A2(new_n2234_), .ZN(new_n2235_));
  INV_X1    g2171(.A(new_n2234_), .ZN(new_n2236_));
  NAND3_X1  g2172(.A1(new_n2228_), .A2(new_n2232_), .A3(new_n2236_), .ZN(new_n2237_));
  NAND3_X1  g2173(.A1(new_n2119_), .A2(new_n2235_), .A3(new_n2237_), .ZN(new_n2238_));
  NAND2_X1  g2174(.A1(new_n2235_), .A2(new_n2237_), .ZN(new_n2239_));
  NAND2_X1  g2175(.A1(new_n2239_), .A2(new_n2118_), .ZN(new_n2240_));
  NAND2_X1  g2176(.A1(new_n2238_), .A2(new_n2240_), .ZN(new_n2241_));
  NOR2_X1   g2177(.A1(new_n113_), .A2(new_n1741_), .ZN(new_n2242_));
  NAND2_X1  g2178(.A1(new_n2241_), .A2(new_n2242_), .ZN(new_n2243_));
  INV_X1    g2179(.A(new_n2242_), .ZN(new_n2244_));
  NAND3_X1  g2180(.A1(new_n2238_), .A2(new_n2240_), .A3(new_n2244_), .ZN(new_n2245_));
  AOI22_X1  g2181(.A1(new_n2078_), .A2(new_n2080_), .B1(new_n2086_), .B2(new_n2087_), .ZN(new_n2246_));
  AOI21_X1  g2182(.A(new_n2092_), .B1(new_n2085_), .B2(new_n2090_), .ZN(new_n2247_));
  OAI211_X1 g2183(.A(new_n2243_), .B(new_n2245_), .C1(new_n2246_), .C2(new_n2247_), .ZN(new_n2248_));
  NOR2_X1   g2184(.A1(new_n2247_), .A2(new_n2246_), .ZN(new_n2249_));
  INV_X1    g2185(.A(new_n2245_), .ZN(new_n2250_));
  AOI21_X1  g2186(.A(new_n2244_), .B1(new_n2238_), .B2(new_n2240_), .ZN(new_n2251_));
  OAI21_X1  g2187(.A(new_n2249_), .B1(new_n2250_), .B2(new_n2251_), .ZN(new_n2252_));
  AND2_X1   g2188(.A1(new_n2248_), .A2(new_n2252_), .ZN(new_n2253_));
  INV_X1    g2189(.A(new_n2253_), .ZN(new_n2254_));
  NAND2_X1  g2190(.A1(new_n2093_), .A2(new_n2095_), .ZN(new_n2255_));
  NAND2_X1  g2191(.A1(new_n2102_), .A2(new_n2101_), .ZN(new_n2256_));
  NAND2_X1  g2192(.A1(new_n2255_), .A2(new_n2256_), .ZN(new_n2257_));
  AOI21_X1  g2193(.A(new_n2254_), .B1(new_n2114_), .B2(new_n2257_), .ZN(new_n2258_));
  AND2_X1   g2194(.A1(new_n2100_), .A2(new_n2105_), .ZN(new_n2259_));
  AOI21_X1  g2195(.A(new_n2259_), .B1(new_n2107_), .B2(new_n2111_), .ZN(new_n2260_));
  INV_X1    g2196(.A(new_n2257_), .ZN(new_n2261_));
  OAI21_X1  g2197(.A(new_n2254_), .B1(new_n2260_), .B2(new_n2261_), .ZN(new_n2262_));
  AOI21_X1  g2198(.A(new_n2258_), .B1(new_n2254_), .B2(new_n2262_), .ZN(G6180gat));
  AND2_X1   g2199(.A1(new_n2155_), .A2(new_n2157_), .ZN(new_n2264_));
  NOR2_X1   g2200(.A1(new_n2150_), .A2(new_n2153_), .ZN(new_n2265_));
  NOR2_X1   g2201(.A1(new_n2264_), .A2(new_n2265_), .ZN(new_n2266_));
  NOR2_X1   g2202(.A1(new_n1041_), .A2(new_n336_), .ZN(new_n2267_));
  INV_X1    g2203(.A(new_n2267_), .ZN(new_n2268_));
  NAND2_X1  g2204(.A1(new_n2147_), .A2(new_n2149_), .ZN(new_n2269_));
  INV_X1    g2205(.A(new_n2128_), .ZN(new_n2270_));
  OAI21_X1  g2206(.A(new_n2269_), .B1(new_n2143_), .B2(new_n2270_), .ZN(new_n2271_));
  NAND2_X1  g2207(.A1(new_n2138_), .A2(new_n2141_), .ZN(new_n2272_));
  NAND2_X1  g2208(.A1(new_n2133_), .A2(new_n2136_), .ZN(new_n2273_));
  NAND2_X1  g2209(.A1(new_n2272_), .A2(new_n2273_), .ZN(new_n2274_));
  NOR2_X1   g2210(.A1(new_n1805_), .A2(new_n190_), .ZN(new_n2275_));
  INV_X1    g2211(.A(new_n2275_), .ZN(new_n2276_));
  NAND2_X1  g2212(.A1(new_n2274_), .A2(new_n2276_), .ZN(new_n2277_));
  NAND2_X1  g2213(.A1(new_n2277_), .A2(new_n2276_), .ZN(new_n2278_));
  NAND2_X1  g2214(.A1(new_n2274_), .A2(new_n2275_), .ZN(new_n2279_));
  NAND2_X1  g2215(.A1(new_n2278_), .A2(new_n2279_), .ZN(new_n2280_));
  NAND2_X1  g2216(.A1(G239gat), .A2(G375gat), .ZN(new_n2281_));
  XNOR2_X1  g2217(.A(new_n2280_), .B(new_n2281_), .ZN(new_n2282_));
  NOR2_X1   g2218(.A1(new_n2271_), .A2(new_n2282_), .ZN(new_n2283_));
  INV_X1    g2219(.A(new_n2283_), .ZN(new_n2284_));
  NAND2_X1  g2220(.A1(new_n2271_), .A2(new_n2282_), .ZN(new_n2285_));
  AOI21_X1  g2221(.A(new_n2268_), .B1(new_n2284_), .B2(new_n2285_), .ZN(new_n2286_));
  INV_X1    g2222(.A(new_n2285_), .ZN(new_n2287_));
  NOR3_X1   g2223(.A1(new_n2287_), .A2(new_n2283_), .A3(new_n2267_), .ZN(new_n2288_));
  OAI21_X1  g2224(.A(new_n2266_), .B1(new_n2286_), .B2(new_n2288_), .ZN(new_n2289_));
  NOR2_X1   g2225(.A1(new_n2286_), .A2(new_n2288_), .ZN(new_n2290_));
  OAI21_X1  g2226(.A(new_n2290_), .B1(new_n2265_), .B2(new_n2264_), .ZN(new_n2291_));
  NOR2_X1   g2227(.A1(new_n873_), .A2(new_n432_), .ZN(new_n2292_));
  INV_X1    g2228(.A(new_n2292_), .ZN(new_n2293_));
  AND3_X1   g2229(.A1(new_n2289_), .A2(new_n2291_), .A3(new_n2293_), .ZN(new_n2294_));
  AOI21_X1  g2230(.A(new_n2293_), .B1(new_n2289_), .B2(new_n2291_), .ZN(new_n2295_));
  NOR2_X1   g2231(.A1(new_n2294_), .A2(new_n2295_), .ZN(new_n2296_));
  OAI21_X1  g2232(.A(new_n2159_), .B1(new_n2164_), .B2(new_n2165_), .ZN(new_n2297_));
  AND2_X1   g2233(.A1(new_n2163_), .A2(new_n2166_), .ZN(new_n2298_));
  OAI21_X1  g2234(.A(new_n2297_), .B1(new_n2298_), .B2(new_n2168_), .ZN(new_n2299_));
  OR2_X1    g2235(.A1(new_n2296_), .A2(new_n2299_), .ZN(new_n2300_));
  NAND2_X1  g2236(.A1(new_n2296_), .A2(new_n2299_), .ZN(new_n2301_));
  NAND2_X1  g2237(.A1(new_n2300_), .A2(new_n2301_), .ZN(new_n2302_));
  NOR2_X1   g2238(.A1(new_n719_), .A2(new_n544_), .ZN(new_n2303_));
  NAND2_X1  g2239(.A1(new_n2302_), .A2(new_n2303_), .ZN(new_n2304_));
  INV_X1    g2240(.A(new_n2303_), .ZN(new_n2305_));
  NAND3_X1  g2241(.A1(new_n2300_), .A2(new_n2301_), .A3(new_n2305_), .ZN(new_n2306_));
  NAND2_X1  g2242(.A1(new_n2304_), .A2(new_n2306_), .ZN(new_n2307_));
  NOR2_X1   g2243(.A1(new_n2174_), .A2(new_n2175_), .ZN(new_n2308_));
  NOR2_X1   g2244(.A1(new_n2308_), .A2(new_n2120_), .ZN(new_n2309_));
  NOR2_X1   g2245(.A1(new_n2309_), .A2(new_n2179_), .ZN(new_n2310_));
  NAND2_X1  g2246(.A1(new_n2307_), .A2(new_n2310_), .ZN(new_n2311_));
  OAI211_X1 g2247(.A(new_n2304_), .B(new_n2306_), .C1(new_n2309_), .C2(new_n2179_), .ZN(new_n2312_));
  NAND2_X1  g2248(.A1(new_n2311_), .A2(new_n2312_), .ZN(new_n2313_));
  NOR2_X1   g2249(.A1(new_n876_), .A2(new_n673_), .ZN(new_n2314_));
  NAND2_X1  g2250(.A1(new_n2313_), .A2(new_n2314_), .ZN(new_n2315_));
  OAI211_X1 g2251(.A(new_n2311_), .B(new_n2312_), .C1(new_n876_), .C2(new_n673_), .ZN(new_n2316_));
  NAND2_X1  g2252(.A1(new_n2315_), .A2(new_n2316_), .ZN(new_n2317_));
  INV_X1    g2253(.A(new_n2184_), .ZN(new_n2318_));
  NAND2_X1  g2254(.A1(new_n2181_), .A2(new_n2318_), .ZN(new_n2319_));
  INV_X1    g2255(.A(new_n2319_), .ZN(new_n2320_));
  AOI21_X1  g2256(.A(new_n2320_), .B1(new_n2187_), .B2(new_n2190_), .ZN(new_n2321_));
  NAND2_X1  g2257(.A1(new_n2317_), .A2(new_n2321_), .ZN(new_n2322_));
  INV_X1    g2258(.A(new_n2321_), .ZN(new_n2323_));
  NAND3_X1  g2259(.A1(new_n2315_), .A2(new_n2323_), .A3(new_n2316_), .ZN(new_n2324_));
  NAND2_X1  g2260(.A1(new_n2322_), .A2(new_n2324_), .ZN(new_n2325_));
  NOR2_X1   g2261(.A1(new_n889_), .A2(new_n816_), .ZN(new_n2326_));
  NAND2_X1  g2262(.A1(new_n2325_), .A2(new_n2326_), .ZN(new_n2327_));
  INV_X1    g2263(.A(new_n2326_), .ZN(new_n2328_));
  NAND3_X1  g2264(.A1(new_n2322_), .A2(new_n2324_), .A3(new_n2328_), .ZN(new_n2329_));
  AOI21_X1  g2265(.A(new_n2195_), .B1(new_n2189_), .B2(new_n2191_), .ZN(new_n2330_));
  AOI21_X1  g2266(.A(new_n2200_), .B1(new_n2194_), .B2(new_n2198_), .ZN(new_n2331_));
  OAI211_X1 g2267(.A(new_n2327_), .B(new_n2329_), .C1(new_n2330_), .C2(new_n2331_), .ZN(new_n2332_));
  NOR2_X1   g2268(.A1(new_n2331_), .A2(new_n2330_), .ZN(new_n2333_));
  INV_X1    g2269(.A(new_n2329_), .ZN(new_n2334_));
  AOI21_X1  g2270(.A(new_n2328_), .B1(new_n2322_), .B2(new_n2324_), .ZN(new_n2335_));
  OAI21_X1  g2271(.A(new_n2333_), .B1(new_n2334_), .B2(new_n2335_), .ZN(new_n2336_));
  NAND2_X1  g2272(.A1(new_n2332_), .A2(new_n2336_), .ZN(new_n2337_));
  NOR2_X1   g2273(.A1(new_n733_), .A2(new_n980_), .ZN(new_n2338_));
  NAND2_X1  g2274(.A1(new_n2337_), .A2(new_n2338_), .ZN(new_n2339_));
  OAI211_X1 g2275(.A(new_n2332_), .B(new_n2336_), .C1(new_n733_), .C2(new_n980_), .ZN(new_n2340_));
  NAND2_X1  g2276(.A1(new_n2339_), .A2(new_n2340_), .ZN(new_n2341_));
  OAI21_X1  g2277(.A(new_n2203_), .B1(new_n2205_), .B2(new_n2204_), .ZN(new_n2342_));
  NAND2_X1  g2278(.A1(new_n2209_), .A2(new_n2212_), .ZN(new_n2343_));
  NAND3_X1  g2279(.A1(new_n2341_), .A2(new_n2342_), .A3(new_n2343_), .ZN(new_n2344_));
  NAND2_X1  g2280(.A1(new_n2343_), .A2(new_n2342_), .ZN(new_n2345_));
  NAND3_X1  g2281(.A1(new_n2339_), .A2(new_n2340_), .A3(new_n2345_), .ZN(new_n2346_));
  NAND2_X1  g2282(.A1(new_n2344_), .A2(new_n2346_), .ZN(new_n2347_));
  NOR2_X1   g2283(.A1(new_n276_), .A2(new_n1155_), .ZN(new_n2348_));
  NAND2_X1  g2284(.A1(new_n2347_), .A2(new_n2348_), .ZN(new_n2349_));
  INV_X1    g2285(.A(new_n2348_), .ZN(new_n2350_));
  NAND3_X1  g2286(.A1(new_n2344_), .A2(new_n2346_), .A3(new_n2350_), .ZN(new_n2351_));
  NAND2_X1  g2287(.A1(new_n2349_), .A2(new_n2351_), .ZN(new_n2352_));
  NAND2_X1  g2288(.A1(new_n2221_), .A2(new_n2224_), .ZN(new_n2353_));
  NOR2_X1   g2289(.A1(new_n2218_), .A2(new_n2219_), .ZN(new_n2354_));
  OAI21_X1  g2290(.A(new_n2353_), .B1(new_n2354_), .B2(new_n2217_), .ZN(new_n2355_));
  INV_X1    g2291(.A(new_n2355_), .ZN(new_n2356_));
  NAND2_X1  g2292(.A1(new_n2352_), .A2(new_n2356_), .ZN(new_n2357_));
  NAND3_X1  g2293(.A1(new_n2349_), .A2(new_n2351_), .A3(new_n2355_), .ZN(new_n2358_));
  NAND2_X1  g2294(.A1(new_n2357_), .A2(new_n2358_), .ZN(new_n2359_));
  NOR2_X1   g2295(.A1(new_n205_), .A2(new_n1345_), .ZN(new_n2360_));
  NAND2_X1  g2296(.A1(new_n2359_), .A2(new_n2360_), .ZN(new_n2361_));
  INV_X1    g2297(.A(new_n2360_), .ZN(new_n2362_));
  NAND3_X1  g2298(.A1(new_n2357_), .A2(new_n2358_), .A3(new_n2362_), .ZN(new_n2363_));
  NAND2_X1  g2299(.A1(new_n2361_), .A2(new_n2363_), .ZN(new_n2364_));
  NAND2_X1  g2300(.A1(new_n2233_), .A2(new_n2236_), .ZN(new_n2365_));
  NOR2_X1   g2301(.A1(new_n2230_), .A2(new_n2231_), .ZN(new_n2366_));
  OAI21_X1  g2302(.A(new_n2365_), .B1(new_n2366_), .B2(new_n2229_), .ZN(new_n2367_));
  INV_X1    g2303(.A(new_n2367_), .ZN(new_n2368_));
  NAND2_X1  g2304(.A1(new_n2364_), .A2(new_n2368_), .ZN(new_n2369_));
  NAND3_X1  g2305(.A1(new_n2361_), .A2(new_n2363_), .A3(new_n2367_), .ZN(new_n2370_));
  NAND2_X1  g2306(.A1(new_n2369_), .A2(new_n2370_), .ZN(new_n2371_));
  NOR2_X1   g2307(.A1(new_n146_), .A2(new_n1741_), .ZN(new_n2372_));
  NAND2_X1  g2308(.A1(new_n2371_), .A2(new_n2372_), .ZN(new_n2373_));
  INV_X1    g2309(.A(new_n2372_), .ZN(new_n2374_));
  NAND3_X1  g2310(.A1(new_n2369_), .A2(new_n2370_), .A3(new_n2374_), .ZN(new_n2375_));
  NAND2_X1  g2311(.A1(new_n2239_), .A2(new_n2119_), .ZN(new_n2376_));
  INV_X1    g2312(.A(new_n2376_), .ZN(new_n2377_));
  AOI21_X1  g2313(.A(new_n2242_), .B1(new_n2238_), .B2(new_n2240_), .ZN(new_n2378_));
  OAI211_X1 g2314(.A(new_n2373_), .B(new_n2375_), .C1(new_n2377_), .C2(new_n2378_), .ZN(new_n2379_));
  NOR2_X1   g2315(.A1(new_n2378_), .A2(new_n2377_), .ZN(new_n2380_));
  AND3_X1   g2316(.A1(new_n2369_), .A2(new_n2370_), .A3(new_n2374_), .ZN(new_n2381_));
  AOI21_X1  g2317(.A(new_n2374_), .B1(new_n2369_), .B2(new_n2370_), .ZN(new_n2382_));
  OAI21_X1  g2318(.A(new_n2380_), .B1(new_n2381_), .B2(new_n2382_), .ZN(new_n2383_));
  NAND2_X1  g2319(.A1(new_n2379_), .A2(new_n2383_), .ZN(new_n2384_));
  NOR2_X1   g2320(.A1(new_n2250_), .A2(new_n2251_), .ZN(new_n2385_));
  NOR2_X1   g2321(.A1(new_n2385_), .A2(new_n2249_), .ZN(new_n2386_));
  INV_X1    g2322(.A(new_n2386_), .ZN(new_n2387_));
  AOI21_X1  g2323(.A(new_n2384_), .B1(new_n2262_), .B2(new_n2387_), .ZN(new_n2388_));
  AOI21_X1  g2324(.A(new_n2253_), .B1(new_n2114_), .B2(new_n2257_), .ZN(new_n2389_));
  OAI21_X1  g2325(.A(new_n2384_), .B1(new_n2389_), .B2(new_n2386_), .ZN(new_n2390_));
  AOI21_X1  g2326(.A(new_n2388_), .B1(new_n2384_), .B2(new_n2390_), .ZN(G6190gat));
  NAND2_X1  g2327(.A1(new_n2341_), .A2(new_n2345_), .ZN(new_n2392_));
  NAND2_X1  g2328(.A1(new_n2347_), .A2(new_n2350_), .ZN(new_n2393_));
  NAND2_X1  g2329(.A1(new_n2302_), .A2(new_n2305_), .ZN(new_n2394_));
  OAI21_X1  g2330(.A(new_n2299_), .B1(new_n2295_), .B2(new_n2294_), .ZN(new_n2395_));
  NAND2_X1  g2331(.A1(new_n2394_), .A2(new_n2395_), .ZN(new_n2396_));
  INV_X1    g2332(.A(new_n2396_), .ZN(new_n2397_));
  AND2_X1   g2333(.A1(new_n2289_), .A2(new_n2291_), .ZN(new_n2398_));
  NOR2_X1   g2334(.A1(new_n2398_), .A2(new_n2292_), .ZN(new_n2399_));
  INV_X1    g2335(.A(new_n2399_), .ZN(new_n2400_));
  NOR2_X1   g2336(.A1(new_n1041_), .A2(new_n432_), .ZN(new_n2401_));
  NAND2_X1  g2337(.A1(new_n2280_), .A2(new_n2281_), .ZN(new_n2402_));
  NAND2_X1  g2338(.A1(new_n2402_), .A2(new_n2277_), .ZN(new_n2403_));
  NOR2_X1   g2339(.A1(new_n1805_), .A2(new_n253_), .ZN(new_n2404_));
  INV_X1    g2340(.A(new_n2404_), .ZN(new_n2405_));
  NAND2_X1  g2341(.A1(new_n2403_), .A2(new_n2405_), .ZN(new_n2406_));
  NAND2_X1  g2342(.A1(new_n2406_), .A2(new_n2405_), .ZN(new_n2407_));
  NAND2_X1  g2343(.A1(new_n2403_), .A2(new_n2404_), .ZN(new_n2408_));
  NAND2_X1  g2344(.A1(new_n2407_), .A2(new_n2408_), .ZN(new_n2409_));
  NOR2_X1   g2345(.A1(new_n1220_), .A2(new_n336_), .ZN(new_n2410_));
  NOR2_X1   g2346(.A1(new_n2409_), .A2(new_n2410_), .ZN(new_n2411_));
  INV_X1    g2347(.A(new_n2410_), .ZN(new_n2412_));
  AOI21_X1  g2348(.A(new_n2412_), .B1(new_n2407_), .B2(new_n2408_), .ZN(new_n2413_));
  NOR2_X1   g2349(.A1(new_n2411_), .A2(new_n2413_), .ZN(new_n2414_));
  OAI21_X1  g2350(.A(new_n2268_), .B1(new_n2287_), .B2(new_n2283_), .ZN(new_n2415_));
  INV_X1    g2351(.A(new_n2282_), .ZN(new_n2416_));
  NAND2_X1  g2352(.A1(new_n2416_), .A2(new_n2271_), .ZN(new_n2417_));
  NAND2_X1  g2353(.A1(new_n2415_), .A2(new_n2417_), .ZN(new_n2418_));
  NAND2_X1  g2354(.A1(new_n2414_), .A2(new_n2418_), .ZN(new_n2419_));
  INV_X1    g2355(.A(new_n2419_), .ZN(new_n2420_));
  NOR2_X1   g2356(.A1(new_n2414_), .A2(new_n2418_), .ZN(new_n2421_));
  OAI21_X1  g2357(.A(new_n2401_), .B1(new_n2420_), .B2(new_n2421_), .ZN(new_n2422_));
  INV_X1    g2358(.A(new_n2421_), .ZN(new_n2423_));
  INV_X1    g2359(.A(new_n2401_), .ZN(new_n2424_));
  NAND3_X1  g2360(.A1(new_n2423_), .A2(new_n2419_), .A3(new_n2424_), .ZN(new_n2425_));
  NAND2_X1  g2361(.A1(new_n2422_), .A2(new_n2425_), .ZN(new_n2426_));
  NOR2_X1   g2362(.A1(new_n2266_), .A2(new_n2290_), .ZN(new_n2427_));
  INV_X1    g2363(.A(new_n2427_), .ZN(new_n2428_));
  NAND3_X1  g2364(.A1(new_n2400_), .A2(new_n2426_), .A3(new_n2428_), .ZN(new_n2429_));
  INV_X1    g2365(.A(new_n2426_), .ZN(new_n2430_));
  OAI21_X1  g2366(.A(new_n2430_), .B1(new_n2399_), .B2(new_n2427_), .ZN(new_n2431_));
  NAND2_X1  g2367(.A1(new_n2429_), .A2(new_n2431_), .ZN(new_n2432_));
  NOR2_X1   g2368(.A1(new_n873_), .A2(new_n544_), .ZN(new_n2433_));
  NAND2_X1  g2369(.A1(new_n2432_), .A2(new_n2433_), .ZN(new_n2434_));
  OAI211_X1 g2370(.A(new_n2429_), .B(new_n2431_), .C1(new_n873_), .C2(new_n544_), .ZN(new_n2435_));
  NAND2_X1  g2371(.A1(new_n2434_), .A2(new_n2435_), .ZN(new_n2436_));
  NAND2_X1  g2372(.A1(new_n2397_), .A2(new_n2436_), .ZN(new_n2437_));
  AND2_X1   g2373(.A1(new_n2434_), .A2(new_n2435_), .ZN(new_n2438_));
  NAND2_X1  g2374(.A1(new_n2438_), .A2(new_n2396_), .ZN(new_n2439_));
  NOR2_X1   g2375(.A1(new_n719_), .A2(new_n673_), .ZN(new_n2440_));
  INV_X1    g2376(.A(new_n2440_), .ZN(new_n2441_));
  AND3_X1   g2377(.A1(new_n2437_), .A2(new_n2439_), .A3(new_n2441_), .ZN(new_n2442_));
  AOI21_X1  g2378(.A(new_n2441_), .B1(new_n2437_), .B2(new_n2439_), .ZN(new_n2443_));
  NOR2_X1   g2379(.A1(new_n2442_), .A2(new_n2443_), .ZN(new_n2444_));
  AOI21_X1  g2380(.A(new_n2314_), .B1(new_n2311_), .B2(new_n2312_), .ZN(new_n2445_));
  AOI21_X1  g2381(.A(new_n2310_), .B1(new_n2304_), .B2(new_n2306_), .ZN(new_n2446_));
  NOR2_X1   g2382(.A1(new_n2445_), .A2(new_n2446_), .ZN(new_n2447_));
  INV_X1    g2383(.A(new_n2447_), .ZN(new_n2448_));
  NAND2_X1  g2384(.A1(new_n2444_), .A2(new_n2448_), .ZN(new_n2449_));
  OAI21_X1  g2385(.A(new_n2447_), .B1(new_n2442_), .B2(new_n2443_), .ZN(new_n2450_));
  NAND2_X1  g2386(.A1(G171gat), .A2(G460gat), .ZN(new_n2451_));
  AND3_X1   g2387(.A1(new_n2449_), .A2(new_n2450_), .A3(new_n2451_), .ZN(new_n2452_));
  AOI21_X1  g2388(.A(new_n2451_), .B1(new_n2449_), .B2(new_n2450_), .ZN(new_n2453_));
  NOR2_X1   g2389(.A1(new_n2452_), .A2(new_n2453_), .ZN(new_n2454_));
  AOI21_X1  g2390(.A(new_n2321_), .B1(new_n2315_), .B2(new_n2316_), .ZN(new_n2455_));
  AOI21_X1  g2391(.A(new_n2326_), .B1(new_n2322_), .B2(new_n2324_), .ZN(new_n2456_));
  OAI21_X1  g2392(.A(new_n2454_), .B1(new_n2455_), .B2(new_n2456_), .ZN(new_n2457_));
  NOR2_X1   g2393(.A1(new_n2456_), .A2(new_n2455_), .ZN(new_n2458_));
  OAI21_X1  g2394(.A(new_n2458_), .B1(new_n2452_), .B2(new_n2453_), .ZN(new_n2459_));
  NAND2_X1  g2395(.A1(new_n2457_), .A2(new_n2459_), .ZN(new_n2460_));
  NOR2_X1   g2396(.A1(new_n889_), .A2(new_n980_), .ZN(new_n2461_));
  NAND2_X1  g2397(.A1(new_n2460_), .A2(new_n2461_), .ZN(new_n2462_));
  INV_X1    g2398(.A(new_n2461_), .ZN(new_n2463_));
  NAND3_X1  g2399(.A1(new_n2457_), .A2(new_n2459_), .A3(new_n2463_), .ZN(new_n2464_));
  NAND2_X1  g2400(.A1(new_n2462_), .A2(new_n2464_), .ZN(new_n2465_));
  AOI21_X1  g2401(.A(new_n2338_), .B1(new_n2332_), .B2(new_n2336_), .ZN(new_n2466_));
  AOI21_X1  g2402(.A(new_n2333_), .B1(new_n2327_), .B2(new_n2329_), .ZN(new_n2467_));
  NOR2_X1   g2403(.A1(new_n2466_), .A2(new_n2467_), .ZN(new_n2468_));
  NAND2_X1  g2404(.A1(new_n2465_), .A2(new_n2468_), .ZN(new_n2469_));
  OAI211_X1 g2405(.A(new_n2462_), .B(new_n2464_), .C1(new_n2467_), .C2(new_n2466_), .ZN(new_n2470_));
  NOR2_X1   g2406(.A1(new_n733_), .A2(new_n1155_), .ZN(new_n2471_));
  INV_X1    g2407(.A(new_n2471_), .ZN(new_n2472_));
  AND3_X1   g2408(.A1(new_n2469_), .A2(new_n2470_), .A3(new_n2472_), .ZN(new_n2473_));
  AOI21_X1  g2409(.A(new_n2472_), .B1(new_n2469_), .B2(new_n2470_), .ZN(new_n2474_));
  OAI211_X1 g2410(.A(new_n2392_), .B(new_n2393_), .C1(new_n2473_), .C2(new_n2474_), .ZN(new_n2475_));
  INV_X1    g2411(.A(new_n2474_), .ZN(new_n2476_));
  NAND2_X1  g2412(.A1(new_n2393_), .A2(new_n2392_), .ZN(new_n2477_));
  NAND3_X1  g2413(.A1(new_n2469_), .A2(new_n2470_), .A3(new_n2472_), .ZN(new_n2478_));
  NAND3_X1  g2414(.A1(new_n2476_), .A2(new_n2477_), .A3(new_n2478_), .ZN(new_n2479_));
  NAND2_X1  g2415(.A1(new_n2475_), .A2(new_n2479_), .ZN(new_n2480_));
  INV_X1    g2416(.A(new_n2480_), .ZN(new_n2481_));
  NOR2_X1   g2417(.A1(new_n276_), .A2(new_n1345_), .ZN(new_n2482_));
  INV_X1    g2418(.A(new_n2482_), .ZN(new_n2483_));
  NAND2_X1  g2419(.A1(new_n2481_), .A2(new_n2483_), .ZN(new_n2484_));
  AOI21_X1  g2420(.A(new_n2483_), .B1(new_n2475_), .B2(new_n2479_), .ZN(new_n2485_));
  INV_X1    g2421(.A(new_n2485_), .ZN(new_n2486_));
  NAND2_X1  g2422(.A1(new_n2359_), .A2(new_n2362_), .ZN(new_n2487_));
  NAND2_X1  g2423(.A1(new_n2352_), .A2(new_n2355_), .ZN(new_n2488_));
  NAND2_X1  g2424(.A1(new_n2487_), .A2(new_n2488_), .ZN(new_n2489_));
  NAND3_X1  g2425(.A1(new_n2484_), .A2(new_n2486_), .A3(new_n2489_), .ZN(new_n2490_));
  NOR2_X1   g2426(.A1(new_n2480_), .A2(new_n2482_), .ZN(new_n2491_));
  OAI211_X1 g2427(.A(new_n2488_), .B(new_n2487_), .C1(new_n2491_), .C2(new_n2485_), .ZN(new_n2492_));
  NAND2_X1  g2428(.A1(new_n2490_), .A2(new_n2492_), .ZN(new_n2493_));
  NOR2_X1   g2429(.A1(new_n205_), .A2(new_n1741_), .ZN(new_n2494_));
  NAND2_X1  g2430(.A1(new_n2493_), .A2(new_n2494_), .ZN(new_n2495_));
  NAND2_X1  g2431(.A1(new_n2371_), .A2(new_n2374_), .ZN(new_n2496_));
  NAND2_X1  g2432(.A1(new_n2364_), .A2(new_n2367_), .ZN(new_n2497_));
  NAND2_X1  g2433(.A1(new_n2496_), .A2(new_n2497_), .ZN(new_n2498_));
  AOI21_X1  g2434(.A(new_n2494_), .B1(new_n2490_), .B2(new_n2492_), .ZN(new_n2499_));
  OAI211_X1 g2435(.A(new_n2495_), .B(new_n2498_), .C1(new_n2494_), .C2(new_n2499_), .ZN(new_n2500_));
  INV_X1    g2436(.A(new_n2494_), .ZN(new_n2501_));
  AND3_X1   g2437(.A1(new_n2490_), .A2(new_n2492_), .A3(new_n2501_), .ZN(new_n2502_));
  AOI21_X1  g2438(.A(new_n2501_), .B1(new_n2490_), .B2(new_n2492_), .ZN(new_n2503_));
  OAI211_X1 g2439(.A(new_n2497_), .B(new_n2496_), .C1(new_n2502_), .C2(new_n2503_), .ZN(new_n2504_));
  AND2_X1   g2440(.A1(new_n2500_), .A2(new_n2504_), .ZN(new_n2505_));
  INV_X1    g2441(.A(new_n2505_), .ZN(new_n2506_));
  NOR2_X1   g2442(.A1(new_n2381_), .A2(new_n2382_), .ZN(new_n2507_));
  NOR2_X1   g2443(.A1(new_n2507_), .A2(new_n2380_), .ZN(new_n2508_));
  INV_X1    g2444(.A(new_n2508_), .ZN(new_n2509_));
  AOI21_X1  g2445(.A(new_n2506_), .B1(new_n2390_), .B2(new_n2509_), .ZN(new_n2510_));
  AND2_X1   g2446(.A1(new_n2379_), .A2(new_n2383_), .ZN(new_n2511_));
  AOI21_X1  g2447(.A(new_n2511_), .B1(new_n2262_), .B2(new_n2387_), .ZN(new_n2512_));
  OAI21_X1  g2448(.A(new_n2506_), .B1(new_n2512_), .B2(new_n2508_), .ZN(new_n2513_));
  AOI21_X1  g2449(.A(new_n2510_), .B1(new_n2513_), .B2(new_n2506_), .ZN(G6200gat));
  AOI21_X1  g2450(.A(new_n2505_), .B1(new_n2390_), .B2(new_n2509_), .ZN(new_n2515_));
  OAI21_X1  g2451(.A(new_n2498_), .B1(new_n2502_), .B2(new_n2503_), .ZN(new_n2516_));
  INV_X1    g2452(.A(new_n2516_), .ZN(new_n2517_));
  NOR2_X1   g2453(.A1(new_n2515_), .A2(new_n2517_), .ZN(new_n2518_));
  NOR2_X1   g2454(.A1(new_n876_), .A2(new_n980_), .ZN(new_n2519_));
  NAND2_X1  g2455(.A1(new_n2409_), .A2(new_n2412_), .ZN(new_n2520_));
  NAND2_X1  g2456(.A1(new_n2520_), .A2(new_n2406_), .ZN(new_n2521_));
  NOR2_X1   g2457(.A1(new_n1805_), .A2(new_n336_), .ZN(new_n2522_));
  OR2_X1    g2458(.A1(new_n2521_), .A2(new_n2522_), .ZN(new_n2523_));
  NAND2_X1  g2459(.A1(new_n2521_), .A2(new_n2522_), .ZN(new_n2524_));
  NAND2_X1  g2460(.A1(new_n2523_), .A2(new_n2524_), .ZN(new_n2525_));
  AOI21_X1  g2461(.A(new_n2525_), .B1(G239gat), .B2(G409gat), .ZN(new_n2526_));
  NAND2_X1  g2462(.A1(G239gat), .A2(G409gat), .ZN(new_n2527_));
  AOI21_X1  g2463(.A(new_n2527_), .B1(new_n2523_), .B2(new_n2524_), .ZN(new_n2528_));
  NOR2_X1   g2464(.A1(new_n2526_), .A2(new_n2528_), .ZN(new_n2529_));
  INV_X1    g2465(.A(new_n2414_), .ZN(new_n2530_));
  NAND2_X1  g2466(.A1(new_n2530_), .A2(new_n2418_), .ZN(new_n2531_));
  INV_X1    g2467(.A(new_n2531_), .ZN(new_n2532_));
  AOI21_X1  g2468(.A(new_n2401_), .B1(new_n2423_), .B2(new_n2419_), .ZN(new_n2533_));
  OAI21_X1  g2469(.A(new_n2529_), .B1(new_n2532_), .B2(new_n2533_), .ZN(new_n2534_));
  INV_X1    g2470(.A(new_n2533_), .ZN(new_n2535_));
  OAI211_X1 g2471(.A(new_n2535_), .B(new_n2531_), .C1(new_n2526_), .C2(new_n2528_), .ZN(new_n2536_));
  NAND2_X1  g2472(.A1(G222gat), .A2(G426gat), .ZN(new_n2537_));
  NAND3_X1  g2473(.A1(new_n2534_), .A2(new_n2536_), .A3(new_n2537_), .ZN(new_n2538_));
  INV_X1    g2474(.A(new_n2538_), .ZN(new_n2539_));
  AOI21_X1  g2475(.A(new_n2537_), .B1(new_n2534_), .B2(new_n2536_), .ZN(new_n2540_));
  NOR2_X1   g2476(.A1(new_n2539_), .A2(new_n2540_), .ZN(new_n2541_));
  AOI21_X1  g2477(.A(new_n2430_), .B1(new_n2400_), .B2(new_n2428_), .ZN(new_n2542_));
  AOI21_X1  g2478(.A(new_n2433_), .B1(new_n2429_), .B2(new_n2431_), .ZN(new_n2543_));
  OAI21_X1  g2479(.A(new_n2541_), .B1(new_n2542_), .B2(new_n2543_), .ZN(new_n2544_));
  NOR2_X1   g2480(.A1(new_n2543_), .A2(new_n2542_), .ZN(new_n2545_));
  OAI21_X1  g2481(.A(new_n2545_), .B1(new_n2540_), .B2(new_n2539_), .ZN(new_n2546_));
  NAND2_X1  g2482(.A1(new_n2544_), .A2(new_n2546_), .ZN(new_n2547_));
  NOR2_X1   g2483(.A1(new_n873_), .A2(new_n673_), .ZN(new_n2548_));
  NAND2_X1  g2484(.A1(new_n2547_), .A2(new_n2548_), .ZN(new_n2549_));
  AOI21_X1  g2485(.A(new_n2548_), .B1(new_n2544_), .B2(new_n2546_), .ZN(new_n2550_));
  OAI21_X1  g2486(.A(new_n2549_), .B1(new_n2548_), .B2(new_n2550_), .ZN(new_n2551_));
  INV_X1    g2487(.A(new_n2551_), .ZN(new_n2552_));
  NOR2_X1   g2488(.A1(new_n2397_), .A2(new_n2438_), .ZN(new_n2553_));
  AOI21_X1  g2489(.A(new_n2440_), .B1(new_n2437_), .B2(new_n2439_), .ZN(new_n2554_));
  OAI21_X1  g2490(.A(new_n2552_), .B1(new_n2553_), .B2(new_n2554_), .ZN(new_n2555_));
  INV_X1    g2491(.A(new_n2554_), .ZN(new_n2556_));
  INV_X1    g2492(.A(new_n2553_), .ZN(new_n2557_));
  NAND3_X1  g2493(.A1(new_n2551_), .A2(new_n2556_), .A3(new_n2557_), .ZN(new_n2558_));
  NAND2_X1  g2494(.A1(new_n2555_), .A2(new_n2558_), .ZN(new_n2559_));
  NOR2_X1   g2495(.A1(new_n719_), .A2(new_n816_), .ZN(new_n2560_));
  NAND2_X1  g2496(.A1(new_n2559_), .A2(new_n2560_), .ZN(new_n2561_));
  AOI21_X1  g2497(.A(new_n2560_), .B1(new_n2555_), .B2(new_n2558_), .ZN(new_n2562_));
  OAI21_X1  g2498(.A(new_n2561_), .B1(new_n2560_), .B2(new_n2562_), .ZN(new_n2563_));
  AOI22_X1  g2499(.A1(new_n2449_), .A2(new_n2450_), .B1(G171gat), .B2(G460gat), .ZN(new_n2564_));
  NOR2_X1   g2500(.A1(new_n2444_), .A2(new_n2447_), .ZN(new_n2565_));
  NOR2_X1   g2501(.A1(new_n2564_), .A2(new_n2565_), .ZN(new_n2566_));
  NOR2_X1   g2502(.A1(new_n2563_), .A2(new_n2566_), .ZN(new_n2567_));
  INV_X1    g2503(.A(new_n2560_), .ZN(new_n2568_));
  AND3_X1   g2504(.A1(new_n2555_), .A2(new_n2558_), .A3(new_n2568_), .ZN(new_n2569_));
  AOI21_X1  g2505(.A(new_n2568_), .B1(new_n2555_), .B2(new_n2558_), .ZN(new_n2570_));
  NOR2_X1   g2506(.A1(new_n2569_), .A2(new_n2570_), .ZN(new_n2571_));
  INV_X1    g2507(.A(new_n2566_), .ZN(new_n2572_));
  NOR2_X1   g2508(.A1(new_n2571_), .A2(new_n2572_), .ZN(new_n2573_));
  OAI21_X1  g2509(.A(new_n2519_), .B1(new_n2567_), .B2(new_n2573_), .ZN(new_n2574_));
  NAND2_X1  g2510(.A1(new_n2563_), .A2(new_n2566_), .ZN(new_n2575_));
  NAND2_X1  g2511(.A1(new_n2571_), .A2(new_n2572_), .ZN(new_n2576_));
  INV_X1    g2512(.A(new_n2519_), .ZN(new_n2577_));
  NAND3_X1  g2513(.A1(new_n2575_), .A2(new_n2576_), .A3(new_n2577_), .ZN(new_n2578_));
  NAND2_X1  g2514(.A1(new_n2574_), .A2(new_n2578_), .ZN(new_n2579_));
  NOR2_X1   g2515(.A1(new_n2454_), .A2(new_n2458_), .ZN(new_n2580_));
  INV_X1    g2516(.A(new_n2580_), .ZN(new_n2581_));
  NAND2_X1  g2517(.A1(new_n2460_), .A2(new_n2463_), .ZN(new_n2582_));
  NAND3_X1  g2518(.A1(new_n2579_), .A2(new_n2581_), .A3(new_n2582_), .ZN(new_n2583_));
  NAND2_X1  g2519(.A1(new_n2582_), .A2(new_n2581_), .ZN(new_n2584_));
  NAND3_X1  g2520(.A1(new_n2584_), .A2(new_n2574_), .A3(new_n2578_), .ZN(new_n2585_));
  NAND2_X1  g2521(.A1(new_n2583_), .A2(new_n2585_), .ZN(new_n2586_));
  NOR2_X1   g2522(.A1(new_n889_), .A2(new_n1155_), .ZN(new_n2587_));
  NAND2_X1  g2523(.A1(new_n2586_), .A2(new_n2587_), .ZN(new_n2588_));
  INV_X1    g2524(.A(new_n2587_), .ZN(new_n2589_));
  NAND3_X1  g2525(.A1(new_n2583_), .A2(new_n2585_), .A3(new_n2589_), .ZN(new_n2590_));
  NAND2_X1  g2526(.A1(new_n2588_), .A2(new_n2590_), .ZN(new_n2591_));
  AOI21_X1  g2527(.A(new_n2471_), .B1(new_n2469_), .B2(new_n2470_), .ZN(new_n2592_));
  AOI21_X1  g2528(.A(new_n2468_), .B1(new_n2462_), .B2(new_n2464_), .ZN(new_n2593_));
  NOR2_X1   g2529(.A1(new_n2592_), .A2(new_n2593_), .ZN(new_n2594_));
  NAND2_X1  g2530(.A1(new_n2591_), .A2(new_n2594_), .ZN(new_n2595_));
  OAI211_X1 g2531(.A(new_n2588_), .B(new_n2590_), .C1(new_n2593_), .C2(new_n2592_), .ZN(new_n2596_));
  NAND2_X1  g2532(.A1(new_n2595_), .A2(new_n2596_), .ZN(new_n2597_));
  NOR2_X1   g2533(.A1(new_n733_), .A2(new_n1345_), .ZN(new_n2598_));
  NAND2_X1  g2534(.A1(new_n2597_), .A2(new_n2598_), .ZN(new_n2599_));
  INV_X1    g2535(.A(new_n2598_), .ZN(new_n2600_));
  NAND3_X1  g2536(.A1(new_n2595_), .A2(new_n2596_), .A3(new_n2600_), .ZN(new_n2601_));
  NAND2_X1  g2537(.A1(new_n2599_), .A2(new_n2601_), .ZN(new_n2602_));
  NOR2_X1   g2538(.A1(new_n2481_), .A2(new_n2482_), .ZN(new_n2603_));
  AOI22_X1  g2539(.A1(new_n2476_), .A2(new_n2478_), .B1(new_n2392_), .B2(new_n2393_), .ZN(new_n2604_));
  NOR2_X1   g2540(.A1(new_n2603_), .A2(new_n2604_), .ZN(new_n2605_));
  NAND2_X1  g2541(.A1(new_n2602_), .A2(new_n2605_), .ZN(new_n2606_));
  OAI211_X1 g2542(.A(new_n2599_), .B(new_n2601_), .C1(new_n2604_), .C2(new_n2603_), .ZN(new_n2607_));
  NAND2_X1  g2543(.A1(new_n2606_), .A2(new_n2607_), .ZN(new_n2608_));
  NOR2_X1   g2544(.A1(new_n276_), .A2(new_n1741_), .ZN(new_n2609_));
  NAND2_X1  g2545(.A1(new_n2608_), .A2(new_n2609_), .ZN(new_n2610_));
  OAI211_X1 g2546(.A(new_n2606_), .B(new_n2607_), .C1(new_n276_), .C2(new_n1741_), .ZN(new_n2611_));
  NAND2_X1  g2547(.A1(new_n2610_), .A2(new_n2611_), .ZN(new_n2612_));
  OAI21_X1  g2548(.A(new_n2489_), .B1(new_n2491_), .B2(new_n2485_), .ZN(new_n2613_));
  INV_X1    g2549(.A(new_n2613_), .ZN(new_n2614_));
  NOR2_X1   g2550(.A1(new_n2499_), .A2(new_n2614_), .ZN(new_n2615_));
  NAND2_X1  g2551(.A1(new_n2612_), .A2(new_n2615_), .ZN(new_n2616_));
  OAI211_X1 g2552(.A(new_n2610_), .B(new_n2611_), .C1(new_n2614_), .C2(new_n2499_), .ZN(new_n2617_));
  NAND2_X1  g2553(.A1(new_n2616_), .A2(new_n2617_), .ZN(new_n2618_));
  INV_X1    g2554(.A(new_n2618_), .ZN(new_n2619_));
  XNOR2_X1  g2555(.A(new_n2518_), .B(new_n2619_), .ZN(G6210gat));
  NOR2_X1   g2556(.A1(new_n719_), .A2(new_n980_), .ZN(new_n2621_));
  AOI22_X1  g2557(.A1(new_n2534_), .A2(new_n2536_), .B1(G222gat), .B2(G426gat), .ZN(new_n2622_));
  AOI21_X1  g2558(.A(new_n2529_), .B1(new_n2531_), .B2(new_n2535_), .ZN(new_n2623_));
  NOR2_X1   g2559(.A1(new_n2622_), .A2(new_n2623_), .ZN(new_n2624_));
  INV_X1    g2560(.A(new_n2624_), .ZN(new_n2625_));
  NAND2_X1  g2561(.A1(new_n2525_), .A2(new_n2527_), .ZN(new_n2626_));
  AOI21_X1  g2562(.A(new_n2522_), .B1(new_n2520_), .B2(new_n2406_), .ZN(new_n2627_));
  INV_X1    g2563(.A(new_n2627_), .ZN(new_n2628_));
  NAND2_X1  g2564(.A1(new_n2626_), .A2(new_n2628_), .ZN(new_n2629_));
  NOR2_X1   g2565(.A1(new_n1805_), .A2(new_n432_), .ZN(new_n2630_));
  INV_X1    g2566(.A(new_n2630_), .ZN(new_n2631_));
  NAND2_X1  g2567(.A1(new_n2629_), .A2(new_n2631_), .ZN(new_n2632_));
  NAND2_X1  g2568(.A1(new_n2632_), .A2(new_n2631_), .ZN(new_n2633_));
  NAND2_X1  g2569(.A1(new_n2629_), .A2(new_n2630_), .ZN(new_n2634_));
  NAND2_X1  g2570(.A1(G239gat), .A2(G426gat), .ZN(new_n2635_));
  AND3_X1   g2571(.A1(new_n2633_), .A2(new_n2634_), .A3(new_n2635_), .ZN(new_n2636_));
  AOI21_X1  g2572(.A(new_n2635_), .B1(new_n2633_), .B2(new_n2634_), .ZN(new_n2637_));
  NOR2_X1   g2573(.A1(new_n2636_), .A2(new_n2637_), .ZN(new_n2638_));
  NAND2_X1  g2574(.A1(new_n2625_), .A2(new_n2638_), .ZN(new_n2639_));
  INV_X1    g2575(.A(new_n2638_), .ZN(new_n2640_));
  NAND2_X1  g2576(.A1(new_n2640_), .A2(new_n2624_), .ZN(new_n2641_));
  NAND2_X1  g2577(.A1(new_n2639_), .A2(new_n2641_), .ZN(new_n2642_));
  NAND2_X1  g2578(.A1(G222gat), .A2(G443gat), .ZN(new_n2643_));
  XNOR2_X1  g2579(.A(new_n2642_), .B(new_n2643_), .ZN(new_n2644_));
  INV_X1    g2580(.A(new_n2644_), .ZN(new_n2645_));
  NOR2_X1   g2581(.A1(new_n2541_), .A2(new_n2545_), .ZN(new_n2646_));
  NOR2_X1   g2582(.A1(new_n2550_), .A2(new_n2646_), .ZN(new_n2647_));
  NAND2_X1  g2583(.A1(new_n2645_), .A2(new_n2647_), .ZN(new_n2648_));
  OAI21_X1  g2584(.A(new_n2644_), .B1(new_n2646_), .B2(new_n2550_), .ZN(new_n2649_));
  NOR2_X1   g2585(.A1(new_n873_), .A2(new_n816_), .ZN(new_n2650_));
  INV_X1    g2586(.A(new_n2650_), .ZN(new_n2651_));
  AND3_X1   g2587(.A1(new_n2648_), .A2(new_n2649_), .A3(new_n2651_), .ZN(new_n2652_));
  AOI21_X1  g2588(.A(new_n2651_), .B1(new_n2648_), .B2(new_n2649_), .ZN(new_n2653_));
  OR2_X1    g2589(.A1(new_n2652_), .A2(new_n2653_), .ZN(new_n2654_));
  AOI21_X1  g2590(.A(new_n2552_), .B1(new_n2557_), .B2(new_n2556_), .ZN(new_n2655_));
  NOR2_X1   g2591(.A1(new_n2562_), .A2(new_n2655_), .ZN(new_n2656_));
  NOR2_X1   g2592(.A1(new_n2654_), .A2(new_n2656_), .ZN(new_n2657_));
  OR2_X1    g2593(.A1(new_n2562_), .A2(new_n2655_), .ZN(new_n2658_));
  NOR2_X1   g2594(.A1(new_n2652_), .A2(new_n2653_), .ZN(new_n2659_));
  NOR2_X1   g2595(.A1(new_n2658_), .A2(new_n2659_), .ZN(new_n2660_));
  OAI21_X1  g2596(.A(new_n2621_), .B1(new_n2657_), .B2(new_n2660_), .ZN(new_n2661_));
  NAND2_X1  g2597(.A1(new_n2654_), .A2(new_n2656_), .ZN(new_n2662_));
  NAND2_X1  g2598(.A1(new_n2658_), .A2(new_n2659_), .ZN(new_n2663_));
  AOI21_X1  g2599(.A(new_n2621_), .B1(new_n2662_), .B2(new_n2663_), .ZN(new_n2664_));
  OAI21_X1  g2600(.A(new_n2661_), .B1(new_n2664_), .B2(new_n2621_), .ZN(new_n2665_));
  NAND2_X1  g2601(.A1(new_n2563_), .A2(new_n2572_), .ZN(new_n2666_));
  OAI21_X1  g2602(.A(new_n2577_), .B1(new_n2567_), .B2(new_n2573_), .ZN(new_n2667_));
  NAND3_X1  g2603(.A1(new_n2665_), .A2(new_n2666_), .A3(new_n2667_), .ZN(new_n2668_));
  INV_X1    g2604(.A(new_n2621_), .ZN(new_n2669_));
  AOI21_X1  g2605(.A(new_n2669_), .B1(new_n2662_), .B2(new_n2663_), .ZN(new_n2670_));
  OAI21_X1  g2606(.A(new_n2669_), .B1(new_n2657_), .B2(new_n2660_), .ZN(new_n2671_));
  AOI21_X1  g2607(.A(new_n2670_), .B1(new_n2671_), .B2(new_n2669_), .ZN(new_n2672_));
  NAND2_X1  g2608(.A1(new_n2667_), .A2(new_n2666_), .ZN(new_n2673_));
  NAND2_X1  g2609(.A1(new_n2672_), .A2(new_n2673_), .ZN(new_n2674_));
  NOR2_X1   g2610(.A1(new_n876_), .A2(new_n1155_), .ZN(new_n2675_));
  INV_X1    g2611(.A(new_n2675_), .ZN(new_n2676_));
  NAND3_X1  g2612(.A1(new_n2668_), .A2(new_n2674_), .A3(new_n2676_), .ZN(new_n2677_));
  INV_X1    g2613(.A(new_n2677_), .ZN(new_n2678_));
  NAND2_X1  g2614(.A1(new_n2579_), .A2(new_n2584_), .ZN(new_n2679_));
  INV_X1    g2615(.A(new_n2679_), .ZN(new_n2680_));
  AOI21_X1  g2616(.A(new_n2680_), .B1(new_n2586_), .B2(new_n2589_), .ZN(new_n2681_));
  AOI21_X1  g2617(.A(new_n2676_), .B1(new_n2668_), .B2(new_n2674_), .ZN(new_n2682_));
  NOR3_X1   g2618(.A1(new_n2678_), .A2(new_n2681_), .A3(new_n2682_), .ZN(new_n2683_));
  INV_X1    g2619(.A(new_n2683_), .ZN(new_n2684_));
  NOR2_X1   g2620(.A1(new_n889_), .A2(new_n1345_), .ZN(new_n2685_));
  INV_X1    g2621(.A(new_n2685_), .ZN(new_n2686_));
  NOR2_X1   g2622(.A1(new_n2678_), .A2(new_n2682_), .ZN(new_n2687_));
  NOR2_X1   g2623(.A1(new_n2687_), .A2(new_n2681_), .ZN(new_n2688_));
  OAI211_X1 g2624(.A(new_n2684_), .B(new_n2686_), .C1(new_n2688_), .C2(new_n2687_), .ZN(new_n2689_));
  INV_X1    g2625(.A(new_n2681_), .ZN(new_n2690_));
  NOR2_X1   g2626(.A1(new_n2687_), .A2(new_n2690_), .ZN(new_n2691_));
  OAI21_X1  g2627(.A(new_n2685_), .B1(new_n2691_), .B2(new_n2683_), .ZN(new_n2692_));
  NAND2_X1  g2628(.A1(new_n2689_), .A2(new_n2692_), .ZN(new_n2693_));
  NAND2_X1  g2629(.A1(new_n2597_), .A2(new_n2600_), .ZN(new_n2694_));
  OAI21_X1  g2630(.A(new_n2591_), .B1(new_n2593_), .B2(new_n2592_), .ZN(new_n2695_));
  NAND2_X1  g2631(.A1(new_n2694_), .A2(new_n2695_), .ZN(new_n2696_));
  INV_X1    g2632(.A(new_n2696_), .ZN(new_n2697_));
  NAND2_X1  g2633(.A1(new_n2693_), .A2(new_n2697_), .ZN(new_n2698_));
  NAND3_X1  g2634(.A1(new_n2696_), .A2(new_n2689_), .A3(new_n2692_), .ZN(new_n2699_));
  NAND2_X1  g2635(.A1(new_n2698_), .A2(new_n2699_), .ZN(new_n2700_));
  NOR2_X1   g2636(.A1(new_n733_), .A2(new_n1741_), .ZN(new_n2701_));
  NAND2_X1  g2637(.A1(new_n2700_), .A2(new_n2701_), .ZN(new_n2702_));
  OAI211_X1 g2638(.A(new_n2698_), .B(new_n2699_), .C1(new_n733_), .C2(new_n1741_), .ZN(new_n2703_));
  NAND2_X1  g2639(.A1(new_n2702_), .A2(new_n2703_), .ZN(new_n2704_));
  AOI21_X1  g2640(.A(new_n2609_), .B1(new_n2606_), .B2(new_n2607_), .ZN(new_n2705_));
  AOI21_X1  g2641(.A(new_n2605_), .B1(new_n2599_), .B2(new_n2601_), .ZN(new_n2706_));
  NOR2_X1   g2642(.A1(new_n2705_), .A2(new_n2706_), .ZN(new_n2707_));
  NAND2_X1  g2643(.A1(new_n2704_), .A2(new_n2707_), .ZN(new_n2708_));
  OAI211_X1 g2644(.A(new_n2702_), .B(new_n2703_), .C1(new_n2706_), .C2(new_n2705_), .ZN(new_n2709_));
  NAND2_X1  g2645(.A1(new_n2708_), .A2(new_n2709_), .ZN(new_n2710_));
  OAI21_X1  g2646(.A(new_n2618_), .B1(new_n2515_), .B2(new_n2517_), .ZN(new_n2711_));
  AOI21_X1  g2647(.A(new_n2615_), .B1(new_n2610_), .B2(new_n2611_), .ZN(new_n2712_));
  INV_X1    g2648(.A(new_n2712_), .ZN(new_n2713_));
  AOI21_X1  g2649(.A(new_n2710_), .B1(new_n2711_), .B2(new_n2713_), .ZN(new_n2714_));
  AOI21_X1  g2650(.A(new_n2619_), .B1(new_n2513_), .B2(new_n2516_), .ZN(new_n2715_));
  OAI21_X1  g2651(.A(new_n2710_), .B1(new_n2715_), .B2(new_n2712_), .ZN(new_n2716_));
  AOI21_X1  g2652(.A(new_n2714_), .B1(new_n2716_), .B2(new_n2710_), .ZN(G6220gat));
  INV_X1    g2653(.A(new_n2710_), .ZN(new_n2718_));
  AOI21_X1  g2654(.A(new_n2718_), .B1(new_n2711_), .B2(new_n2713_), .ZN(new_n2719_));
  AOI21_X1  g2655(.A(new_n2707_), .B1(new_n2702_), .B2(new_n2703_), .ZN(new_n2720_));
  NOR2_X1   g2656(.A1(new_n2719_), .A2(new_n2720_), .ZN(new_n2721_));
  AOI21_X1  g2657(.A(new_n2675_), .B1(new_n2668_), .B2(new_n2674_), .ZN(new_n2722_));
  NAND2_X1  g2658(.A1(new_n2665_), .A2(new_n2673_), .ZN(new_n2723_));
  INV_X1    g2659(.A(new_n2723_), .ZN(new_n2724_));
  OR2_X1    g2660(.A1(new_n2722_), .A2(new_n2724_), .ZN(new_n2725_));
  AOI21_X1  g2661(.A(new_n2664_), .B1(new_n2654_), .B2(new_n2658_), .ZN(new_n2726_));
  NAND2_X1  g2662(.A1(G205gat), .A2(G477gat), .ZN(new_n2727_));
  NAND2_X1  g2663(.A1(new_n2633_), .A2(new_n2634_), .ZN(new_n2728_));
  NAND2_X1  g2664(.A1(new_n2728_), .A2(new_n2635_), .ZN(new_n2729_));
  NAND2_X1  g2665(.A1(new_n2729_), .A2(new_n2632_), .ZN(new_n2730_));
  NOR2_X1   g2666(.A1(new_n1805_), .A2(new_n544_), .ZN(new_n2731_));
  INV_X1    g2667(.A(new_n2731_), .ZN(new_n2732_));
  NAND2_X1  g2668(.A1(new_n2730_), .A2(new_n2732_), .ZN(new_n2733_));
  NAND2_X1  g2669(.A1(new_n2733_), .A2(new_n2732_), .ZN(new_n2734_));
  NAND2_X1  g2670(.A1(new_n2730_), .A2(new_n2731_), .ZN(new_n2735_));
  NAND2_X1  g2671(.A1(new_n2734_), .A2(new_n2735_), .ZN(new_n2736_));
  NOR2_X1   g2672(.A1(new_n1220_), .A2(new_n673_), .ZN(new_n2737_));
  AND2_X1   g2673(.A1(new_n2736_), .A2(new_n2737_), .ZN(new_n2738_));
  NOR2_X1   g2674(.A1(new_n2624_), .A2(new_n2638_), .ZN(new_n2739_));
  AOI21_X1  g2675(.A(new_n2739_), .B1(new_n2642_), .B2(new_n2643_), .ZN(new_n2740_));
  NOR2_X1   g2676(.A1(new_n2736_), .A2(new_n2737_), .ZN(new_n2741_));
  OR3_X1    g2677(.A1(new_n2738_), .A2(new_n2740_), .A3(new_n2741_), .ZN(new_n2742_));
  OAI21_X1  g2678(.A(new_n2740_), .B1(new_n2738_), .B2(new_n2741_), .ZN(new_n2743_));
  NAND2_X1  g2679(.A1(new_n2742_), .A2(new_n2743_), .ZN(new_n2744_));
  NOR2_X1   g2680(.A1(new_n1041_), .A2(new_n816_), .ZN(new_n2745_));
  NOR2_X1   g2681(.A1(new_n2744_), .A2(new_n2745_), .ZN(new_n2746_));
  INV_X1    g2682(.A(new_n2745_), .ZN(new_n2747_));
  AOI21_X1  g2683(.A(new_n2747_), .B1(new_n2742_), .B2(new_n2743_), .ZN(new_n2748_));
  NOR2_X1   g2684(.A1(new_n2746_), .A2(new_n2748_), .ZN(new_n2749_));
  NOR2_X1   g2685(.A1(new_n2644_), .A2(new_n2647_), .ZN(new_n2750_));
  AOI21_X1  g2686(.A(new_n2650_), .B1(new_n2648_), .B2(new_n2649_), .ZN(new_n2751_));
  OAI21_X1  g2687(.A(new_n2749_), .B1(new_n2750_), .B2(new_n2751_), .ZN(new_n2752_));
  NOR2_X1   g2688(.A1(new_n2751_), .A2(new_n2750_), .ZN(new_n2753_));
  OAI21_X1  g2689(.A(new_n2753_), .B1(new_n2748_), .B2(new_n2746_), .ZN(new_n2754_));
  AOI21_X1  g2690(.A(new_n2727_), .B1(new_n2752_), .B2(new_n2754_), .ZN(new_n2755_));
  AND3_X1   g2691(.A1(new_n2752_), .A2(new_n2754_), .A3(new_n2727_), .ZN(new_n2756_));
  OAI21_X1  g2692(.A(new_n2726_), .B1(new_n2755_), .B2(new_n2756_), .ZN(new_n2757_));
  OAI21_X1  g2693(.A(new_n2671_), .B1(new_n2659_), .B2(new_n2656_), .ZN(new_n2758_));
  NOR2_X1   g2694(.A1(new_n2756_), .A2(new_n2755_), .ZN(new_n2759_));
  NAND2_X1  g2695(.A1(new_n2758_), .A2(new_n2759_), .ZN(new_n2760_));
  NAND2_X1  g2696(.A1(G188gat), .A2(G494gat), .ZN(new_n2761_));
  AND3_X1   g2697(.A1(new_n2757_), .A2(new_n2760_), .A3(new_n2761_), .ZN(new_n2762_));
  AOI21_X1  g2698(.A(new_n2761_), .B1(new_n2757_), .B2(new_n2760_), .ZN(new_n2763_));
  NOR2_X1   g2699(.A1(new_n2762_), .A2(new_n2763_), .ZN(new_n2764_));
  NAND2_X1  g2700(.A1(new_n2725_), .A2(new_n2764_), .ZN(new_n2765_));
  NOR2_X1   g2701(.A1(new_n2722_), .A2(new_n2724_), .ZN(new_n2766_));
  OAI21_X1  g2702(.A(new_n2766_), .B1(new_n2762_), .B2(new_n2763_), .ZN(new_n2767_));
  NAND2_X1  g2703(.A1(new_n2765_), .A2(new_n2767_), .ZN(new_n2768_));
  AOI21_X1  g2704(.A(new_n2768_), .B1(G171gat), .B2(G511gat), .ZN(new_n2769_));
  NAND2_X1  g2705(.A1(G171gat), .A2(G511gat), .ZN(new_n2770_));
  AOI21_X1  g2706(.A(new_n2770_), .B1(new_n2765_), .B2(new_n2767_), .ZN(new_n2771_));
  NOR2_X1   g2707(.A1(new_n2769_), .A2(new_n2771_), .ZN(new_n2772_));
  NOR2_X1   g2708(.A1(new_n2691_), .A2(new_n2683_), .ZN(new_n2773_));
  NOR2_X1   g2709(.A1(new_n2773_), .A2(new_n2685_), .ZN(new_n2774_));
  OAI21_X1  g2710(.A(new_n2772_), .B1(new_n2688_), .B2(new_n2774_), .ZN(new_n2775_));
  NOR2_X1   g2711(.A1(new_n2774_), .A2(new_n2688_), .ZN(new_n2776_));
  OAI21_X1  g2712(.A(new_n2776_), .B1(new_n2771_), .B2(new_n2769_), .ZN(new_n2777_));
  NAND2_X1  g2713(.A1(new_n2775_), .A2(new_n2777_), .ZN(new_n2778_));
  NOR2_X1   g2714(.A1(new_n889_), .A2(new_n1741_), .ZN(new_n2779_));
  XNOR2_X1  g2715(.A(new_n2778_), .B(new_n2779_), .ZN(new_n2780_));
  AOI21_X1  g2716(.A(new_n2701_), .B1(new_n2698_), .B2(new_n2699_), .ZN(new_n2781_));
  AOI21_X1  g2717(.A(new_n2697_), .B1(new_n2692_), .B2(new_n2689_), .ZN(new_n2782_));
  NOR2_X1   g2718(.A1(new_n2781_), .A2(new_n2782_), .ZN(new_n2783_));
  INV_X1    g2719(.A(new_n2783_), .ZN(new_n2784_));
  XNOR2_X1  g2720(.A(new_n2780_), .B(new_n2784_), .ZN(new_n2785_));
  XNOR2_X1  g2721(.A(new_n2721_), .B(new_n2785_), .ZN(G6230gat));
  NOR2_X1   g2722(.A1(new_n873_), .A2(new_n1155_), .ZN(new_n2787_));
  INV_X1    g2723(.A(new_n2787_), .ZN(new_n2788_));
  INV_X1    g2724(.A(new_n2736_), .ZN(new_n2789_));
  OAI21_X1  g2725(.A(new_n2733_), .B1(new_n2789_), .B2(new_n2737_), .ZN(new_n2790_));
  NOR2_X1   g2726(.A1(new_n1805_), .A2(new_n673_), .ZN(new_n2791_));
  INV_X1    g2727(.A(new_n2791_), .ZN(new_n2792_));
  NAND2_X1  g2728(.A1(new_n2790_), .A2(new_n2792_), .ZN(new_n2793_));
  NAND2_X1  g2729(.A1(new_n2793_), .A2(new_n2792_), .ZN(new_n2794_));
  NAND2_X1  g2730(.A1(new_n2790_), .A2(new_n2791_), .ZN(new_n2795_));
  NAND2_X1  g2731(.A1(new_n2794_), .A2(new_n2795_), .ZN(new_n2796_));
  AOI21_X1  g2732(.A(new_n2796_), .B1(G239gat), .B2(G460gat), .ZN(new_n2797_));
  NAND2_X1  g2733(.A1(G239gat), .A2(G460gat), .ZN(new_n2798_));
  AOI21_X1  g2734(.A(new_n2798_), .B1(new_n2794_), .B2(new_n2795_), .ZN(new_n2799_));
  NOR2_X1   g2735(.A1(new_n2797_), .A2(new_n2799_), .ZN(new_n2800_));
  NOR2_X1   g2736(.A1(new_n2738_), .A2(new_n2741_), .ZN(new_n2801_));
  NOR2_X1   g2737(.A1(new_n2801_), .A2(new_n2740_), .ZN(new_n2802_));
  AOI21_X1  g2738(.A(new_n2802_), .B1(new_n2744_), .B2(new_n2747_), .ZN(new_n2803_));
  INV_X1    g2739(.A(new_n2803_), .ZN(new_n2804_));
  NOR2_X1   g2740(.A1(new_n2800_), .A2(new_n2804_), .ZN(new_n2805_));
  INV_X1    g2741(.A(new_n2805_), .ZN(new_n2806_));
  NAND2_X1  g2742(.A1(new_n2800_), .A2(new_n2804_), .ZN(new_n2807_));
  NOR2_X1   g2743(.A1(new_n1041_), .A2(new_n980_), .ZN(new_n2808_));
  INV_X1    g2744(.A(new_n2808_), .ZN(new_n2809_));
  AND3_X1   g2745(.A1(new_n2806_), .A2(new_n2807_), .A3(new_n2809_), .ZN(new_n2810_));
  AOI21_X1  g2746(.A(new_n2809_), .B1(new_n2806_), .B2(new_n2807_), .ZN(new_n2811_));
  NOR2_X1   g2747(.A1(new_n2810_), .A2(new_n2811_), .ZN(new_n2812_));
  NOR2_X1   g2748(.A1(new_n2749_), .A2(new_n2753_), .ZN(new_n2813_));
  NAND2_X1  g2749(.A1(new_n2752_), .A2(new_n2754_), .ZN(new_n2814_));
  AOI21_X1  g2750(.A(new_n2813_), .B1(new_n2814_), .B2(new_n2727_), .ZN(new_n2815_));
  INV_X1    g2751(.A(new_n2815_), .ZN(new_n2816_));
  NOR2_X1   g2752(.A1(new_n2812_), .A2(new_n2816_), .ZN(new_n2817_));
  INV_X1    g2753(.A(new_n2817_), .ZN(new_n2818_));
  NAND2_X1  g2754(.A1(new_n2812_), .A2(new_n2816_), .ZN(new_n2819_));
  AOI21_X1  g2755(.A(new_n2788_), .B1(new_n2818_), .B2(new_n2819_), .ZN(new_n2820_));
  INV_X1    g2756(.A(new_n2819_), .ZN(new_n2821_));
  NOR3_X1   g2757(.A1(new_n2821_), .A2(new_n2817_), .A3(new_n2787_), .ZN(new_n2822_));
  NOR2_X1   g2758(.A1(new_n2820_), .A2(new_n2822_), .ZN(new_n2823_));
  NOR2_X1   g2759(.A1(new_n2726_), .A2(new_n2759_), .ZN(new_n2824_));
  AOI22_X1  g2760(.A1(new_n2757_), .A2(new_n2760_), .B1(G188gat), .B2(G494gat), .ZN(new_n2825_));
  OAI21_X1  g2761(.A(new_n2823_), .B1(new_n2824_), .B2(new_n2825_), .ZN(new_n2826_));
  NOR2_X1   g2762(.A1(new_n2825_), .A2(new_n2824_), .ZN(new_n2827_));
  OAI21_X1  g2763(.A(new_n2827_), .B1(new_n2822_), .B2(new_n2820_), .ZN(new_n2828_));
  NAND2_X1  g2764(.A1(G188gat), .A2(G511gat), .ZN(new_n2829_));
  AND3_X1   g2765(.A1(new_n2826_), .A2(new_n2828_), .A3(new_n2829_), .ZN(new_n2830_));
  AOI21_X1  g2766(.A(new_n2829_), .B1(new_n2826_), .B2(new_n2828_), .ZN(new_n2831_));
  NOR2_X1   g2767(.A1(new_n2830_), .A2(new_n2831_), .ZN(new_n2832_));
  AND2_X1   g2768(.A1(new_n2768_), .A2(new_n2770_), .ZN(new_n2833_));
  NOR2_X1   g2769(.A1(new_n2764_), .A2(new_n2766_), .ZN(new_n2834_));
  OAI21_X1  g2770(.A(new_n2832_), .B1(new_n2833_), .B2(new_n2834_), .ZN(new_n2835_));
  NOR2_X1   g2771(.A1(new_n2833_), .A2(new_n2834_), .ZN(new_n2836_));
  OAI21_X1  g2772(.A(new_n2836_), .B1(new_n2830_), .B2(new_n2831_), .ZN(new_n2837_));
  NAND2_X1  g2773(.A1(new_n2835_), .A2(new_n2837_), .ZN(new_n2838_));
  NAND2_X1  g2774(.A1(G171gat), .A2(G528gat), .ZN(new_n2839_));
  XNOR2_X1  g2775(.A(new_n2838_), .B(new_n2839_), .ZN(new_n2840_));
  OAI21_X1  g2776(.A(new_n2778_), .B1(new_n889_), .B2(new_n1741_), .ZN(new_n2841_));
  OAI21_X1  g2777(.A(new_n2841_), .B1(new_n2772_), .B2(new_n2776_), .ZN(new_n2842_));
  INV_X1    g2778(.A(new_n2842_), .ZN(new_n2843_));
  XNOR2_X1  g2779(.A(new_n2840_), .B(new_n2843_), .ZN(new_n2844_));
  INV_X1    g2780(.A(new_n2844_), .ZN(new_n2845_));
  XNOR2_X1  g2781(.A(new_n2780_), .B(new_n2783_), .ZN(new_n2846_));
  OAI21_X1  g2782(.A(new_n2846_), .B1(new_n2719_), .B2(new_n2720_), .ZN(new_n2847_));
  NAND2_X1  g2783(.A1(new_n2780_), .A2(new_n2784_), .ZN(new_n2848_));
  AOI21_X1  g2784(.A(new_n2845_), .B1(new_n2847_), .B2(new_n2848_), .ZN(new_n2849_));
  INV_X1    g2785(.A(new_n2720_), .ZN(new_n2850_));
  AOI21_X1  g2786(.A(new_n2785_), .B1(new_n2716_), .B2(new_n2850_), .ZN(new_n2851_));
  INV_X1    g2787(.A(new_n2848_), .ZN(new_n2852_));
  OAI21_X1  g2788(.A(new_n2845_), .B1(new_n2851_), .B2(new_n2852_), .ZN(new_n2853_));
  AOI21_X1  g2789(.A(new_n2849_), .B1(new_n2853_), .B2(new_n2845_), .ZN(G6240gat));
  AOI21_X1  g2790(.A(new_n2844_), .B1(new_n2847_), .B2(new_n2848_), .ZN(new_n2855_));
  NOR2_X1   g2791(.A1(new_n2840_), .A2(new_n2843_), .ZN(new_n2856_));
  NOR2_X1   g2792(.A1(new_n2855_), .A2(new_n2856_), .ZN(new_n2857_));
  AOI21_X1  g2793(.A(new_n2808_), .B1(new_n2806_), .B2(new_n2807_), .ZN(new_n2858_));
  NOR2_X1   g2794(.A1(new_n2800_), .A2(new_n2803_), .ZN(new_n2859_));
  NOR2_X1   g2795(.A1(new_n2858_), .A2(new_n2859_), .ZN(new_n2860_));
  INV_X1    g2796(.A(new_n2860_), .ZN(new_n2861_));
  NAND2_X1  g2797(.A1(new_n2796_), .A2(new_n2798_), .ZN(new_n2862_));
  NAND2_X1  g2798(.A1(new_n2862_), .A2(new_n2793_), .ZN(new_n2863_));
  NOR2_X1   g2799(.A1(new_n1805_), .A2(new_n816_), .ZN(new_n2864_));
  XNOR2_X1  g2800(.A(new_n2863_), .B(new_n2864_), .ZN(new_n2865_));
  NOR2_X1   g2801(.A1(new_n1220_), .A2(new_n980_), .ZN(new_n2866_));
  INV_X1    g2802(.A(new_n2866_), .ZN(new_n2867_));
  XNOR2_X1  g2803(.A(new_n2865_), .B(new_n2867_), .ZN(new_n2868_));
  OR2_X1    g2804(.A1(new_n2861_), .A2(new_n2868_), .ZN(new_n2869_));
  NAND2_X1  g2805(.A1(new_n2861_), .A2(new_n2868_), .ZN(new_n2870_));
  NAND2_X1  g2806(.A1(new_n2869_), .A2(new_n2870_), .ZN(new_n2871_));
  AOI21_X1  g2807(.A(new_n2871_), .B1(G222gat), .B2(G494gat), .ZN(new_n2872_));
  NAND2_X1  g2808(.A1(G222gat), .A2(G494gat), .ZN(new_n2873_));
  AOI21_X1  g2809(.A(new_n2873_), .B1(new_n2869_), .B2(new_n2870_), .ZN(new_n2874_));
  NOR2_X1   g2810(.A1(new_n2872_), .A2(new_n2874_), .ZN(new_n2875_));
  AOI21_X1  g2811(.A(new_n2787_), .B1(new_n2818_), .B2(new_n2819_), .ZN(new_n2876_));
  NOR2_X1   g2812(.A1(new_n2812_), .A2(new_n2815_), .ZN(new_n2877_));
  NOR2_X1   g2813(.A1(new_n2876_), .A2(new_n2877_), .ZN(new_n2878_));
  XNOR2_X1  g2814(.A(new_n2875_), .B(new_n2878_), .ZN(new_n2879_));
  NOR2_X1   g2815(.A1(new_n873_), .A2(new_n1345_), .ZN(new_n2880_));
  XOR2_X1   g2816(.A(new_n2879_), .B(new_n2880_), .Z(new_n2881_));
  AOI22_X1  g2817(.A1(new_n2826_), .A2(new_n2828_), .B1(G188gat), .B2(G511gat), .ZN(new_n2882_));
  NOR2_X1   g2818(.A1(new_n2823_), .A2(new_n2827_), .ZN(new_n2883_));
  NOR2_X1   g2819(.A1(new_n2882_), .A2(new_n2883_), .ZN(new_n2884_));
  NAND2_X1  g2820(.A1(new_n2881_), .A2(new_n2884_), .ZN(new_n2885_));
  XNOR2_X1  g2821(.A(new_n2879_), .B(new_n2880_), .ZN(new_n2886_));
  OAI21_X1  g2822(.A(new_n2886_), .B1(new_n2883_), .B2(new_n2882_), .ZN(new_n2887_));
  NAND2_X1  g2823(.A1(G188gat), .A2(G528gat), .ZN(new_n2888_));
  AND3_X1   g2824(.A1(new_n2885_), .A2(new_n2887_), .A3(new_n2888_), .ZN(new_n2889_));
  AOI21_X1  g2825(.A(new_n2888_), .B1(new_n2885_), .B2(new_n2887_), .ZN(new_n2890_));
  NOR2_X1   g2826(.A1(new_n2889_), .A2(new_n2890_), .ZN(new_n2891_));
  NOR2_X1   g2827(.A1(new_n2832_), .A2(new_n2836_), .ZN(new_n2892_));
  AOI21_X1  g2828(.A(new_n2892_), .B1(new_n2838_), .B2(new_n2839_), .ZN(new_n2893_));
  XNOR2_X1  g2829(.A(new_n2891_), .B(new_n2893_), .ZN(new_n2894_));
  XNOR2_X1  g2830(.A(new_n2857_), .B(new_n2894_), .ZN(G6250gat));
  NOR2_X1   g2831(.A1(new_n2879_), .A2(new_n2880_), .ZN(new_n2896_));
  NOR2_X1   g2832(.A1(new_n2875_), .A2(new_n2878_), .ZN(new_n2897_));
  NOR2_X1   g2833(.A1(new_n2896_), .A2(new_n2897_), .ZN(new_n2898_));
  INV_X1    g2834(.A(new_n2898_), .ZN(new_n2899_));
  NAND2_X1  g2835(.A1(new_n2871_), .A2(new_n2873_), .ZN(new_n2900_));
  OAI21_X1  g2836(.A(new_n2900_), .B1(new_n2868_), .B2(new_n2860_), .ZN(new_n2901_));
  NAND2_X1  g2837(.A1(new_n2865_), .A2(new_n2867_), .ZN(new_n2902_));
  OAI21_X1  g2838(.A(new_n2863_), .B1(new_n1805_), .B2(new_n816_), .ZN(new_n2903_));
  NAND2_X1  g2839(.A1(new_n2902_), .A2(new_n2903_), .ZN(new_n2904_));
  NAND2_X1  g2840(.A1(G256gat), .A2(G477gat), .ZN(new_n2905_));
  XNOR2_X1  g2841(.A(new_n2904_), .B(new_n2905_), .ZN(new_n2906_));
  NOR2_X1   g2842(.A1(new_n1220_), .A2(new_n1155_), .ZN(new_n2907_));
  XNOR2_X1  g2843(.A(new_n2906_), .B(new_n2907_), .ZN(new_n2908_));
  INV_X1    g2844(.A(new_n2908_), .ZN(new_n2909_));
  XNOR2_X1  g2845(.A(new_n2901_), .B(new_n2909_), .ZN(new_n2910_));
  NOR2_X1   g2846(.A1(new_n1041_), .A2(new_n1345_), .ZN(new_n2911_));
  XNOR2_X1  g2847(.A(new_n2910_), .B(new_n2911_), .ZN(new_n2912_));
  OR2_X1    g2848(.A1(new_n2899_), .A2(new_n2912_), .ZN(new_n2913_));
  NAND2_X1  g2849(.A1(new_n2899_), .A2(new_n2912_), .ZN(new_n2914_));
  NAND2_X1  g2850(.A1(G205gat), .A2(G528gat), .ZN(new_n2915_));
  AND3_X1   g2851(.A1(new_n2913_), .A2(new_n2914_), .A3(new_n2915_), .ZN(new_n2916_));
  AOI21_X1  g2852(.A(new_n2915_), .B1(new_n2913_), .B2(new_n2914_), .ZN(new_n2917_));
  NOR2_X1   g2853(.A1(new_n2916_), .A2(new_n2917_), .ZN(new_n2918_));
  NAND2_X1  g2854(.A1(new_n2885_), .A2(new_n2887_), .ZN(new_n2919_));
  NAND2_X1  g2855(.A1(new_n2919_), .A2(new_n2888_), .ZN(new_n2920_));
  OAI21_X1  g2856(.A(new_n2920_), .B1(new_n2886_), .B2(new_n2884_), .ZN(new_n2921_));
  XOR2_X1   g2857(.A(new_n2918_), .B(new_n2921_), .Z(new_n2922_));
  INV_X1    g2858(.A(new_n2922_), .ZN(new_n2923_));
  XOR2_X1   g2859(.A(new_n2891_), .B(new_n2893_), .Z(new_n2924_));
  OAI21_X1  g2860(.A(new_n2924_), .B1(new_n2855_), .B2(new_n2856_), .ZN(new_n2925_));
  NOR2_X1   g2861(.A1(new_n2891_), .A2(new_n2893_), .ZN(new_n2926_));
  INV_X1    g2862(.A(new_n2926_), .ZN(new_n2927_));
  AOI21_X1  g2863(.A(new_n2923_), .B1(new_n2925_), .B2(new_n2927_), .ZN(new_n2928_));
  INV_X1    g2864(.A(new_n2856_), .ZN(new_n2929_));
  AOI21_X1  g2865(.A(new_n2894_), .B1(new_n2853_), .B2(new_n2929_), .ZN(new_n2930_));
  OAI21_X1  g2866(.A(new_n2923_), .B1(new_n2930_), .B2(new_n2926_), .ZN(new_n2931_));
  AOI21_X1  g2867(.A(new_n2928_), .B1(new_n2931_), .B2(new_n2923_), .ZN(G6260gat));
  AOI21_X1  g2868(.A(new_n2922_), .B1(new_n2925_), .B2(new_n2927_), .ZN(new_n2933_));
  OAI21_X1  g2869(.A(new_n2921_), .B1(new_n2917_), .B2(new_n2916_), .ZN(new_n2934_));
  INV_X1    g2870(.A(new_n2934_), .ZN(new_n2935_));
  NOR2_X1   g2871(.A1(new_n2933_), .A2(new_n2935_), .ZN(new_n2936_));
  NAND2_X1  g2872(.A1(new_n2913_), .A2(new_n2914_), .ZN(new_n2937_));
  NAND2_X1  g2873(.A1(new_n2937_), .A2(new_n2915_), .ZN(new_n2938_));
  OAI21_X1  g2874(.A(new_n2938_), .B1(new_n2912_), .B2(new_n2898_), .ZN(new_n2939_));
  NAND2_X1  g2875(.A1(new_n2901_), .A2(new_n2909_), .ZN(new_n2940_));
  OAI21_X1  g2876(.A(new_n2940_), .B1(new_n2910_), .B2(new_n2911_), .ZN(new_n2941_));
  NAND2_X1  g2877(.A1(new_n2904_), .A2(new_n2905_), .ZN(new_n2942_));
  OAI21_X1  g2878(.A(new_n2942_), .B1(new_n2906_), .B2(new_n2907_), .ZN(new_n2943_));
  NOR2_X1   g2879(.A1(new_n1805_), .A2(new_n1155_), .ZN(new_n2944_));
  XNOR2_X1  g2880(.A(new_n2943_), .B(new_n2944_), .ZN(new_n2945_));
  NOR2_X1   g2881(.A1(new_n1220_), .A2(new_n1345_), .ZN(new_n2946_));
  INV_X1    g2882(.A(new_n2946_), .ZN(new_n2947_));
  XNOR2_X1  g2883(.A(new_n2945_), .B(new_n2947_), .ZN(new_n2948_));
  XNOR2_X1  g2884(.A(new_n2941_), .B(new_n2948_), .ZN(new_n2949_));
  NOR2_X1   g2885(.A1(new_n1041_), .A2(new_n1741_), .ZN(new_n2950_));
  XNOR2_X1  g2886(.A(new_n2949_), .B(new_n2950_), .ZN(new_n2951_));
  XNOR2_X1  g2887(.A(new_n2939_), .B(new_n2951_), .ZN(new_n2952_));
  XNOR2_X1  g2888(.A(new_n2936_), .B(new_n2952_), .ZN(G6270gat));
  INV_X1    g2889(.A(new_n2950_), .ZN(new_n2954_));
  NAND2_X1  g2890(.A1(new_n2949_), .A2(new_n2954_), .ZN(new_n2955_));
  INV_X1    g2891(.A(new_n2948_), .ZN(new_n2956_));
  NAND2_X1  g2892(.A1(new_n2941_), .A2(new_n2956_), .ZN(new_n2957_));
  NAND2_X1  g2893(.A1(new_n2955_), .A2(new_n2957_), .ZN(new_n2958_));
  NAND2_X1  g2894(.A1(new_n2945_), .A2(new_n2947_), .ZN(new_n2959_));
  OAI21_X1  g2895(.A(new_n2943_), .B1(new_n1805_), .B2(new_n1155_), .ZN(new_n2960_));
  NAND2_X1  g2896(.A1(new_n2959_), .A2(new_n2960_), .ZN(new_n2961_));
  NAND2_X1  g2897(.A1(G256gat), .A2(G511gat), .ZN(new_n2962_));
  XNOR2_X1  g2898(.A(new_n2961_), .B(new_n2962_), .ZN(new_n2963_));
  NOR2_X1   g2899(.A1(new_n1220_), .A2(new_n1741_), .ZN(new_n2964_));
  XNOR2_X1  g2900(.A(new_n2963_), .B(new_n2964_), .ZN(new_n2965_));
  XOR2_X1   g2901(.A(new_n2958_), .B(new_n2965_), .Z(new_n2966_));
  INV_X1    g2902(.A(new_n2966_), .ZN(new_n2967_));
  INV_X1    g2903(.A(new_n2952_), .ZN(new_n2968_));
  OAI21_X1  g2904(.A(new_n2968_), .B1(new_n2933_), .B2(new_n2935_), .ZN(new_n2969_));
  NAND2_X1  g2905(.A1(new_n2939_), .A2(new_n2951_), .ZN(new_n2970_));
  AOI21_X1  g2906(.A(new_n2967_), .B1(new_n2969_), .B2(new_n2970_), .ZN(new_n2971_));
  AOI21_X1  g2907(.A(new_n2952_), .B1(new_n2931_), .B2(new_n2934_), .ZN(new_n2972_));
  INV_X1    g2908(.A(new_n2970_), .ZN(new_n2973_));
  OAI21_X1  g2909(.A(new_n2967_), .B1(new_n2972_), .B2(new_n2973_), .ZN(new_n2974_));
  AOI21_X1  g2910(.A(new_n2971_), .B1(new_n2974_), .B2(new_n2967_), .ZN(G6280gat));
  NOR2_X1   g2911(.A1(new_n1805_), .A2(new_n1741_), .ZN(new_n2976_));
  OR2_X1    g2912(.A1(new_n2963_), .A2(new_n2964_), .ZN(new_n2977_));
  NAND2_X1  g2913(.A1(new_n2961_), .A2(new_n2962_), .ZN(new_n2978_));
  AOI21_X1  g2914(.A(new_n2976_), .B1(new_n2977_), .B2(new_n2978_), .ZN(new_n2979_));
  INV_X1    g2915(.A(new_n2958_), .ZN(new_n2980_));
  NOR2_X1   g2916(.A1(new_n2980_), .A2(new_n2965_), .ZN(new_n2981_));
  INV_X1    g2917(.A(new_n2981_), .ZN(new_n2982_));
  NAND2_X1  g2918(.A1(new_n2974_), .A2(new_n2982_), .ZN(new_n2983_));
  NAND2_X1  g2919(.A1(new_n2977_), .A2(new_n2978_), .ZN(new_n2984_));
  XOR2_X1   g2920(.A(new_n2984_), .B(new_n2976_), .Z(new_n2985_));
  INV_X1    g2921(.A(new_n2985_), .ZN(new_n2986_));
  AOI21_X1  g2922(.A(new_n2979_), .B1(new_n2983_), .B2(new_n2986_), .ZN(G6287gat));
  AOI21_X1  g2923(.A(new_n2986_), .B1(new_n2974_), .B2(new_n2982_), .ZN(new_n2988_));
  AOI21_X1  g2924(.A(new_n2966_), .B1(new_n2969_), .B2(new_n2970_), .ZN(new_n2989_));
  NOR3_X1   g2925(.A1(new_n2989_), .A2(new_n2981_), .A3(new_n2985_), .ZN(new_n2990_));
  NOR2_X1   g2926(.A1(new_n2988_), .A2(new_n2990_), .ZN(G6288gat));
endmodule


