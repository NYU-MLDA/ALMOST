//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT82), .ZN(new_n203_));
  INV_X1    g002(.A(G71gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G99gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  AOI22_X1  g010(.A1(new_n207_), .A2(new_n208_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT24), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT81), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n216_), .A2(new_n219_), .A3(KEYINPUT81), .A4(new_n220_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n212_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(G169gat), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n219_), .B(new_n220_), .C1(G183gat), .C2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n206_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n231_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G15gat), .B(G43gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT83), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT30), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT31), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n236_), .A2(new_n240_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G141gat), .ZN(new_n245_));
  INV_X1    g044(.A(G148gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G141gat), .A2(G148gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G155gat), .B(G162gat), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n252_), .B2(KEYINPUT1), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT2), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n247_), .A2(KEYINPUT3), .B1(new_n254_), .B2(new_n248_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT85), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT85), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n258_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT84), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G141gat), .A2(G148gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NOR4_X1   g063(.A1(KEYINPUT84), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n255_), .B(new_n260_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT86), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT84), .B1(new_n247_), .B2(KEYINPUT3), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n262_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n271_), .A2(KEYINPUT86), .A3(new_n260_), .A4(new_n255_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n252_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n253_), .B1(new_n273_), .B2(KEYINPUT87), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT87), .ZN(new_n275_));
  AOI211_X1 g074(.A(new_n275_), .B(new_n252_), .C1(new_n268_), .C2(new_n272_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n235_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n266_), .A2(new_n267_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n248_), .A2(new_n254_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT86), .B1(new_n282_), .B2(new_n260_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n251_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n275_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n273_), .A2(KEYINPUT87), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n285_), .A2(new_n234_), .A3(new_n286_), .A4(new_n253_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G225gat), .A2(G233gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n277_), .A2(new_n287_), .A3(KEYINPUT4), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n291_), .B(new_n235_), .C1(new_n274_), .C2(new_n276_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n288_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n289_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G29gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G85gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT0), .B(G57gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n289_), .B(new_n299_), .C1(new_n290_), .C2(new_n294_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n244_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G78gat), .B(G106gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT89), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT29), .B1(new_n274_), .B2(new_n276_), .ZN(new_n309_));
  INV_X1    g108(.A(G228gat), .ZN(new_n310_));
  INV_X1    g109(.A(G233gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(G197gat), .A2(G204gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G197gat), .A2(G204gat), .ZN(new_n317_));
  AND2_X1   g116(.A1(KEYINPUT88), .A2(KEYINPUT21), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n317_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT21), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n314_), .A2(new_n316_), .A3(new_n317_), .A4(new_n318_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n309_), .A2(new_n313_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n313_), .B1(new_n309_), .B2(new_n326_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n308_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n329_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n327_), .A3(new_n307_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n332_), .A3(KEYINPUT90), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n285_), .A2(new_n286_), .A3(new_n253_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT28), .B1(new_n334_), .B2(KEYINPUT29), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n274_), .A2(KEYINPUT29), .A3(new_n276_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT28), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G22gat), .B(G50gat), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n335_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT90), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n331_), .A2(new_n327_), .A3(new_n343_), .A4(new_n307_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n333_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT91), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n332_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n340_), .A2(new_n341_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n331_), .A2(new_n327_), .A3(KEYINPUT91), .A4(new_n307_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n306_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .A4(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n345_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT100), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  INV_X1    g153(.A(new_n221_), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n212_), .A2(new_n355_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n357_), .B2(new_n326_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n225_), .A2(new_n325_), .A3(new_n229_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n362_), .B(KEYINPUT92), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n230_), .A2(new_n326_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT93), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n325_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT93), .ZN(new_n370_));
  INV_X1    g169(.A(new_n362_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n354_), .B1(new_n356_), .B2(new_n325_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n365_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT95), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n378_), .B(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n374_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n378_), .B(new_n379_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(new_n365_), .A3(new_n373_), .ZN(new_n384_));
  AOI211_X1 g183(.A(new_n353_), .B(KEYINPUT27), .C1(new_n382_), .C2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n384_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT100), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n370_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n372_), .B1(new_n369_), .B2(KEYINPUT93), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OAI22_X1  g190(.A1(new_n391_), .A2(new_n371_), .B1(new_n364_), .B2(new_n360_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n383_), .A2(KEYINPUT98), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT98), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n381_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT99), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n384_), .A2(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n383_), .A2(new_n365_), .A3(new_n373_), .A4(KEYINPUT99), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n396_), .A2(new_n398_), .A3(KEYINPUT27), .A4(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n385_), .B1(new_n388_), .B2(new_n400_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n305_), .A2(new_n352_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n292_), .A2(new_n288_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n277_), .A2(new_n287_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(KEYINPUT4), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n277_), .A2(new_n287_), .A3(new_n293_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n300_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT96), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n277_), .A2(new_n287_), .A3(KEYINPUT4), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(new_n288_), .A3(new_n292_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT96), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n300_), .A4(new_n406_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n386_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT33), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n302_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n409_), .A2(new_n293_), .A3(new_n292_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n417_), .A2(KEYINPUT33), .A3(new_n289_), .A4(new_n299_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n413_), .A2(new_n414_), .A3(new_n416_), .A4(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n383_), .A2(KEYINPUT32), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(new_n374_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n392_), .B2(new_n420_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n302_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n299_), .B1(new_n417_), .B2(new_n289_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT97), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT97), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n303_), .A2(new_n427_), .A3(new_n422_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n419_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n352_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n401_), .B1(new_n345_), .B2(new_n351_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n304_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n402_), .B1(new_n434_), .B2(new_n243_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G29gat), .B(G36gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT76), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G43gat), .B(G50gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G15gat), .B(G22gat), .ZN(new_n441_));
  INV_X1    g240(.A(G1gat), .ZN(new_n442_));
  INV_X1    g241(.A(G8gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT14), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G8gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n440_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n439_), .B(KEYINPUT15), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n447_), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n439_), .B(new_n447_), .Z(new_n453_));
  INV_X1    g252(.A(new_n449_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n450_), .A2(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G113gat), .B(G141gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(G169gat), .B(G197gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n458_), .A2(KEYINPUT80), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n455_), .B(new_n459_), .Z(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n435_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G57gat), .B(G64gat), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n463_), .A2(KEYINPUT11), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(KEYINPUT11), .ZN(new_n465_));
  XOR2_X1   g264(.A(G71gat), .B(G78gat), .Z(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n465_), .A2(new_n466_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G231gat), .A2(G233gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n469_), .B(new_n470_), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT79), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(new_n447_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G127gat), .B(G155gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT16), .ZN(new_n475_));
  XOR2_X1   g274(.A(G183gat), .B(G211gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n473_), .A2(KEYINPUT17), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n477_), .B(KEYINPUT17), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n479_), .B1(new_n473_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G190gat), .B(G218gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G134gat), .B(G162gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n485_), .A2(KEYINPUT36), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT6), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G106gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT10), .B(G99gat), .Z(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT9), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT65), .B(G92gat), .ZN(new_n496_));
  INV_X1    g295(.A(G85gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  AND2_X1   g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(KEYINPUT9), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n494_), .B1(new_n500_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT67), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT8), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n502_), .A2(new_n501_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT7), .ZN(new_n509_));
  INV_X1    g308(.A(G99gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n492_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n507_), .B(new_n508_), .C1(new_n491_), .C2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT68), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n491_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT69), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n511_), .A2(new_n517_), .A3(new_n512_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(KEYINPUT69), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n488_), .A2(new_n490_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT68), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .A4(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(KEYINPUT70), .A3(new_n508_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT8), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT70), .B1(new_n522_), .B2(new_n508_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n514_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n506_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT77), .B1(new_n527_), .B2(new_n440_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT77), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n506_), .A2(new_n526_), .A3(new_n529_), .A4(new_n439_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n451_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G232gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT75), .B(KEYINPUT35), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n528_), .A2(new_n530_), .A3(new_n531_), .A4(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n534_), .A2(new_n535_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(KEYINPUT78), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(KEYINPUT78), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n541_), .B1(new_n537_), .B2(new_n542_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n486_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n545_), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n485_), .B(KEYINPUT36), .Z(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n543_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT37), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n549_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n482_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G120gat), .B(G148gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT73), .Z(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT64), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n506_), .A2(new_n526_), .A3(new_n469_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n469_), .B1(new_n506_), .B2(new_n526_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n564_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT71), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT71), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n570_), .B(new_n564_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n567_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(KEYINPUT12), .A3(new_n565_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n567_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n564_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n561_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n566_), .A2(new_n567_), .A3(new_n575_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n576_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n563_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n559_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n571_), .A4(new_n569_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n578_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n554_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n462_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n442_), .A3(new_n303_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT38), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n587_), .A2(new_n461_), .A3(new_n482_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT101), .ZN(new_n596_));
  INV_X1    g395(.A(new_n550_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n596_), .B1(new_n435_), .B2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n352_), .A2(new_n401_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(new_n304_), .A3(new_n244_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n429_), .A2(new_n430_), .B1(new_n432_), .B2(new_n304_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n600_), .B1(new_n601_), .B2(new_n244_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(KEYINPUT101), .A3(new_n550_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n595_), .B1(new_n598_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G1gat), .B1(new_n605_), .B2(new_n304_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n593_), .A2(new_n606_), .ZN(G1324gat));
  AND3_X1   g406(.A1(new_n602_), .A2(KEYINPUT101), .A3(new_n550_), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT101), .B1(new_n602_), .B2(new_n550_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n401_), .B(new_n594_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT102), .ZN(new_n611_));
  OAI21_X1  g410(.A(G8gat), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT102), .B1(new_n604_), .B2(new_n401_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT39), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n604_), .A2(KEYINPUT102), .A3(new_n401_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n610_), .A2(new_n611_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .A4(G8gat), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n591_), .A2(new_n443_), .A3(new_n401_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(KEYINPUT40), .A3(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1325gat));
  OAI21_X1  g424(.A(G15gat), .B1(new_n605_), .B2(new_n243_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n627_), .ZN(new_n629_));
  OR3_X1    g428(.A1(new_n590_), .A2(G15gat), .A3(new_n243_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(G1326gat));
  OR3_X1    g430(.A1(new_n590_), .A2(G22gat), .A3(new_n430_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G22gat), .B1(new_n605_), .B2(new_n430_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(KEYINPUT42), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(KEYINPUT42), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n632_), .B1(new_n634_), .B2(new_n635_), .ZN(G1327gat));
  NAND2_X1  g435(.A1(new_n551_), .A2(new_n553_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT43), .B1(new_n435_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  INV_X1    g438(.A(new_n637_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n602_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n460_), .B(new_n482_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT104), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT44), .B1(new_n642_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n647_), .B(new_n644_), .C1(new_n638_), .C2(new_n641_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n646_), .A2(new_n648_), .A3(new_n304_), .ZN(new_n649_));
  INV_X1    g448(.A(G29gat), .ZN(new_n650_));
  INV_X1    g449(.A(new_n482_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n550_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n462_), .A2(new_n588_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n303_), .A2(new_n650_), .ZN(new_n654_));
  OAI22_X1  g453(.A1(new_n649_), .A2(new_n650_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(new_n401_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n653_), .A2(G36gat), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT45), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n646_), .A2(new_n648_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(new_n401_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n602_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n639_), .B1(new_n602_), .B2(new_n640_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n645_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n647_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n645_), .B(KEYINPUT44), .C1(new_n665_), .C2(new_n666_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n668_), .A2(new_n662_), .A3(new_n401_), .A4(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G36gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n661_), .B1(new_n664_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT46), .B(new_n661_), .C1(new_n664_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1329gat));
  NAND3_X1  g475(.A1(new_n663_), .A2(G43gat), .A3(new_n244_), .ZN(new_n677_));
  INV_X1    g476(.A(G43gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n678_), .B1(new_n653_), .B2(new_n243_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g480(.A1(new_n663_), .A2(KEYINPUT107), .A3(new_n352_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G50gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT107), .B1(new_n663_), .B2(new_n352_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n430_), .A2(G50gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT108), .ZN(new_n686_));
  OAI22_X1  g485(.A1(new_n683_), .A2(new_n684_), .B1(new_n653_), .B2(new_n686_), .ZN(G1331gat));
  NAND2_X1  g486(.A1(new_n598_), .A2(new_n603_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n588_), .A2(new_n460_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n651_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT109), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n688_), .A2(new_n692_), .A3(new_n651_), .A4(new_n689_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n303_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G57gat), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n689_), .A2(new_n602_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n554_), .ZN(new_n697_));
  OR3_X1    g496(.A1(new_n697_), .A2(G57gat), .A3(new_n304_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n695_), .A2(KEYINPUT110), .A3(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1332gat));
  OR3_X1    g502(.A1(new_n697_), .A2(G64gat), .A3(new_n658_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n691_), .A2(new_n401_), .A3(new_n693_), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(G64gat), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(G64gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(G1333gat));
  NAND3_X1  g508(.A1(new_n691_), .A2(new_n244_), .A3(new_n693_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT49), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(G71gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G71gat), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n244_), .A2(new_n204_), .ZN(new_n714_));
  OAI22_X1  g513(.A1(new_n712_), .A2(new_n713_), .B1(new_n697_), .B2(new_n714_), .ZN(G1334gat));
  OR3_X1    g514(.A1(new_n697_), .A2(G78gat), .A3(new_n430_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n691_), .A2(new_n352_), .A3(new_n693_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT50), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(new_n718_), .A3(G78gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n717_), .B2(G78gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1335gat));
  AND2_X1   g520(.A1(new_n696_), .A2(new_n652_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n303_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n642_), .A2(KEYINPUT112), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n642_), .A2(KEYINPUT112), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n588_), .A2(new_n460_), .A3(new_n651_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n303_), .A2(G85gat), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT113), .Z(new_n730_));
  AOI21_X1  g529(.A(new_n723_), .B1(new_n728_), .B2(new_n730_), .ZN(G1336gat));
  AOI21_X1  g530(.A(G92gat), .B1(new_n722_), .B2(new_n401_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n658_), .A2(new_n496_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n728_), .B2(new_n733_), .ZN(G1337gat));
  OAI21_X1  g533(.A(G99gat), .B1(new_n727_), .B2(new_n243_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n722_), .A2(new_n244_), .A3(new_n493_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT114), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT51), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n740_), .A3(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1338gat));
  NAND3_X1  g541(.A1(new_n722_), .A2(new_n492_), .A3(new_n352_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n726_), .A2(new_n352_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT115), .B1(new_n745_), .B2(new_n492_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n665_), .A2(new_n666_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n747_), .B(G106gat), .C1(new_n748_), .C2(new_n744_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n746_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n743_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT53), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n743_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1339gat));
  INV_X1    g556(.A(KEYINPUT59), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n554_), .A2(new_n461_), .A3(new_n588_), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n460_), .A2(new_n583_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n574_), .A2(new_n564_), .A3(new_n576_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n577_), .B1(new_n764_), .B2(KEYINPUT55), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n766_), .B(new_n564_), .C1(new_n574_), .C2(new_n576_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n561_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n764_), .A2(KEYINPUT55), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n581_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n767_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n561_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n763_), .B1(new_n770_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT117), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n452_), .A2(new_n448_), .A3(new_n454_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n458_), .B1(new_n453_), .B2(new_n449_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT118), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n458_), .B2(new_n455_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n578_), .A2(new_n583_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n776_), .B2(KEYINPUT117), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT57), .B(new_n550_), .C1(new_n778_), .C2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n768_), .A2(new_n769_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n561_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n783_), .A2(new_n583_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT119), .B(new_n788_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n770_), .B2(new_n775_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT58), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n796_), .A3(new_n640_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n460_), .B(new_n583_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n798_), .A2(new_n799_), .B1(new_n784_), .B2(new_n783_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n597_), .B1(new_n800_), .B2(new_n777_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n787_), .B(new_n797_), .C1(new_n801_), .C2(KEYINPUT57), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n762_), .B1(new_n802_), .B2(new_n482_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n599_), .A2(new_n303_), .A3(new_n244_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n758_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n787_), .A2(new_n797_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n798_), .A2(new_n799_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(new_n777_), .A3(new_n785_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT57), .B1(new_n808_), .B2(new_n550_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n482_), .B1(new_n806_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n761_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n804_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(KEYINPUT59), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n461_), .B1(new_n805_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(G113gat), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n460_), .A2(new_n815_), .ZN(new_n817_));
  OAI22_X1  g616(.A1(new_n814_), .A2(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(G1340gat));
  AOI21_X1  g617(.A(new_n588_), .B1(new_n805_), .B2(new_n813_), .ZN(new_n819_));
  INV_X1    g618(.A(G120gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT120), .B1(new_n820_), .B2(KEYINPUT60), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n588_), .B2(KEYINPUT60), .ZN(new_n822_));
  MUX2_X1   g621(.A(KEYINPUT120), .B(new_n821_), .S(new_n822_), .Z(new_n823_));
  OAI22_X1  g622(.A1(new_n819_), .A2(new_n820_), .B1(new_n816_), .B2(new_n823_), .ZN(G1341gat));
  NAND2_X1  g623(.A1(new_n805_), .A2(new_n813_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n482_), .A2(KEYINPUT121), .ZN(new_n826_));
  MUX2_X1   g625(.A(KEYINPUT121), .B(new_n826_), .S(G127gat), .Z(new_n827_));
  INV_X1    g626(.A(G127gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n811_), .A2(new_n651_), .A3(new_n812_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n825_), .A2(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(G1342gat));
  XOR2_X1   g629(.A(KEYINPUT122), .B(G134gat), .Z(new_n831_));
  NAND2_X1  g630(.A1(new_n640_), .A2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT123), .ZN(new_n833_));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n811_), .A2(new_n597_), .A3(new_n812_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n825_), .A2(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(G1343gat));
  AND2_X1   g635(.A1(new_n432_), .A2(new_n303_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n811_), .A2(new_n243_), .A3(new_n460_), .A4(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g638(.A1(new_n811_), .A2(new_n243_), .A3(new_n587_), .A4(new_n837_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g640(.A1(new_n811_), .A2(new_n243_), .A3(new_n651_), .A4(new_n837_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT61), .B(G155gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1346gat));
  NOR2_X1   g643(.A1(new_n803_), .A2(new_n244_), .ZN(new_n845_));
  INV_X1    g644(.A(G162gat), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n597_), .A4(new_n837_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n845_), .A2(new_n640_), .A3(new_n837_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n846_), .ZN(G1347gat));
  INV_X1    g648(.A(KEYINPUT22), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n305_), .A2(new_n352_), .A3(new_n658_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n811_), .A2(new_n850_), .A3(new_n460_), .A4(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n854_));
  INV_X1    g653(.A(new_n851_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n803_), .A2(new_n461_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n856_), .B2(new_n850_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n214_), .B1(new_n856_), .B2(new_n854_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n853_), .B1(new_n857_), .B2(new_n858_), .ZN(G1348gat));
  NOR2_X1   g658(.A1(new_n803_), .A2(new_n855_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n587_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g661(.A(new_n860_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n863_), .A2(new_n207_), .A3(new_n482_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G183gat), .B1(new_n860_), .B2(new_n651_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1350gat));
  OAI21_X1  g665(.A(G190gat), .B1(new_n863_), .B2(new_n637_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n860_), .A2(new_n208_), .A3(new_n597_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1351gat));
  NOR3_X1   g668(.A1(new_n430_), .A2(new_n303_), .A3(new_n658_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n811_), .A2(new_n243_), .A3(new_n460_), .A4(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n872_));
  NOR2_X1   g671(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT125), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n871_), .A2(new_n872_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1352gat));
  NAND2_X1  g676(.A1(new_n811_), .A2(new_n243_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n870_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n587_), .A3(new_n881_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n878_), .A2(new_n588_), .A3(new_n879_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT126), .B(G204gat), .Z(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1353gat));
  XNOR2_X1  g684(.A(KEYINPUT63), .B(G211gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n880_), .A2(new_n651_), .A3(new_n886_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n878_), .A2(new_n482_), .A3(new_n879_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(G1354gat));
  NAND2_X1  g689(.A1(new_n880_), .A2(new_n597_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT127), .B(G218gat), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n637_), .A2(new_n892_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n891_), .A2(new_n892_), .B1(new_n880_), .B2(new_n893_), .ZN(G1355gat));
endmodule


