//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n205_), .B(KEYINPUT36), .Z(new_n206_));
  XNOR2_X1  g005(.A(G85gat), .B(G92gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT9), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT10), .B(G99gat), .Z(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT9), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n209_), .A2(new_n212_), .A3(new_n215_), .A4(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AOI211_X1 g024(.A(KEYINPUT8), .B(new_n207_), .C1(new_n225_), .C2(new_n220_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n211_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n218_), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n222_), .B(new_n230_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n227_), .B1(new_n233_), .B2(new_n208_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n221_), .B1(new_n226_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G29gat), .B(G36gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G43gat), .B(G50gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n236_), .B(KEYINPUT69), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n235_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT35), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G232gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT34), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n245_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n235_), .A2(KEYINPUT65), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n252_), .B(new_n221_), .C1(new_n226_), .C2(new_n234_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n241_), .A2(new_n243_), .A3(KEYINPUT15), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT15), .B1(new_n241_), .B2(new_n243_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n251_), .B(new_n253_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n249_), .A2(new_n246_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n257_), .A2(new_n258_), .ZN(new_n261_));
  OAI211_X1 g060(.A(KEYINPUT71), .B(new_n206_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n259_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT71), .B1(new_n267_), .B2(new_n206_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n202_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n206_), .B(KEYINPUT70), .Z(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(KEYINPUT37), .A3(new_n265_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G1gat), .B(G8gat), .ZN(new_n275_));
  INV_X1    g074(.A(G1gat), .ZN(new_n276_));
  OR2_X1    g075(.A1(KEYINPUT72), .A2(G8gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(KEYINPUT72), .A2(G8gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT14), .ZN(new_n280_));
  OR3_X1    g079(.A1(new_n279_), .A2(KEYINPUT73), .A3(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT73), .B1(new_n279_), .B2(new_n280_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G15gat), .B(G22gat), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n275_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n275_), .ZN(new_n287_));
  AOI211_X1 g086(.A(new_n284_), .B(new_n287_), .C1(new_n281_), .C2(new_n282_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G57gat), .B(G64gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G71gat), .B(G78gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT11), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(KEYINPUT11), .ZN(new_n293_));
  INV_X1    g092(.A(new_n291_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n290_), .A2(KEYINPUT11), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n292_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G231gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n289_), .B(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G127gat), .B(G155gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G183gat), .B(G211gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT17), .B1(new_n300_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n305_), .B1(new_n300_), .B2(KEYINPUT75), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OAI211_X1 g107(.A(KEYINPUT17), .B(new_n305_), .C1(new_n300_), .C2(KEYINPUT75), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n274_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT76), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT98), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G228gat), .A2(G233gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT90), .ZN(new_n316_));
  INV_X1    g115(.A(G141gat), .ZN(new_n317_));
  INV_X1    g116(.A(G148gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(G155gat), .B2(G162gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT91), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(G155gat), .A3(G162gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT92), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT92), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n320_), .B1(new_n323_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n316_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n319_), .A2(KEYINPUT3), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n333_), .B2(new_n315_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n332_), .B1(new_n334_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT29), .B1(new_n330_), .B2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G197gat), .B(G204gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT95), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G211gat), .B(G218gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT21), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n343_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n341_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n314_), .B1(new_n340_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT96), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT96), .B1(new_n347_), .B2(new_n350_), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n314_), .B(KEYINPUT94), .Z(new_n356_));
  AND3_X1   g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n323_), .A2(new_n329_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n320_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n339_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT93), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT93), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n330_), .B2(new_n339_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n364_), .A3(KEYINPUT29), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n352_), .B1(new_n357_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT97), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n352_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n365_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT97), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n367_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n369_), .A2(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n362_), .A2(new_n364_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT28), .B1(new_n377_), .B2(KEYINPUT29), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT29), .B1(new_n362_), .B2(new_n364_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G22gat), .B(G50gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n382_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n379_), .A2(new_n380_), .ZN(new_n385_));
  AOI211_X1 g184(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n362_), .C2(new_n364_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n370_), .B(new_n368_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n313_), .B1(new_n376_), .B2(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n383_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n391_), .A2(KEYINPUT98), .A3(new_n369_), .A4(new_n375_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n347_), .A2(new_n350_), .A3(KEYINPUT96), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n344_), .A2(new_n349_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT21), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n353_), .B1(new_n396_), .B2(new_n346_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G169gat), .A2(G176gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT22), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(G169gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(KEYINPUT87), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT87), .B1(new_n402_), .B2(G169gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(G176gat), .B1(new_n402_), .B2(G169gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n401_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT79), .B(G183gat), .Z(new_n410_));
  INV_X1    g209(.A(G190gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G183gat), .A2(G190gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n414_), .A2(KEYINPUT23), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT86), .B(KEYINPUT23), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n409_), .A2(KEYINPUT88), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(KEYINPUT88), .B2(new_n409_), .ZN(new_n419_));
  INV_X1    g218(.A(G169gat), .ZN(new_n420_));
  INV_X1    g219(.A(G176gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(KEYINPUT83), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(G169gat), .B2(G176gat), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(KEYINPUT24), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n413_), .A2(KEYINPUT23), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n416_), .B2(new_n413_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n410_), .A2(KEYINPUT25), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n410_), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT25), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n434_), .A2(KEYINPUT81), .ZN(new_n435_));
  INV_X1    g234(.A(G183gat), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(KEYINPUT81), .B2(new_n434_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT26), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT82), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n439_), .B2(new_n411_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT82), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n435_), .A2(new_n437_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n432_), .A2(new_n433_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n425_), .A2(new_n401_), .A3(KEYINPUT24), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n444_), .A2(new_n445_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n429_), .B(new_n443_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n419_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n398_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT19), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n404_), .A2(new_n407_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(G183gat), .A2(G190gat), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n401_), .B(new_n455_), .C1(new_n428_), .C2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n399_), .A2(KEYINPUT24), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n458_), .A2(KEYINPUT100), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(KEYINPUT100), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n425_), .A3(new_n460_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n461_), .B(new_n417_), .C1(KEYINPUT24), .C2(new_n425_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT26), .B(G190gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT99), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT25), .B(G183gat), .Z(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n457_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n450_), .B(new_n454_), .C1(new_n351_), .C2(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n448_), .B(new_n419_), .C1(new_n394_), .C2(new_n397_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n453_), .B1(new_n468_), .B2(new_n351_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT101), .B1(new_n472_), .B2(new_n452_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT101), .ZN(new_n474_));
  INV_X1    g273(.A(new_n452_), .ZN(new_n475_));
  AOI211_X1 g274(.A(new_n474_), .B(new_n475_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n469_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT18), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G64gat), .B(G92gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G127gat), .B(G134gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT89), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G113gat), .B(G120gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n361_), .A3(new_n360_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n362_), .A2(new_n364_), .A3(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G225gat), .A2(G233gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G29gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(G85gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT0), .B(G57gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT4), .ZN(new_n498_));
  INV_X1    g297(.A(new_n491_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n499_), .B1(new_n490_), .B2(KEYINPUT4), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n492_), .B(new_n497_), .C1(new_n498_), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT33), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT33), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT4), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n505_), .B(new_n491_), .C1(KEYINPUT4), .C2(new_n490_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n489_), .A2(new_n490_), .A3(new_n499_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n507_), .A2(new_n496_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n501_), .A2(new_n504_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n481_), .B(new_n469_), .C1(new_n473_), .C2(new_n476_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n483_), .A2(new_n503_), .A3(new_n509_), .A4(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n373_), .A2(new_n367_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n388_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n383_), .A2(new_n387_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n481_), .A2(KEYINPUT32), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n469_), .B(new_n516_), .C1(new_n473_), .C2(new_n476_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n470_), .A2(new_n475_), .A3(new_n471_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n468_), .B2(new_n351_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n398_), .B2(new_n449_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n518_), .B1(new_n521_), .B2(new_n475_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(KEYINPUT32), .A3(new_n481_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n498_), .A2(new_n500_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n497_), .B1(new_n524_), .B2(new_n492_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n517_), .B(new_n523_), .C1(new_n525_), .C2(new_n502_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n393_), .A2(new_n511_), .A3(new_n515_), .A4(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G71gat), .B(G99gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G43gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n449_), .B(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n530_), .A2(new_n488_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n488_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G227gat), .A2(G233gat), .ZN(new_n533_));
  INV_X1    g332(.A(G15gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT30), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT31), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OR3_X1    g337(.A1(new_n531_), .A2(new_n532_), .A3(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n538_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT27), .B1(new_n483_), .B2(new_n510_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n524_), .A2(new_n492_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n496_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n501_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n522_), .A2(new_n482_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n510_), .A2(KEYINPUT27), .A3(new_n546_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n542_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n390_), .A2(new_n392_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n527_), .B(new_n541_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n542_), .A2(new_n547_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n545_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n541_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n551_), .A2(new_n549_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n297_), .B(new_n221_), .C1(new_n226_), .C2(new_n234_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT66), .B(KEYINPUT12), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n295_), .A2(new_n296_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n235_), .A2(new_n292_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT12), .B(new_n292_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n251_), .A2(new_n253_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n561_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT67), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n561_), .A2(new_n564_), .A3(KEYINPUT67), .A4(new_n565_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n226_), .A2(new_n234_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT64), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n221_), .A4(new_n297_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n556_), .A2(KEYINPUT64), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n560_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(G230gat), .A3(G233gat), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n568_), .A2(new_n569_), .A3(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT5), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n580_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n568_), .A2(new_n569_), .A3(new_n575_), .A4(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n583_), .A2(KEYINPUT68), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(KEYINPUT68), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n581_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n583_), .B(KEYINPUT68), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(KEYINPUT13), .A3(new_n581_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n283_), .A2(new_n285_), .A3(new_n275_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n282_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n279_), .A2(KEYINPUT73), .A3(new_n280_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n285_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n287_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n592_), .B(new_n596_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G229gat), .A2(G233gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n244_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT78), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n596_), .A2(new_n244_), .A3(new_n592_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT77), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n598_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n289_), .A2(KEYINPUT77), .A3(new_n244_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n597_), .A2(KEYINPUT78), .A3(new_n600_), .A4(new_n598_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n603_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G169gat), .B(G197gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n603_), .A2(new_n609_), .A3(new_n610_), .A4(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n591_), .A2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n555_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n312_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n276_), .A3(new_n545_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT103), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT38), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n625_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n620_), .B(KEYINPUT104), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n266_), .A2(new_n268_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n550_), .B2(new_n554_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n628_), .A2(new_n310_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n276_), .B1(new_n631_), .B2(new_n545_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT105), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n626_), .A2(new_n627_), .A3(new_n633_), .ZN(G1324gat));
  XNOR2_X1  g433(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n635_));
  INV_X1    g434(.A(new_n551_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(G8gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT39), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n622_), .A2(new_n277_), .A3(new_n278_), .A4(new_n636_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n635_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n638_), .A2(KEYINPUT39), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n637_), .B2(G8gat), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n640_), .B(new_n635_), .C1(new_n642_), .C2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n641_), .A2(new_n646_), .ZN(G1325gat));
  AOI21_X1  g446(.A(new_n534_), .B1(new_n631_), .B2(new_n553_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT41), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n622_), .A2(new_n534_), .A3(new_n553_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n549_), .B(KEYINPUT107), .Z(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n631_), .B2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT42), .Z(new_n656_));
  NAND3_X1  g455(.A1(new_n622_), .A2(new_n652_), .A3(new_n654_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1327gat));
  INV_X1    g457(.A(new_n629_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n310_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n621_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G29gat), .B1(new_n661_), .B2(new_n545_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n310_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n274_), .B1(new_n550_), .B2(new_n554_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(KEYINPUT108), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n274_), .B(new_n668_), .C1(new_n550_), .C2(new_n554_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n628_), .B(new_n663_), .C1(new_n666_), .C2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n668_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n555_), .A2(new_n273_), .A3(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n675_), .A2(KEYINPUT44), .A3(new_n628_), .A4(new_n663_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n672_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n545_), .A2(G29gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n662_), .B1(new_n677_), .B2(new_n678_), .ZN(G1328gat));
  NAND3_X1  g478(.A1(new_n672_), .A2(new_n636_), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G36gat), .ZN(new_n681_));
  NOR2_X1   g480(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n551_), .A2(G36gat), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n661_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT45), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n661_), .A2(new_n686_), .A3(new_n683_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n682_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n681_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1329gat));
  NAND4_X1  g490(.A1(new_n672_), .A2(new_n676_), .A3(G43gat), .A4(new_n553_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n661_), .A2(new_n553_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(G43gat), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g494(.A1(new_n653_), .A2(G50gat), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT112), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n661_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n699_));
  INV_X1    g498(.A(new_n549_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n672_), .A2(new_n676_), .A3(new_n699_), .A4(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(G50gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n672_), .A2(new_n700_), .A3(new_n676_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT110), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT111), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  AND4_X1   g504(.A1(KEYINPUT111), .A2(new_n704_), .A3(G50gat), .A4(new_n701_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n698_), .B1(new_n705_), .B2(new_n706_), .ZN(G1331gat));
  INV_X1    g506(.A(new_n591_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n708_), .A2(new_n618_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n555_), .A2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n312_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n545_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n630_), .A2(new_n310_), .A3(new_n709_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n552_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1332gat));
  OAI21_X1  g515(.A(G64gat), .B1(new_n714_), .B2(new_n551_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT48), .ZN(new_n718_));
  INV_X1    g517(.A(G64gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n711_), .A2(new_n719_), .A3(new_n636_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n714_), .B2(new_n541_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  INV_X1    g522(.A(G71gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n711_), .A2(new_n724_), .A3(new_n553_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1334gat));
  OAI21_X1  g525(.A(G78gat), .B1(new_n714_), .B2(new_n653_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT50), .ZN(new_n728_));
  INV_X1    g527(.A(G78gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n711_), .A2(new_n729_), .A3(new_n654_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1335gat));
  NAND3_X1  g530(.A1(new_n675_), .A2(new_n663_), .A3(new_n709_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G85gat), .B1(new_n732_), .B2(new_n552_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n710_), .A2(new_n660_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n213_), .A3(new_n545_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1336gat));
  OAI21_X1  g535(.A(G92gat), .B1(new_n732_), .B2(new_n551_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n214_), .A3(new_n636_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1337gat));
  OAI21_X1  g538(.A(G99gat), .B1(new_n732_), .B2(new_n541_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT114), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT51), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n734_), .A2(new_n210_), .A3(new_n553_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT113), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT113), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n740_), .B(new_n742_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n741_), .A2(KEYINPUT51), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(G1338gat));
  NAND3_X1  g547(.A1(new_n734_), .A2(new_n211_), .A3(new_n700_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n675_), .A2(new_n663_), .A3(new_n700_), .A4(new_n709_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(G106gat), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n751_), .B1(new_n750_), .B2(G106gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n749_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g555(.A1(new_n551_), .A2(new_n549_), .A3(new_n545_), .A4(new_n553_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT58), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n568_), .A2(new_n760_), .A3(new_n569_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n565_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n561_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(KEYINPUT55), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n759_), .B1(new_n765_), .B2(new_n580_), .ZN(new_n766_));
  AOI211_X1 g565(.A(KEYINPUT56), .B(new_n582_), .C1(new_n761_), .C2(new_n764_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n606_), .A2(new_n598_), .A3(new_n608_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n597_), .A2(new_n607_), .A3(new_n600_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n615_), .A3(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n617_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(KEYINPUT116), .C1(new_n584_), .C2(new_n585_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n768_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT116), .B1(new_n589_), .B2(new_n772_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT117), .B(new_n758_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n772_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(new_n773_), .A3(new_n768_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n758_), .B1(new_n781_), .B2(KEYINPUT117), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n777_), .A2(new_n782_), .A3(new_n274_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n765_), .A2(new_n580_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(KEYINPUT56), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n582_), .B1(new_n761_), .B2(new_n764_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n759_), .B1(new_n787_), .B2(KEYINPUT115), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n786_), .A2(new_n788_), .A3(new_n618_), .A4(new_n589_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n586_), .A2(new_n772_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n629_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT57), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n663_), .B1(new_n783_), .B2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n269_), .A2(new_n619_), .A3(new_n310_), .A4(new_n272_), .ZN(new_n794_));
  OR3_X1    g593(.A1(new_n794_), .A2(KEYINPUT54), .A3(new_n591_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT54), .B1(new_n794_), .B2(new_n591_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n757_), .B1(new_n793_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT118), .ZN(new_n799_));
  INV_X1    g598(.A(new_n757_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n791_), .A2(KEYINPUT57), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n802_), .B(new_n629_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT117), .B1(new_n774_), .B2(new_n775_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT58), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n273_), .A3(new_n776_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n310_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n797_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n800_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n799_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(G113gat), .B1(new_n813_), .B2(new_n618_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n798_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n810_), .A2(new_n817_), .A3(KEYINPUT59), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n810_), .B2(KEYINPUT59), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n816_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT120), .B(new_n816_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n618_), .A2(KEYINPUT121), .A3(G113gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(KEYINPUT121), .B2(G113gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n814_), .B1(new_n824_), .B2(new_n826_), .ZN(G1340gat));
  NOR2_X1   g626(.A1(new_n708_), .A2(KEYINPUT60), .ZN(new_n828_));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  MUX2_X1   g628(.A(KEYINPUT60), .B(new_n828_), .S(new_n829_), .Z(new_n830_));
  NAND3_X1  g629(.A1(new_n799_), .A2(new_n812_), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n591_), .B1(new_n810_), .B2(KEYINPUT59), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT119), .B1(new_n798_), .B2(new_n815_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n810_), .A2(new_n817_), .A3(KEYINPUT59), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n835_), .B2(new_n829_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT122), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n831_), .C1(new_n835_), .C2(new_n829_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1341gat));
  AOI21_X1  g639(.A(G127gat), .B1(new_n813_), .B2(new_n310_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n310_), .A2(G127gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n824_), .B2(new_n842_), .ZN(G1342gat));
  AOI21_X1  g642(.A(G134gat), .B1(new_n813_), .B2(new_n629_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n273_), .A2(G134gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n824_), .B2(new_n845_), .ZN(G1343gat));
  NAND2_X1  g645(.A1(new_n793_), .A2(new_n797_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n636_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n700_), .A3(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n619_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n317_), .ZN(G1344gat));
  NOR2_X1   g650(.A1(new_n849_), .A2(new_n708_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(new_n318_), .ZN(G1345gat));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n849_), .B2(new_n663_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n808_), .A2(new_n809_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n549_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n857_), .A2(KEYINPUT123), .A3(new_n310_), .A4(new_n848_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1346gat));
  OAI21_X1  g660(.A(G162gat), .B1(new_n849_), .B2(new_n274_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n659_), .A2(G162gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n849_), .B2(new_n863_), .ZN(G1347gat));
  NAND3_X1  g663(.A1(new_n636_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n653_), .B(new_n866_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n420_), .A2(KEYINPUT22), .ZN(new_n868_));
  OR4_X1    g667(.A1(new_n619_), .A2(new_n867_), .A3(new_n403_), .A4(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n847_), .A2(new_n618_), .A3(new_n653_), .A4(new_n866_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(G169gat), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n870_), .B(G169gat), .C1(new_n867_), .C2(new_n619_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n869_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n869_), .B(new_n877_), .C1(new_n872_), .C2(new_n874_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1348gat));
  OR2_X1    g678(.A1(new_n867_), .A2(new_n708_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n856_), .A2(new_n700_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n865_), .A2(new_n421_), .A3(new_n708_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n880_), .A2(new_n421_), .B1(new_n881_), .B2(new_n882_), .ZN(G1349gat));
  NOR2_X1   g682(.A1(new_n856_), .A2(new_n654_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n866_), .A2(new_n310_), .A3(new_n466_), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT125), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n884_), .A2(KEYINPUT125), .A3(new_n885_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n881_), .A2(new_n310_), .A3(new_n866_), .ZN(new_n888_));
  AOI211_X1 g687(.A(new_n886_), .B(new_n887_), .C1(new_n410_), .C2(new_n888_), .ZN(G1350gat));
  OAI21_X1  g688(.A(G190gat), .B1(new_n867_), .B2(new_n274_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n659_), .A2(new_n465_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n867_), .B2(new_n891_), .ZN(G1351gat));
  NAND3_X1  g691(.A1(new_n636_), .A2(new_n552_), .A3(new_n541_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n857_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n619_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n708_), .ZN(new_n898_));
  AND2_X1   g697(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n899_));
  NOR2_X1   g698(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n898_), .B2(new_n900_), .ZN(G1353gat));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  AND2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n895_), .A2(new_n663_), .A3(new_n903_), .A4(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n895_), .B2(new_n663_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n906_), .A2(KEYINPUT127), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(KEYINPUT127), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n907_), .B2(new_n908_), .ZN(G1354gat));
  OAI21_X1  g708(.A(G218gat), .B1(new_n895_), .B2(new_n274_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n659_), .A2(G218gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n895_), .B2(new_n911_), .ZN(G1355gat));
endmodule


