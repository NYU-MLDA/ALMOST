//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT66), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n206_));
  XOR2_X1   g005(.A(G71gat), .B(G78gat), .Z(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT10), .B(G99gat), .Z(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G85gat), .B(G92gat), .Z(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n216_));
  INV_X1    g015(.A(G85gat), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  OR3_X1    g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT9), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT6), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n214_), .A2(new_n216_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(new_n221_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n215_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n215_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n225_), .B1(KEYINPUT65), .B2(new_n221_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n221_), .A2(KEYINPUT65), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n229_), .B1(new_n233_), .B2(new_n228_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n209_), .A2(new_n222_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n222_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n206_), .A2(new_n207_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n206_), .A2(new_n207_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n238_), .B2(new_n205_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G230gat), .A2(G233gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G120gat), .B(G148gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G176gat), .B(G204gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n236_), .A2(KEYINPUT12), .A3(new_n239_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT12), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n240_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n236_), .A2(KEYINPUT67), .A3(new_n239_), .A4(KEYINPUT12), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n253_), .A2(new_n255_), .A3(new_n235_), .A4(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n244_), .B(new_n250_), .C1(new_n257_), .C2(new_n243_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n236_), .A2(new_n239_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n254_), .B2(new_n240_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n262_), .A2(new_n242_), .A3(new_n256_), .A4(new_n253_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n263_), .A2(KEYINPUT69), .A3(new_n244_), .A4(new_n250_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n244_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n249_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n265_), .A2(KEYINPUT13), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT13), .B1(new_n265_), .B2(new_n267_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n202_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n267_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT13), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n265_), .A2(KEYINPUT13), .A3(new_n267_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(KEYINPUT70), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G29gat), .B(G36gat), .Z(new_n277_));
  XOR2_X1   g076(.A(G43gat), .B(G50gat), .Z(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  XNOR2_X1  g078(.A(G15gat), .B(G22gat), .ZN(new_n280_));
  INV_X1    g079(.A(G1gat), .ZN(new_n281_));
  INV_X1    g080(.A(G8gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT14), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G1gat), .B(G8gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n279_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT78), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(G229gat), .A3(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n279_), .B(KEYINPUT15), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n286_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G229gat), .A2(G233gat), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n292_), .B(new_n293_), .C1(new_n286_), .C2(new_n279_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G113gat), .B(G141gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT79), .ZN(new_n296_));
  XOR2_X1   g095(.A(G169gat), .B(G197gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n289_), .A2(new_n294_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n289_), .B2(new_n294_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n276_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G232gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT35), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT72), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n279_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n234_), .A2(new_n222_), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT74), .B1(new_n308_), .B2(new_n309_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n290_), .B1(new_n234_), .B2(new_n222_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n312_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G190gat), .B(G218gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT73), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G134gat), .B(G162gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(KEYINPUT36), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n291_), .A2(new_n236_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n326_), .A2(new_n311_), .A3(new_n314_), .A4(new_n315_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(KEYINPUT36), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n318_), .A2(new_n325_), .A3(new_n327_), .A4(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n325_), .B1(new_n318_), .B2(new_n327_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n329_), .B1(new_n330_), .B2(KEYINPUT75), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n332_));
  AOI211_X1 g131(.A(new_n332_), .B(new_n325_), .C1(new_n318_), .C2(new_n327_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n305_), .B(KEYINPUT37), .C1(new_n331_), .C2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n318_), .A2(new_n327_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n324_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n329_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n337_), .A2(KEYINPUT37), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n332_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n330_), .A2(KEYINPUT75), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n329_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n305_), .B1(new_n342_), .B2(KEYINPUT37), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n286_), .ZN(new_n345_));
  INV_X1    g144(.A(G231gat), .ZN(new_n346_));
  INV_X1    g145(.A(G233gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n209_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n239_), .A2(new_n348_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n345_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n209_), .A2(new_n349_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n239_), .A2(new_n348_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT77), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n286_), .A3(new_n353_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G127gat), .B(G155gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT16), .ZN(new_n363_));
  XOR2_X1   g162(.A(G183gat), .B(G211gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT17), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n365_), .B(KEYINPUT17), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n356_), .A2(new_n360_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n344_), .A2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT88), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT90), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT89), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT2), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384_));
  INV_X1    g183(.A(G141gat), .ZN(new_n385_));
  INV_X1    g184(.A(G148gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n377_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n378_), .A2(new_n380_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT89), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(KEYINPUT90), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n376_), .B1(new_n391_), .B2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n378_), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n375_), .B(KEYINPUT1), .Z(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(new_n374_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n398_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405_));
  XOR2_X1   g204(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n376_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n383_), .A2(new_n377_), .A3(new_n390_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT90), .B1(new_n395_), .B2(new_n396_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n403_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n406_), .B1(new_n414_), .B2(KEYINPUT29), .ZN(new_n415_));
  INV_X1    g214(.A(G228gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(new_n347_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(KEYINPUT29), .ZN(new_n419_));
  XOR2_X1   g218(.A(G211gat), .B(G218gat), .Z(new_n420_));
  OR2_X1    g219(.A1(G197gat), .A2(G204gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G197gat), .A2(G204gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT21), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(KEYINPUT92), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n420_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n423_), .A2(new_n424_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G211gat), .B(G218gat), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n429_), .A2(new_n421_), .A3(new_n422_), .A4(new_n425_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n418_), .B1(new_n419_), .B2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n404_), .A2(new_n405_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n427_), .A2(KEYINPUT93), .A3(new_n428_), .A4(new_n430_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n418_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n408_), .B(new_n415_), .C1(new_n433_), .C2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n417_), .B1(new_n434_), .B2(new_n431_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n415_), .A2(new_n408_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n442_), .B(new_n443_), .C1(new_n434_), .C2(new_n439_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G22gat), .B(G50gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n441_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G183gat), .A2(G190gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT23), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n456_), .B(new_n457_), .C1(G183gat), .C2(G190gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459_));
  OR2_X1    g258(.A1(KEYINPUT83), .A2(G176gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(KEYINPUT83), .A2(G176gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT22), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(G169gat), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n460_), .B(new_n461_), .C1(new_n463_), .C2(KEYINPUT82), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465_));
  INV_X1    g264(.A(G169gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT22), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n462_), .A2(G169gat), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n465_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n458_), .B(new_n459_), .C1(new_n464_), .C2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(G169gat), .A2(G176gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(KEYINPUT24), .A3(new_n459_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT25), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT25), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n477_));
  INV_X1    g276(.A(G190gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT26), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT26), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G190gat), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n475_), .A2(new_n477_), .A3(new_n479_), .A4(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n454_), .A2(KEYINPUT23), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n455_), .A2(G183gat), .A3(G190gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT24), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n483_), .A2(new_n484_), .B1(new_n485_), .B2(new_n471_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n473_), .B(new_n482_), .C1(new_n486_), .C2(KEYINPUT81), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n471_), .A2(new_n485_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n455_), .B1(G183gat), .B2(G190gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n454_), .A2(KEYINPUT23), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT81), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n470_), .B1(new_n487_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT84), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n496_), .B(new_n470_), .C1(new_n487_), .C2(new_n493_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G227gat), .A2(G233gat), .ZN(new_n499_));
  INV_X1    g298(.A(G15gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT30), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n498_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G127gat), .B(G134gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT85), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT85), .ZN(new_n507_));
  INV_X1    g306(.A(G127gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(G134gat), .ZN(new_n509_));
  INV_X1    g308(.A(G134gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(G127gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n507_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G113gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(G120gat), .ZN(new_n514_));
  INV_X1    g313(.A(G120gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n515_), .A2(G113gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT86), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(G113gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(G120gat), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT86), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AND4_X1   g320(.A1(new_n506_), .A2(new_n512_), .A3(new_n517_), .A4(new_n521_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n506_), .A2(new_n512_), .B1(new_n517_), .B2(new_n521_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n504_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n506_), .A2(new_n512_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n517_), .A2(new_n521_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT87), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n503_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G71gat), .B(G99gat), .ZN(new_n530_));
  INV_X1    g329(.A(G43gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT31), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n529_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G1gat), .B(G29gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G85gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT0), .B(G57gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  INV_X1    g337(.A(KEYINPUT4), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n524_), .B(new_n527_), .C1(new_n403_), .C2(new_n398_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n525_), .A2(new_n526_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n506_), .A2(new_n512_), .A3(new_n517_), .A4(new_n521_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n412_), .A2(new_n543_), .A3(new_n413_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n539_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G225gat), .A2(G233gat), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n506_), .A2(new_n512_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n521_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n520_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n504_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n551_), .B1(new_n504_), .B2(new_n543_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT4), .B1(new_n552_), .B2(new_n414_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n545_), .A2(new_n546_), .A3(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n544_), .B1(new_n528_), .B2(new_n404_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n546_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n538_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT99), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(KEYINPUT4), .ZN(new_n560_));
  INV_X1    g359(.A(new_n546_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n553_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n538_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n564_), .A3(new_n556_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n558_), .A2(new_n559_), .A3(new_n565_), .ZN(new_n566_));
  OAI211_X1 g365(.A(KEYINPUT99), .B(new_n538_), .C1(new_n554_), .C2(new_n557_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n534_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT100), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n460_), .A2(new_n461_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n467_), .A2(new_n468_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(new_n459_), .A3(new_n458_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT25), .B(G183gat), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n479_), .A2(new_n481_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n473_), .A2(new_n456_), .A3(new_n457_), .A4(new_n488_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n575_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n571_), .B1(new_n582_), .B2(new_n432_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n495_), .A2(new_n436_), .A3(new_n437_), .A4(new_n497_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G226gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(new_n584_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT20), .B1(new_n582_), .B2(new_n432_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n498_), .A2(new_n593_), .A3(new_n438_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n593_), .B1(new_n498_), .B2(new_n438_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n592_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n590_), .B1(new_n596_), .B2(new_n587_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G8gat), .B(G36gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G64gat), .B(G92gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n570_), .B1(new_n597_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT27), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n588_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n497_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n482_), .A2(new_n473_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n491_), .A2(new_n492_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n486_), .A2(KEYINPUT81), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n496_), .B1(new_n610_), .B2(new_n470_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n438_), .B1(new_n606_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT96), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n498_), .A2(new_n593_), .A3(new_n438_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n591_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n605_), .B1(new_n615_), .B2(new_n588_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n604_), .B1(new_n616_), .B2(new_n602_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n589_), .B1(new_n615_), .B2(new_n588_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n602_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(KEYINPUT100), .A3(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n603_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n603_), .A2(new_n617_), .A3(KEYINPUT101), .A4(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n588_), .B(new_n592_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n605_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(new_n602_), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n602_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT103), .B1(new_n625_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n633_));
  INV_X1    g432(.A(new_n631_), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n633_), .B(new_n634_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n453_), .B(new_n569_), .C1(new_n632_), .C2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n558_), .A2(KEYINPUT33), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n638_), .B(new_n538_), .C1(new_n554_), .C2(new_n557_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n629_), .A2(new_n630_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n546_), .B1(new_n545_), .B2(new_n553_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n642_), .B(new_n564_), .C1(new_n555_), .C2(new_n546_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n640_), .A2(new_n641_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n627_), .A2(new_n628_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n602_), .A2(KEYINPUT32), .ZN(new_n646_));
  MUX2_X1   g445(.A(new_n597_), .B(new_n645_), .S(new_n646_), .Z(new_n647_));
  AOI22_X1  g446(.A1(new_n644_), .A2(KEYINPUT98), .B1(new_n568_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n640_), .A2(new_n641_), .A3(new_n649_), .A4(new_n643_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n452_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n566_), .A2(new_n567_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n452_), .ZN(new_n653_));
  AOI211_X1 g452(.A(new_n634_), .B(new_n653_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n534_), .B1(new_n651_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n636_), .A2(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n304_), .A2(new_n372_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT104), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n304_), .A2(new_n656_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n372_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n652_), .A2(G1gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n658_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n658_), .A2(KEYINPUT38), .A3(new_n662_), .A4(new_n663_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n303_), .A2(new_n371_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n337_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n636_), .B2(new_n655_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G1gat), .B1(new_n672_), .B2(new_n652_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n666_), .A2(new_n667_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1324gat));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n632_), .A2(new_n635_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n671_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  AND4_X1   g479(.A1(new_n677_), .A2(new_n679_), .A3(new_n680_), .A4(G8gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n282_), .B1(KEYINPUT106), .B2(KEYINPUT39), .ZN(new_n682_));
  AOI22_X1  g481(.A1(new_n679_), .A2(new_n682_), .B1(new_n677_), .B2(new_n680_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n658_), .A2(new_n662_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n678_), .A2(new_n282_), .ZN(new_n685_));
  OAI22_X1  g484(.A1(new_n681_), .A2(new_n683_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI221_X1 g487(.A(KEYINPUT40), .B1(new_n684_), .B2(new_n685_), .C1(new_n681_), .C2(new_n683_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1325gat));
  INV_X1    g489(.A(new_n534_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n500_), .B1(new_n671_), .B2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT41), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n657_), .A2(new_n500_), .A3(new_n691_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1326gat));
  OAI21_X1  g494(.A(G22gat), .B1(new_n672_), .B2(new_n453_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT42), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n453_), .A2(G22gat), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT107), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n657_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1327gat));
  INV_X1    g500(.A(new_n371_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n303_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n656_), .B2(new_n344_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n339_), .A2(new_n343_), .ZN(new_n706_));
  AOI211_X1 g505(.A(KEYINPUT43), .B(new_n706_), .C1(new_n636_), .C2(new_n655_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n703_), .B(KEYINPUT44), .C1(new_n705_), .C2(new_n707_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n710_), .A2(G29gat), .A3(new_n568_), .A4(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(G29gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n303_), .B1(new_n655_), .B2(new_n636_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n702_), .A2(new_n337_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n716_), .B2(new_n652_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n712_), .A2(new_n717_), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n710_), .A2(new_n678_), .A3(new_n711_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G36gat), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n632_), .A2(new_n635_), .A3(G36gat), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n714_), .A2(new_n721_), .A3(new_n715_), .A4(new_n722_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n304_), .A2(new_n656_), .A3(new_n715_), .A4(new_n722_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT108), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n723_), .A2(new_n725_), .A3(KEYINPUT45), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT45), .B1(new_n723_), .B2(new_n725_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n720_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n720_), .A2(KEYINPUT46), .A3(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1329gat));
  NAND4_X1  g532(.A1(new_n710_), .A2(G43gat), .A3(new_n691_), .A4(new_n711_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n531_), .B1(new_n716_), .B2(new_n534_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(G1330gat));
  NAND3_X1  g537(.A1(new_n710_), .A2(new_n452_), .A3(new_n711_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n739_), .A2(KEYINPUT110), .A3(G50gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT110), .B1(new_n739_), .B2(G50gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n453_), .A2(G50gat), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT111), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n740_), .A2(new_n741_), .B1(new_n716_), .B2(new_n743_), .ZN(G1331gat));
  NAND3_X1  g543(.A1(new_n368_), .A2(new_n301_), .A3(new_n370_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n276_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n670_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(G57gat), .A3(new_n568_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT113), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n656_), .A2(new_n301_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT112), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n270_), .A2(new_n275_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n372_), .A3(new_n568_), .ZN(new_n755_));
  INV_X1    g554(.A(G57gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n750_), .B1(new_n755_), .B2(new_n756_), .ZN(G1332gat));
  NAND2_X1  g556(.A1(new_n748_), .A2(new_n678_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G64gat), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT114), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n758_), .A2(new_n761_), .A3(G64gat), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n760_), .A2(KEYINPUT48), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n754_), .A2(new_n372_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n678_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n768_), .A2(G64gat), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n765_), .B(new_n766_), .C1(new_n767_), .C2(new_n769_), .ZN(G1333gat));
  NOR2_X1   g569(.A1(new_n534_), .A2(G71gat), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT115), .ZN(new_n772_));
  OAI21_X1  g571(.A(G71gat), .B1(new_n747_), .B2(new_n534_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(KEYINPUT49), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(KEYINPUT49), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n767_), .A2(new_n772_), .B1(new_n774_), .B2(new_n775_), .ZN(G1334gat));
  OR2_X1    g575(.A1(new_n453_), .A2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(G78gat), .B1(new_n747_), .B2(new_n453_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(KEYINPUT50), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(KEYINPUT50), .ZN(new_n780_));
  OAI22_X1  g579(.A1(new_n767_), .A2(new_n777_), .B1(new_n779_), .B2(new_n780_), .ZN(G1335gat));
  NOR3_X1   g580(.A1(new_n276_), .A2(new_n702_), .A3(new_n302_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n652_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n754_), .A2(new_n715_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n568_), .A2(new_n217_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(G1336gat));
  OAI21_X1  g586(.A(G92gat), .B1(new_n783_), .B2(new_n768_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n678_), .A2(new_n218_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n785_), .B2(new_n789_), .ZN(G1337gat));
  AND2_X1   g589(.A1(new_n691_), .A2(new_n210_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n752_), .A2(new_n753_), .A3(new_n715_), .A4(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n691_), .B(new_n782_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n793_), .A2(new_n794_), .A3(G99gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n793_), .B2(G99gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g597(.A1(new_n453_), .A2(G106gat), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n752_), .A2(new_n753_), .A3(new_n715_), .A4(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n452_), .B(new_n782_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(G106gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(G106gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n243_), .B2(KEYINPUT119), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n257_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n807_), .B2(new_n243_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n262_), .A2(new_n256_), .A3(new_n253_), .A4(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n249_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n809_), .A2(new_n811_), .A3(KEYINPUT56), .A4(new_n249_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n299_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n288_), .A2(new_n293_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n293_), .B1(new_n313_), .B2(new_n345_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n298_), .B1(new_n292_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n816_), .A2(new_n265_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n814_), .A2(new_n815_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(KEYINPUT58), .A3(new_n823_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n344_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT120), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n826_), .A2(new_n344_), .A3(new_n831_), .A4(new_n828_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n302_), .A2(new_n827_), .B1(new_n271_), .B2(new_n823_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n669_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n816_), .A2(new_n302_), .A3(new_n265_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n822_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT57), .B(new_n337_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n830_), .A2(new_n832_), .A3(new_n835_), .A4(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n371_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n745_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n368_), .A2(new_n301_), .A3(new_n370_), .A4(KEYINPUT117), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n706_), .A2(new_n273_), .A3(new_n845_), .A4(new_n274_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n841_), .B1(new_n846_), .B2(KEYINPUT54), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(KEYINPUT54), .ZN(new_n848_));
  AND4_X1   g647(.A1(new_n273_), .A2(new_n274_), .A3(new_n844_), .A4(new_n843_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n849_), .A2(KEYINPUT118), .A3(new_n850_), .A4(new_n706_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n848_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n840_), .A2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n678_), .A2(new_n452_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n534_), .A2(new_n652_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n835_), .A2(new_n829_), .A3(new_n838_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n371_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT122), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n862_), .A3(new_n371_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n852_), .A3(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n856_), .A2(KEYINPUT59), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n858_), .A2(KEYINPUT59), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n513_), .B1(new_n866_), .B2(new_n302_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n858_), .A2(KEYINPUT121), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n853_), .A2(new_n869_), .A3(new_n857_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n301_), .A2(G113gat), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n868_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT123), .B1(new_n867_), .B2(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n848_), .A2(new_n851_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n874_), .A2(new_n847_), .B1(new_n839_), .B2(new_n371_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT59), .B1(new_n875_), .B2(new_n856_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n864_), .A2(new_n865_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n302_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G113gat), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n868_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n873_), .A2(new_n882_), .ZN(G1340gat));
  AND2_X1   g682(.A1(new_n868_), .A2(new_n870_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n515_), .B1(new_n276_), .B2(KEYINPUT60), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n884_), .B(new_n885_), .C1(KEYINPUT60), .C2(new_n515_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n866_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G120gat), .B1(new_n887_), .B2(new_n276_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1341gat));
  OAI21_X1  g688(.A(G127gat), .B1(new_n887_), .B2(new_n371_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n884_), .A2(new_n508_), .A3(new_n702_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1342gat));
  OAI21_X1  g691(.A(G134gat), .B1(new_n887_), .B2(new_n706_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n884_), .A2(new_n510_), .A3(new_n669_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1343gat));
  NOR4_X1   g694(.A1(new_n678_), .A2(new_n652_), .A3(new_n453_), .A4(new_n691_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n853_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n301_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n385_), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n276_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n386_), .ZN(G1345gat));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n371_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT61), .B(G155gat), .Z(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n897_), .B2(new_n706_), .ZN(new_n905_));
  INV_X1    g704(.A(G162gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n669_), .A2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n897_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1347gat));
  NAND2_X1  g709(.A1(new_n678_), .A2(new_n569_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n452_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n864_), .A2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n466_), .B1(new_n913_), .B2(new_n302_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n914_), .A2(KEYINPUT62), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n573_), .A3(new_n302_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(KEYINPUT62), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(G1348gat));
  NAND2_X1  g717(.A1(new_n853_), .A2(new_n453_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n753_), .A2(G176gat), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n919_), .A2(new_n911_), .A3(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n913_), .A2(new_n753_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n572_), .ZN(G1349gat));
  OR3_X1    g722(.A1(new_n919_), .A2(new_n371_), .A3(new_n911_), .ZN(new_n924_));
  INV_X1    g723(.A(G183gat), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n702_), .A2(new_n578_), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n924_), .A2(new_n925_), .B1(new_n913_), .B2(new_n926_), .ZN(G1350gat));
  NAND4_X1  g726(.A1(new_n913_), .A2(new_n669_), .A3(new_n479_), .A4(new_n481_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n913_), .A2(new_n344_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n478_), .ZN(G1351gat));
  NAND3_X1  g729(.A1(new_n534_), .A2(new_n652_), .A3(new_n452_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT125), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n768_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n853_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n302_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g736(.A1(new_n934_), .A2(new_n276_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n938_), .B(new_n939_), .ZN(G1353gat));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n371_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n935_), .A2(new_n941_), .A3(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n941_), .B1(new_n935_), .B2(new_n942_), .ZN(new_n945_));
  OAI22_X1  g744(.A1(new_n944_), .A2(new_n945_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n946_));
  INV_X1    g745(.A(new_n945_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n947_), .A2(new_n948_), .A3(new_n943_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n946_), .A2(new_n949_), .ZN(G1354gat));
  OR3_X1    g749(.A1(new_n934_), .A2(G218gat), .A3(new_n337_), .ZN(new_n951_));
  OAI21_X1  g750(.A(G218gat), .B1(new_n934_), .B2(new_n706_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1355gat));
endmodule


