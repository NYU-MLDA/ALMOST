//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(G176gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR3_X1   g009(.A1(new_n210_), .A2(new_n205_), .A3(new_n204_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n207_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT25), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n213_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT26), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n212_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT83), .B(G176gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT22), .B(G169gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT84), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT84), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n210_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT85), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n203_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n220_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT86), .ZN(new_n235_));
  XOR2_X1   g034(.A(G71gat), .B(G99gat), .Z(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n235_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n239_), .B(new_n242_), .Z(new_n243_));
  XNOR2_X1  g042(.A(G15gat), .B(G43gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT31), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n239_), .B(new_n242_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n246_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G228gat), .ZN(new_n252_));
  INV_X1    g051(.A(G233gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G141gat), .ZN(new_n256_));
  INV_X1    g055(.A(G148gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n257_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(KEYINPUT1), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT87), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OR3_X1    g064(.A1(new_n261_), .A2(KEYINPUT88), .A3(KEYINPUT1), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT88), .B1(new_n261_), .B2(KEYINPUT1), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n263_), .A2(new_n264_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n259_), .B(new_n260_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT89), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(G141gat), .B2(G148gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT3), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n274_), .A2(new_n275_), .B1(new_n258_), .B2(KEYINPUT2), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT90), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n272_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n262_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n261_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n277_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n270_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT29), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT92), .ZN(new_n287_));
  INV_X1    g086(.A(G197gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(G204gat), .ZN(new_n289_));
  INV_X1    g088(.A(G204gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(KEYINPUT92), .A3(G197gat), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n289_), .B(new_n291_), .C1(G197gat), .C2(new_n290_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n286_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT93), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n286_), .A2(new_n292_), .A3(KEYINPUT93), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n292_), .A2(KEYINPUT21), .ZN(new_n298_));
  INV_X1    g097(.A(new_n284_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G197gat), .B(G204gat), .Z(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n300_), .B2(KEYINPUT21), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n255_), .B1(new_n283_), .B2(new_n303_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n295_), .A2(new_n296_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n305_));
  AOI211_X1 g104(.A(new_n254_), .B(new_n305_), .C1(new_n282_), .C2(KEYINPUT29), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G78gat), .B(G106gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(KEYINPUT95), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G22gat), .B(G50gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(KEYINPUT28), .Z(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n282_), .B2(KEYINPUT29), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n272_), .A2(new_n276_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT90), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n318_), .A2(new_n278_), .A3(new_n261_), .A4(new_n279_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n270_), .A4(new_n314_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n310_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n312_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n304_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n306_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n308_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT91), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n322_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n316_), .A2(KEYINPUT91), .A3(new_n321_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n309_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT94), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n307_), .A2(new_n308_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT94), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n334_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n325_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT20), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G190gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n211_), .B1(new_n216_), .B2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n207_), .A2(KEYINPUT96), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT96), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n203_), .B2(new_n206_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n344_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n210_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n232_), .A2(new_n349_), .A3(new_n223_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n342_), .B1(new_n351_), .B2(new_n303_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n234_), .B2(new_n303_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT19), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT97), .B(KEYINPUT18), .Z(new_n357_));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT20), .B1(new_n351_), .B2(new_n303_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n234_), .A2(new_n303_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n355_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n356_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n361_), .B1(new_n356_), .B2(new_n366_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n341_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n356_), .A2(new_n366_), .A3(new_n361_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n225_), .A2(new_n226_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n349_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT85), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n229_), .A3(new_n232_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n305_), .B1(new_n374_), .B2(new_n220_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n355_), .B1(new_n375_), .B2(new_n362_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n352_), .B(new_n365_), .C1(new_n234_), .C2(new_n303_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(KEYINPUT27), .B(new_n370_), .C1(new_n378_), .C2(new_n361_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n369_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT99), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n282_), .A2(KEYINPUT98), .A3(new_n242_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n242_), .A2(KEYINPUT98), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n242_), .A2(KEYINPUT98), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n319_), .A2(new_n384_), .A3(new_n385_), .A4(new_n270_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n382_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n383_), .A2(new_n386_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n242_), .A2(KEYINPUT4), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n388_), .A2(KEYINPUT4), .B1(new_n282_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n387_), .B1(new_n390_), .B2(new_n382_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G1gat), .B(G29gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT0), .ZN(new_n393_));
  INV_X1    g192(.A(G57gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G85gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n391_), .B(new_n396_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n340_), .A2(new_n380_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n361_), .A2(KEYINPUT32), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n356_), .A2(new_n366_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(new_n399_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n390_), .A2(new_n382_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n387_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(new_n396_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n391_), .A2(new_n396_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n402_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n367_), .A2(new_n368_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n382_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n390_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n396_), .B1(new_n388_), .B2(new_n382_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n409_), .B1(new_n405_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n408_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n340_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT100), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n398_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n338_), .B1(new_n337_), .B2(new_n334_), .ZN(new_n422_));
  AND4_X1   g221(.A1(new_n338_), .A2(new_n328_), .A3(new_n332_), .A4(new_n334_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n324_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n391_), .A2(new_n396_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n410_), .B(new_n411_), .C1(new_n425_), .C2(new_n409_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n426_), .B2(new_n408_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT100), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n251_), .B1(new_n421_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n397_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n424_), .A2(new_n380_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n251_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT8), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G99gat), .A2(G106gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(G85gat), .A2(G92gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G85gat), .A2(G92gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n434_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT65), .ZN(new_n448_));
  AND3_X1   g247(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n441_), .A2(KEYINPUT65), .A3(new_n442_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT66), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n438_), .A2(new_n451_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n444_), .A2(new_n445_), .A3(KEYINPUT8), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n438_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT66), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n447_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT64), .B(G85gat), .Z(new_n461_));
  INV_X1    g260(.A(G92gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n460_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n444_), .A2(KEYINPUT9), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n451_), .A2(new_n452_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT10), .B(G99gat), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n467_), .A2(G106gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT67), .B1(new_n459_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n443_), .A2(new_n446_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT8), .ZN(new_n473_));
  INV_X1    g272(.A(new_n458_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n454_), .A2(new_n455_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT67), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(new_n469_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G29gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n471_), .A2(new_n478_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT71), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G232gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT34), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n483_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n487_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n476_), .A2(new_n469_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n481_), .B(KEYINPUT15), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n493_), .A2(new_n489_), .A3(new_n482_), .A4(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n482_), .A2(new_n489_), .A3(new_n496_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G190gat), .B(G218gat), .Z(new_n501_));
  XNOR2_X1  g300(.A(G134gat), .B(G162gat), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n502_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT36), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n500_), .A2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT36), .B1(new_n503_), .B2(new_n504_), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT72), .Z(new_n509_));
  NAND3_X1  g308(.A1(new_n497_), .A2(new_n499_), .A3(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n433_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G57gat), .B(G64gat), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n513_), .A2(KEYINPUT11), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(KEYINPUT11), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G71gat), .B(G78gat), .ZN(new_n516_));
  OR3_X1    g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n516_), .A3(KEYINPUT11), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G15gat), .B(G22gat), .ZN(new_n520_));
  INV_X1    g319(.A(G1gat), .ZN(new_n521_));
  INV_X1    g320(.A(G8gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G8gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n519_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G183gat), .B(G211gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G127gat), .B(G155gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT76), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n530_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(KEYINPUT77), .Z(new_n540_));
  XOR2_X1   g339(.A(new_n535_), .B(KEYINPUT78), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT17), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n542_), .A2(new_n530_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(G230gat), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(new_n253_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n471_), .A2(new_n478_), .A3(new_n519_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT68), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n471_), .A2(new_n478_), .A3(KEYINPUT68), .A4(new_n519_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n519_), .B1(new_n471_), .B2(new_n478_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n546_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n546_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n547_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n519_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n459_), .A2(new_n470_), .A3(KEYINPUT67), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n477_), .B1(new_n476_), .B2(new_n469_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT12), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n494_), .A2(KEYINPUT12), .A3(new_n557_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n556_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G120gat), .B(G148gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT69), .B(G204gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT5), .B(G176gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  NAND3_X1  g368(.A1(new_n553_), .A2(new_n564_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n553_), .B2(new_n564_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(KEYINPUT13), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT13), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n526_), .B(new_n481_), .Z(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n495_), .A2(new_n526_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n527_), .A2(new_n481_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n583_), .A3(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT80), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT79), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n586_), .B(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n512_), .A2(new_n544_), .A3(new_n577_), .A4(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G1gat), .B1(new_n593_), .B2(new_n430_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT101), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n577_), .A2(new_n592_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n506_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT37), .B1(new_n598_), .B2(KEYINPUT73), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n511_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT73), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT37), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n507_), .B(new_n510_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n544_), .B1(new_n600_), .B2(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n433_), .A2(new_n596_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n521_), .A3(new_n397_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT38), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n595_), .A2(new_n608_), .ZN(G1324gat));
  AND2_X1   g408(.A1(new_n369_), .A2(new_n379_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G8gat), .B1(new_n593_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(KEYINPUT102), .A3(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n606_), .A2(new_n522_), .A3(new_n380_), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n615_));
  OAI211_X1 g414(.A(new_n613_), .B(new_n614_), .C1(new_n611_), .C2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT40), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(G1325gat));
  AND2_X1   g417(.A1(new_n247_), .A2(new_n250_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G15gat), .B1(new_n593_), .B2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT41), .Z(new_n621_));
  INV_X1    g420(.A(G15gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n606_), .A2(new_n622_), .A3(new_n251_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(G1326gat));
  OAI21_X1  g423(.A(G22gat), .B1(new_n593_), .B2(new_n340_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT42), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n340_), .A2(G22gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT103), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n606_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(G1327gat));
  INV_X1    g429(.A(new_n511_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n433_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n596_), .A2(new_n544_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n397_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n600_), .A2(new_n604_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n636_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT43), .B1(new_n637_), .B2(KEYINPUT105), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639_));
  INV_X1    g438(.A(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n610_), .A2(new_n424_), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n427_), .A2(KEYINPUT100), .B1(new_n397_), .B2(new_n641_), .ZN(new_n642_));
  AOI211_X1 g441(.A(new_n420_), .B(new_n424_), .C1(new_n408_), .C2(new_n426_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n619_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n251_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n640_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n639_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n638_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n639_), .B(KEYINPUT43), .C1(new_n646_), .C2(new_n647_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n649_), .A2(KEYINPUT44), .A3(new_n633_), .A4(new_n650_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n651_), .A2(G29gat), .A3(new_n397_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n649_), .A2(new_n633_), .A3(new_n650_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n635_), .B1(new_n652_), .B2(new_n655_), .ZN(G1328gat));
  NOR2_X1   g455(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n657_));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n651_), .A2(new_n380_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(new_n655_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n634_), .A2(new_n658_), .A3(new_n380_), .ZN(new_n661_));
  XOR2_X1   g460(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n661_), .B(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n657_), .B1(new_n660_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n655_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n651_), .A2(new_n380_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G36gat), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n657_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n661_), .B(new_n662_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n665_), .A2(new_n671_), .ZN(G1329gat));
  NAND2_X1  g471(.A1(new_n634_), .A2(new_n251_), .ZN(new_n673_));
  INV_X1    g472(.A(G43gat), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n651_), .A2(G43gat), .A3(new_n251_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n666_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n634_), .B2(new_n424_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n651_), .A2(G50gat), .A3(new_n424_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(new_n655_), .ZN(G1331gat));
  INV_X1    g480(.A(new_n592_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n576_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n512_), .A2(new_n544_), .A3(new_n684_), .ZN(new_n685_));
  OR3_X1    g484(.A1(new_n685_), .A2(new_n394_), .A3(new_n430_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n433_), .A2(new_n605_), .A3(new_n683_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n394_), .B1(new_n689_), .B2(new_n430_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n686_), .A2(new_n687_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n688_), .A2(KEYINPUT109), .A3(new_n690_), .A4(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1332gat));
  OAI21_X1  g495(.A(G64gat), .B1(new_n685_), .B2(new_n610_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT48), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n610_), .A2(G64gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n689_), .B2(new_n699_), .ZN(G1333gat));
  OR3_X1    g499(.A1(new_n689_), .A2(G71gat), .A3(new_n619_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G71gat), .B1(new_n685_), .B2(new_n619_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n702_), .A2(KEYINPUT110), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(KEYINPUT110), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(KEYINPUT49), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT49), .B1(new_n703_), .B2(new_n704_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n701_), .B1(new_n705_), .B2(new_n706_), .ZN(G1334gat));
  OAI21_X1  g506(.A(G78gat), .B1(new_n685_), .B2(new_n340_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT50), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n340_), .A2(G78gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n689_), .B2(new_n710_), .ZN(G1335gat));
  INV_X1    g510(.A(new_n544_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n576_), .A2(new_n712_), .A3(new_n682_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT111), .B1(new_n632_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n717_));
  NOR4_X1   g516(.A1(new_n433_), .A2(new_n717_), .A3(new_n713_), .A4(new_n631_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n397_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n713_), .B(KEYINPUT112), .Z(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT105), .B1(new_n637_), .B2(KEYINPUT104), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n646_), .B2(new_n639_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n650_), .B(new_n722_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT113), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n430_), .A2(new_n461_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n721_), .B1(new_n727_), .B2(new_n728_), .ZN(G1336gat));
  NAND3_X1  g528(.A1(new_n720_), .A2(new_n462_), .A3(new_n380_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n727_), .A2(new_n380_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(new_n462_), .ZN(G1337gat));
  OR2_X1    g531(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n619_), .A2(new_n467_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n715_), .B2(new_n718_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT114), .B(new_n734_), .C1(new_n715_), .C2(new_n718_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G99gat), .B1(new_n726_), .B2(new_n619_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n741_));
  AND4_X1   g540(.A1(new_n733_), .A2(new_n739_), .A3(new_n740_), .A4(new_n741_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n737_), .A2(new_n738_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n733_), .B1(new_n743_), .B2(new_n740_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1338gat));
  XNOR2_X1  g544(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n746_));
  OAI21_X1  g545(.A(G106gat), .B1(new_n726_), .B2(new_n340_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT52), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n749_), .B(G106gat), .C1(new_n726_), .C2(new_n340_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n340_), .A2(G106gat), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n746_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n746_), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n757_), .B(new_n754_), .C1(new_n748_), .C2(new_n750_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1339gat));
  INV_X1    g558(.A(KEYINPUT123), .ZN(new_n760_));
  AND2_X1   g559(.A1(KEYINPUT122), .A2(KEYINPUT57), .ZN(new_n761_));
  NOR2_X1   g560(.A1(KEYINPUT122), .A2(KEYINPUT57), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n570_), .A2(new_n592_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n563_), .B1(new_n552_), .B2(KEYINPUT12), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n546_), .B1(new_n551_), .B2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n556_), .A2(new_n562_), .A3(KEYINPUT55), .A4(new_n563_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n769_), .B1(new_n766_), .B2(new_n555_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n768_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n569_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n771_), .A2(KEYINPUT56), .A3(new_n772_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n765_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n578_), .A2(new_n579_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n582_), .A2(new_n583_), .A3(new_n580_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n590_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT119), .Z(new_n781_));
  NOR2_X1   g580(.A1(new_n585_), .A2(new_n590_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n631_), .B(new_n764_), .C1(new_n777_), .C2(new_n785_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n771_), .A2(KEYINPUT56), .A3(new_n772_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n772_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n570_), .B(new_n592_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n511_), .B1(new_n789_), .B2(new_n784_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n790_), .B2(new_n761_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n783_), .A2(new_n570_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT120), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT58), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n787_), .A2(new_n788_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT120), .B(new_n796_), .C1(new_n797_), .C2(new_n792_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n636_), .A2(new_n795_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n791_), .B1(KEYINPUT121), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT121), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n636_), .A2(new_n795_), .A3(new_n801_), .A4(new_n798_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n544_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n574_), .A2(new_n575_), .A3(new_n682_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  OAI22_X1  g604(.A1(new_n605_), .A2(new_n804_), .B1(new_n805_), .B2(KEYINPUT54), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(KEYINPUT54), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT118), .Z(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n806_), .B(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n760_), .B1(new_n803_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n799_), .A2(KEYINPUT121), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n790_), .A2(new_n761_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n812_), .A2(new_n802_), .A3(new_n786_), .A4(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n712_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n806_), .B(new_n808_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(KEYINPUT123), .A3(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n251_), .A2(new_n397_), .A3(new_n431_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n811_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT59), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n813_), .A2(new_n799_), .A3(new_n786_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n712_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n816_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT124), .B1(new_n592_), .B2(G113gat), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n820_), .A2(new_n826_), .A3(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G113gat), .B1(new_n829_), .B2(KEYINPUT124), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n811_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n592_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1340gat));
  NAND2_X1  g632(.A1(new_n820_), .A2(new_n826_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n577_), .B2(G120gat), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n576_), .B1(new_n819_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G120gat), .B1(new_n834_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n831_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1341gat));
  AOI21_X1  g640(.A(KEYINPUT125), .B1(new_n544_), .B2(G127gat), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n820_), .A2(new_n826_), .A3(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(G127gat), .B1(new_n844_), .B2(KEYINPUT125), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n544_), .A3(new_n831_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1342gat));
  INV_X1    g646(.A(G134gat), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n640_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n825_), .B(new_n850_), .C1(new_n819_), .C2(KEYINPUT59), .ZN(new_n851_));
  AOI21_X1  g650(.A(G134gat), .B1(new_n831_), .B2(new_n511_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT126), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n820_), .A2(new_n826_), .A3(new_n849_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT126), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n848_), .B1(new_n819_), .B2(new_n631_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(G1343gat));
  AND2_X1   g657(.A1(new_n811_), .A2(new_n817_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n251_), .A2(new_n430_), .A3(new_n641_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n592_), .A3(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n576_), .A3(new_n860_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n544_), .A3(new_n860_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  NAND2_X1  g666(.A1(new_n859_), .A2(new_n860_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G162gat), .B1(new_n868_), .B2(new_n640_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n631_), .A2(G162gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n868_), .B2(new_n870_), .ZN(G1347gat));
  AOI21_X1  g670(.A(new_n424_), .B1(new_n816_), .B2(new_n824_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n430_), .A2(new_n380_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n619_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G169gat), .B1(new_n875_), .B2(new_n682_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n875_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n222_), .A3(new_n592_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n877_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n880_), .A3(new_n881_), .ZN(G1348gat));
  AND2_X1   g681(.A1(new_n859_), .A2(new_n340_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n577_), .A2(new_n619_), .A3(new_n209_), .A4(new_n873_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n576_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n883_), .A2(new_n884_), .B1(new_n221_), .B2(new_n885_), .ZN(G1349gat));
  INV_X1    g685(.A(new_n216_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n619_), .A2(new_n712_), .A3(new_n873_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n872_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n883_), .A2(new_n888_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n214_), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n875_), .B2(new_n640_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n511_), .A2(new_n343_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n875_), .B2(new_n893_), .ZN(G1351gat));
  NOR3_X1   g693(.A1(new_n251_), .A2(new_n340_), .A3(new_n873_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n859_), .A2(new_n592_), .A3(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g696(.A1(new_n859_), .A2(new_n576_), .A3(new_n895_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT127), .B(G204gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1353gat));
  NAND3_X1  g699(.A1(new_n859_), .A2(new_n544_), .A3(new_n895_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT63), .B(G211gat), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n901_), .B2(new_n904_), .ZN(G1354gat));
  NAND2_X1  g704(.A1(new_n859_), .A2(new_n895_), .ZN(new_n906_));
  OAI21_X1  g705(.A(G218gat), .B1(new_n906_), .B2(new_n640_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n631_), .A2(G218gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n906_), .B2(new_n908_), .ZN(G1355gat));
endmodule


