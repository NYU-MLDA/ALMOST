//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_;
  INV_X1    g000(.A(G106gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(G228gat), .B1(KEYINPUT85), .B2(G233gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n203_), .B1(KEYINPUT85), .B2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT88), .A2(KEYINPUT21), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT87), .B(G204gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G197gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n207_), .B(new_n209_), .C1(G197gat), .C2(G204gat), .ZN(new_n210_));
  INV_X1    g009(.A(G197gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(G204gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n212_), .B(KEYINPUT86), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n211_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n213_), .A2(KEYINPUT21), .A3(new_n214_), .A4(new_n205_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT84), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n204_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G78gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT84), .B1(new_n210_), .B2(new_n215_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n221_), .A2(G78gat), .A3(new_n204_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n202_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n219_), .ZN(new_n224_));
  OAI21_X1  g023(.A(G78gat), .B1(new_n221_), .B2(new_n204_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(G106gat), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n216_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G141gat), .B(G148gat), .Z(new_n229_));
  NAND2_X1  g028(.A1(G155gat), .A2(G162gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT1), .ZN(new_n231_));
  OR2_X1    g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n230_), .A2(KEYINPUT1), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n229_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT82), .Z(new_n236_));
  NOR2_X1   g035(.A1(G141gat), .A2(G148gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT3), .Z(new_n238_));
  NAND2_X1  g037(.A1(G141gat), .A2(G148gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT2), .Z(new_n240_));
  OAI211_X1 g039(.A(new_n230_), .B(new_n232_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n228_), .B1(new_n242_), .B2(KEYINPUT29), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n227_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT83), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n223_), .A2(new_n243_), .A3(new_n226_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n242_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT29), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT28), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G22gat), .B(G50gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n252_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n245_), .A2(new_n246_), .A3(new_n255_), .A4(new_n247_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n253_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n254_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT25), .B(G183gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT26), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT75), .B1(new_n261_), .B2(G190gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G190gat), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n260_), .B(new_n262_), .C1(new_n263_), .C2(KEYINPUT75), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT76), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G176gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT24), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  MUX2_X1   g068(.A(new_n268_), .B(KEYINPUT24), .S(new_n269_), .Z(new_n270_));
  NAND2_X1  g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT23), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n265_), .A2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(G183gat), .B2(G190gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n275_), .A2(KEYINPUT78), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(new_n271_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(new_n278_), .B2(new_n271_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n280_), .A2(KEYINPUT78), .ZN(new_n281_));
  AOI21_X1  g080(.A(G176gat), .B1(KEYINPUT77), .B2(KEYINPUT22), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(new_n266_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n276_), .A2(new_n281_), .A3(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n274_), .A2(new_n284_), .ZN(new_n285_));
  OR3_X1    g084(.A1(new_n285_), .A2(KEYINPUT91), .A3(new_n228_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT91), .B1(new_n285_), .B2(new_n228_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT22), .B(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT89), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT90), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n291_), .A2(new_n267_), .B1(new_n275_), .B2(new_n292_), .ZN(new_n293_));
  OAI221_X1 g092(.A(new_n293_), .B1(new_n292_), .B2(new_n280_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n263_), .A2(new_n260_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n270_), .A2(new_n272_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT20), .B1(new_n297_), .B2(new_n216_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT19), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n288_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT20), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n297_), .B2(new_n216_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n285_), .A2(new_n228_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G8gat), .B(G36gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT18), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G64gat), .B(G92gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n298_), .B1(new_n287_), .B2(new_n286_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n307_), .B1(new_n316_), .B2(new_n302_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT27), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n317_), .B2(new_n313_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n305_), .A2(new_n302_), .A3(new_n306_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(new_n316_), .B2(new_n302_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n314_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n319_), .A2(new_n320_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G71gat), .B(G99gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(G43gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(G15gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n327_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT30), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n285_), .B(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n334_), .A2(KEYINPUT79), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(KEYINPUT79), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n332_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n331_), .B1(new_n334_), .B2(KEYINPUT79), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G127gat), .B(G134gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n340_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(KEYINPUT80), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n339_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n337_), .A2(new_n338_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G1gat), .B(G29gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G85gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT0), .B(G57gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n242_), .A2(new_n346_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n341_), .A2(new_n342_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n236_), .A2(new_n241_), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n360_), .A2(KEYINPUT92), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(KEYINPUT92), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n356_), .A2(new_n364_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n357_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n355_), .B1(new_n363_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n367_), .ZN(new_n370_));
  OAI211_X1 g169(.A(G225gat), .B(G233gat), .C1(new_n370_), .C2(new_n365_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n371_), .A2(new_n354_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n349_), .A2(new_n350_), .A3(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n259_), .A2(new_n325_), .A3(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n313_), .A2(KEYINPUT32), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n323_), .A2(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n373_), .B(new_n377_), .C1(new_n309_), .C2(new_n376_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n363_), .A2(new_n368_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n379_), .A2(KEYINPUT93), .A3(KEYINPUT33), .A4(new_n354_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT93), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n372_), .B2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n372_), .A2(new_n382_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n356_), .A2(new_n359_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n355_), .B1(new_n386_), .B2(new_n357_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n387_), .A2(KEYINPUT94), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(KEYINPUT94), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n357_), .B1(new_n370_), .B2(new_n365_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n315_), .A2(new_n318_), .A3(new_n385_), .A4(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n378_), .B1(new_n384_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n259_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n373_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n325_), .B(new_n395_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n349_), .A2(new_n350_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n375_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G99gat), .A2(G106gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT6), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(G99gat), .A3(G106gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT10), .B(G99gat), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n405_), .B1(new_n406_), .B2(G106gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT64), .ZN(new_n408_));
  OAI211_X1 g207(.A(G85gat), .B(G92gat), .C1(new_n408_), .C2(KEYINPUT9), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n408_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n409_), .A2(new_n410_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n407_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G85gat), .B(G92gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n402_), .A2(new_n404_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT7), .ZN(new_n417_));
  INV_X1    g216(.A(G99gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n202_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n415_), .B1(new_n416_), .B2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n403_), .B1(G99gat), .B2(G106gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n401_), .A2(KEYINPUT6), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n420_), .B(new_n419_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n423_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n415_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n413_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G29gat), .B(G36gat), .Z(new_n433_));
  XOR2_X1   g232(.A(G43gat), .B(G50gat), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n420_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AOI211_X1 g238(.A(new_n423_), .B(new_n414_), .C1(new_n439_), .C2(new_n405_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n428_), .B1(new_n427_), .B2(new_n415_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n431_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n413_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n435_), .B(KEYINPUT15), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n436_), .A2(KEYINPUT69), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n435_), .ZN(new_n447_));
  OR3_X1    g246(.A1(new_n444_), .A2(KEYINPUT69), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT35), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G190gat), .B(G218gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT71), .ZN(new_n452_));
  XOR2_X1   g251(.A(G134gat), .B(G162gat), .Z(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n449_), .A2(new_n450_), .B1(KEYINPUT36), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G232gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT35), .ZN(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n458_));
  XOR2_X1   g257(.A(new_n457_), .B(new_n458_), .Z(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(new_n449_), .B2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n446_), .A2(KEYINPUT70), .A3(new_n448_), .A4(new_n459_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n455_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n454_), .A2(KEYINPUT36), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n455_), .A2(new_n462_), .A3(new_n467_), .A4(new_n463_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n400_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G230gat), .ZN(new_n472_));
  INV_X1    g271(.A(G233gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G64gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n476_));
  XOR2_X1   g275(.A(G71gat), .B(G78gat), .Z(new_n477_));
  OR2_X1    g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n477_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n474_), .B1(new_n432_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n483_));
  INV_X1    g282(.A(new_n481_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n444_), .B2(new_n484_), .ZN(new_n485_));
  AOI211_X1 g284(.A(KEYINPUT12), .B(new_n481_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n482_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n432_), .A2(new_n481_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n424_), .A2(new_n429_), .B1(KEYINPUT65), .B2(KEYINPUT8), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n484_), .B1(new_n490_), .B2(new_n413_), .ZN(new_n491_));
  AOI211_X1 g290(.A(new_n472_), .B(new_n473_), .C1(new_n489_), .C2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G120gat), .B(G148gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(G176gat), .B(G204gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT66), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT66), .B(new_n498_), .C1(new_n488_), .C2(new_n492_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n500_), .A2(KEYINPUT13), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT13), .B1(new_n500_), .B2(new_n501_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(G231gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n481_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G1gat), .B(G8gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT72), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(G22gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n329_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G15gat), .A2(G22gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G1gat), .A2(G8gat), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n512_), .A2(new_n513_), .B1(KEYINPUT14), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n510_), .B(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n507_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n507_), .A2(new_n516_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G127gat), .B(G155gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT16), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G183gat), .B(G211gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n523_), .A2(new_n524_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n517_), .A2(new_n528_), .A3(new_n518_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n510_), .A2(new_n515_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n510_), .A2(new_n515_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n447_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n516_), .A2(new_n435_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT74), .ZN(new_n536_));
  OR3_X1    g335(.A1(new_n516_), .A2(KEYINPUT74), .A3(new_n435_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n536_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n445_), .A2(new_n533_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(new_n535_), .A3(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G169gat), .B(G197gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n540_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n505_), .A2(new_n530_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n471_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT95), .ZN(new_n554_));
  OAI21_X1  g353(.A(G1gat), .B1(new_n554_), .B2(new_n395_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n400_), .A2(new_n551_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n529_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n525_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT73), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT73), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n527_), .A2(new_n560_), .A3(new_n529_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT37), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n469_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n466_), .A2(KEYINPUT37), .A3(new_n468_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n556_), .A2(new_n504_), .A3(new_n563_), .A4(new_n568_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n569_), .A2(G1gat), .A3(new_n395_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n570_), .A2(KEYINPUT38), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(KEYINPUT38), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n555_), .A2(new_n571_), .A3(new_n572_), .ZN(G1324gat));
  OAI21_X1  g372(.A(G8gat), .B1(new_n553_), .B2(new_n325_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT39), .ZN(new_n575_));
  OR3_X1    g374(.A1(new_n569_), .A2(G8gat), .A3(new_n325_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g377(.A(G15gat), .B1(new_n554_), .B2(new_n399_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT41), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT41), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n569_), .A2(G15gat), .A3(new_n399_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT96), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n581_), .A3(new_n583_), .ZN(G1326gat));
  OAI21_X1  g383(.A(G22gat), .B1(new_n554_), .B2(new_n259_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT42), .ZN(new_n586_));
  INV_X1    g385(.A(new_n259_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n511_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n586_), .B1(new_n569_), .B2(new_n588_), .ZN(G1327gat));
  NOR2_X1   g388(.A1(new_n469_), .A2(new_n563_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT101), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(new_n505_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n556_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT102), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT102), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n556_), .A2(new_n595_), .A3(new_n592_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(G29gat), .B1(new_n597_), .B2(new_n373_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n504_), .A2(new_n550_), .A3(new_n562_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT97), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT43), .B1(new_n568_), .B2(KEYINPUT98), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n400_), .B2(new_n568_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n398_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n567_), .B(new_n601_), .C1(new_n604_), .C2(new_n375_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n600_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT99), .B1(new_n606_), .B2(KEYINPUT44), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n605_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n600_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT44), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n375_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n258_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n253_), .A2(new_n256_), .A3(new_n254_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n373_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n617_), .A2(new_n325_), .B1(new_n393_), .B2(new_n259_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n614_), .B1(new_n618_), .B2(new_n398_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n601_), .B1(new_n619_), .B2(new_n567_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n605_), .ZN(new_n621_));
  OAI211_X1 g420(.A(KEYINPUT44), .B(new_n609_), .C1(new_n620_), .C2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n606_), .A2(KEYINPUT100), .A3(KEYINPUT44), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n607_), .A2(new_n613_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n373_), .A2(G29gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n598_), .B1(new_n626_), .B2(new_n627_), .ZN(G1328gat));
  INV_X1    g427(.A(KEYINPUT46), .ZN(new_n629_));
  INV_X1    g428(.A(G36gat), .ZN(new_n630_));
  INV_X1    g429(.A(new_n325_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n626_), .B2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n594_), .A2(new_n630_), .A3(new_n631_), .A4(new_n596_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT45), .Z(new_n634_));
  OAI21_X1  g433(.A(new_n629_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n613_), .A2(new_n607_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n624_), .A2(new_n625_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n631_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G36gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n633_), .B(KEYINPUT45), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(KEYINPUT46), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n635_), .A2(new_n641_), .ZN(G1329gat));
  NAND4_X1  g441(.A1(new_n636_), .A2(new_n637_), .A3(G43gat), .A4(new_n398_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n597_), .A2(new_n398_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT103), .B(G43gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT47), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT47), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n643_), .A2(new_n649_), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(G1330gat));
  INV_X1    g450(.A(G50gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n626_), .B2(new_n587_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n597_), .A2(new_n652_), .A3(new_n587_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT104), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n636_), .A2(new_n637_), .A3(new_n587_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(G50gat), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(new_n654_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n656_), .A2(new_n660_), .ZN(G1331gat));
  NOR2_X1   g460(.A1(new_n400_), .A2(new_n550_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n662_), .A2(new_n505_), .A3(new_n563_), .A4(new_n568_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n395_), .B1(new_n663_), .B2(KEYINPUT105), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n664_), .B1(KEYINPUT105), .B2(new_n663_), .ZN(new_n665_));
  INV_X1    g464(.A(G57gat), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n559_), .A2(new_n561_), .A3(new_n548_), .A4(new_n549_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n504_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n471_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n666_), .B1(new_n373_), .B2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n671_), .B2(new_n666_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n665_), .A2(new_n666_), .B1(new_n670_), .B2(new_n673_), .ZN(G1332gat));
  OAI21_X1  g473(.A(G64gat), .B1(new_n669_), .B2(new_n325_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT48), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n325_), .A2(G64gat), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT107), .Z(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n663_), .B2(new_n678_), .ZN(G1333gat));
  OAI21_X1  g478(.A(G71gat), .B1(new_n669_), .B2(new_n399_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n399_), .A2(G71gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n663_), .B2(new_n683_), .ZN(G1334gat));
  OAI21_X1  g483(.A(G78gat), .B1(new_n669_), .B2(new_n259_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT50), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n587_), .A2(new_n219_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n663_), .B2(new_n687_), .ZN(G1335gat));
  NOR3_X1   g487(.A1(new_n504_), .A2(new_n550_), .A3(new_n563_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G85gat), .B1(new_n692_), .B2(new_n395_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n591_), .A2(new_n504_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n662_), .A2(new_n694_), .ZN(new_n695_));
  OR3_X1    g494(.A1(new_n695_), .A2(G85gat), .A3(new_n395_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1336gat));
  OAI21_X1  g496(.A(G92gat), .B1(new_n692_), .B2(new_n325_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n695_), .ZN(new_n699_));
  INV_X1    g498(.A(G92gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n631_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT109), .Z(G1337gat));
  NOR3_X1   g502(.A1(new_n695_), .A2(new_n399_), .A3(new_n406_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(KEYINPUT51), .ZN(new_n706_));
  OAI21_X1  g505(.A(G99gat), .B1(new_n692_), .B2(new_n399_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n705_), .A2(KEYINPUT51), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n708_), .B(new_n709_), .Z(G1338gat));
  NAND3_X1  g509(.A1(new_n699_), .A2(new_n202_), .A3(new_n587_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT111), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n608_), .A2(KEYINPUT112), .A3(new_n587_), .A4(new_n689_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(G106gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT112), .B1(new_n691_), .B2(new_n587_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n714_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n715_), .A2(G106gat), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(new_n717_), .A3(new_n713_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n712_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT53), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT53), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n712_), .B(new_n724_), .C1(new_n719_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1339gat));
  NOR2_X1   g525(.A1(new_n399_), .A2(new_n395_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(new_n259_), .A3(new_n325_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(KEYINPUT59), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT55), .B(new_n482_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT116), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n491_), .A2(KEYINPUT12), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n444_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT116), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(KEYINPUT55), .A4(new_n482_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n731_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT117), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n489_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n740_));
  AOI22_X1  g539(.A1(new_n739_), .A2(new_n487_), .B1(new_n740_), .B2(new_n474_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n737_), .A2(new_n738_), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n738_), .B1(new_n737_), .B2(new_n741_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n498_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT56), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(KEYINPUT120), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n538_), .B1(new_n516_), .B2(new_n435_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n546_), .B1(new_n541_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n549_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT119), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n488_), .A2(new_n492_), .A3(new_n498_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n498_), .B(new_n757_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n747_), .A2(new_n756_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT58), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n747_), .A2(new_n756_), .A3(KEYINPUT58), .A4(new_n758_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(new_n567_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT115), .B1(new_n551_), .B2(new_n754_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n755_), .A2(new_n550_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(KEYINPUT56), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n744_), .A2(new_n769_), .ZN(new_n770_));
  OAI221_X1 g569(.A(new_n498_), .B1(new_n768_), .B2(KEYINPUT56), .C1(new_n742_), .C2(new_n743_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n500_), .A2(new_n501_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n753_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n469_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n761_), .A2(new_n763_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT57), .B(new_n469_), .C1(new_n772_), .C2(new_n774_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n563_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n667_), .A2(KEYINPUT114), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n551_), .A2(new_n782_), .A3(new_n559_), .A4(new_n561_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n505_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n780_), .B1(new_n568_), .B2(new_n785_), .ZN(new_n786_));
  NOR4_X1   g585(.A1(new_n567_), .A2(new_n505_), .A3(KEYINPUT54), .A4(new_n784_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT122), .B(new_n729_), .C1(new_n779_), .C2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT122), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n775_), .A2(new_n776_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n761_), .A2(new_n567_), .A3(new_n762_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n778_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n788_), .B1(new_n793_), .B2(new_n562_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n729_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n790_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n789_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n793_), .A2(new_n530_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n788_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n728_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G113gat), .B1(new_n802_), .B2(new_n551_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n728_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n530_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n806_), .B2(new_n788_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT121), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n551_), .A2(G113gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n803_), .B1(new_n808_), .B2(new_n809_), .ZN(G1340gat));
  AOI21_X1  g609(.A(new_n504_), .B1(new_n807_), .B2(KEYINPUT59), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n811_), .A2(new_n797_), .A3(KEYINPUT123), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT123), .B1(new_n811_), .B2(new_n797_), .ZN(new_n813_));
  INV_X1    g612(.A(G120gat), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n812_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n504_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(KEYINPUT60), .B2(new_n814_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n808_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT124), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n818_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n811_), .A2(new_n797_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT123), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G120gat), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n820_), .B(new_n821_), .C1(new_n825_), .C2(new_n812_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n819_), .A2(new_n826_), .ZN(G1341gat));
  OAI21_X1  g626(.A(G127gat), .B1(new_n802_), .B2(new_n530_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n562_), .A2(G127gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n808_), .B2(new_n829_), .ZN(G1342gat));
  OAI21_X1  g629(.A(G134gat), .B1(new_n802_), .B2(new_n568_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n469_), .A2(G134gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n808_), .B2(new_n832_), .ZN(G1343gat));
  NAND2_X1  g632(.A1(new_n799_), .A2(new_n800_), .ZN(new_n834_));
  NOR4_X1   g633(.A1(new_n259_), .A2(new_n631_), .A3(new_n395_), .A4(new_n398_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n550_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n505_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g640(.A1(new_n836_), .A2(new_n562_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT61), .B(G155gat), .Z(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1346gat));
  INV_X1    g643(.A(G162gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n836_), .B2(new_n469_), .ZN(new_n846_));
  XOR2_X1   g645(.A(new_n846_), .B(KEYINPUT125), .Z(new_n847_));
  NOR3_X1   g646(.A1(new_n836_), .A2(new_n845_), .A3(new_n568_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1347gat));
  NAND2_X1  g648(.A1(new_n631_), .A2(new_n374_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n794_), .A2(new_n587_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G169gat), .B1(new_n852_), .B2(new_n551_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(KEYINPUT62), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n853_), .A2(KEYINPUT62), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n291_), .A3(new_n550_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(G1348gat));
  AOI21_X1  g656(.A(G176gat), .B1(new_n851_), .B2(new_n505_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n587_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n850_), .A2(new_n267_), .A3(new_n504_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(G1349gat));
  NAND4_X1  g660(.A1(new_n859_), .A2(new_n631_), .A3(new_n374_), .A4(new_n563_), .ZN(new_n862_));
  INV_X1    g661(.A(G183gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n530_), .A2(new_n260_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n862_), .A2(new_n863_), .B1(new_n851_), .B2(new_n864_), .ZN(G1350gat));
  OAI21_X1  g664(.A(G190gat), .B1(new_n852_), .B2(new_n568_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n851_), .A2(new_n263_), .A3(new_n470_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1351gat));
  AND4_X1   g667(.A1(new_n617_), .A2(new_n834_), .A3(new_n631_), .A4(new_n399_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n550_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g670(.A1(new_n869_), .A2(new_n505_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(G204gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n208_), .B2(new_n872_), .ZN(G1353gat));
  NAND2_X1  g673(.A1(new_n869_), .A2(new_n805_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n876_));
  AND2_X1   g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n875_), .A2(new_n876_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n879_), .A2(KEYINPUT126), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(KEYINPUT126), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n878_), .B1(new_n880_), .B2(new_n881_), .ZN(G1354gat));
  AOI21_X1  g681(.A(G218gat), .B1(new_n869_), .B2(new_n470_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n567_), .A2(G218gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT127), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n869_), .B2(new_n885_), .ZN(G1355gat));
endmodule


