//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_;
  AND2_X1   g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT9), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT9), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  INV_X1    g005(.A(G92gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(KEYINPUT64), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n202_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT10), .B(G99gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n209_), .A2(KEYINPUT65), .A3(new_n211_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n214_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G57gat), .B(G64gat), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n225_), .A2(KEYINPUT11), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(KEYINPUT11), .ZN(new_n227_));
  XOR2_X1   g026(.A(G71gat), .B(G78gat), .Z(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n227_), .A2(new_n228_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n221_), .A2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n236_));
  INV_X1    g035(.A(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(G106gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n219_), .A2(KEYINPUT67), .A3(new_n220_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n234_), .A2(new_n235_), .A3(new_n239_), .A4(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n202_), .A2(new_n203_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n232_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n239_), .A2(new_n219_), .A3(new_n235_), .A4(new_n220_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(new_n232_), .A3(new_n242_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT66), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n244_), .A2(new_n247_), .A3(new_n232_), .A4(new_n242_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n224_), .B(new_n231_), .C1(new_n243_), .C2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G230gat), .A2(G233gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n224_), .B1(new_n243_), .B2(new_n249_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n231_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(KEYINPUT12), .A3(new_n256_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n250_), .A2(KEYINPUT69), .A3(new_n251_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n254_), .A2(new_n259_), .A3(new_n260_), .A4(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT70), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n250_), .A2(KEYINPUT69), .A3(new_n251_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT69), .B1(new_n250_), .B2(new_n251_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n255_), .A2(KEYINPUT12), .A3(new_n256_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT12), .B1(new_n255_), .B2(new_n256_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n266_), .A2(new_n267_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n257_), .A2(new_n273_), .A3(new_n250_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n251_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n255_), .A2(KEYINPUT68), .A3(new_n256_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n272_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G120gat), .B(G148gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT5), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(G176gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT13), .ZN(new_n285_));
  INV_X1    g084(.A(new_n283_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n272_), .A2(new_n278_), .A3(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(new_n272_), .B2(new_n278_), .ZN(new_n289_));
  AOI211_X1 g088(.A(new_n277_), .B(new_n283_), .C1(new_n263_), .C2(new_n271_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT13), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G1gat), .B(G29gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G57gat), .B(G85gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G225gat), .A2(G233gat), .ZN(new_n299_));
  AND2_X1   g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n300_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G113gat), .B(G120gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n305_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT89), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n317_), .A2(G141gat), .A3(G148gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT89), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT2), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n317_), .A2(new_n320_), .B1(G141gat), .B2(G148gat), .ZN(new_n321_));
  NOR3_X1   g120(.A1(new_n315_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n302_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n308_), .B(new_n313_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n308_), .ZN(new_n325_));
  OR3_X1    g124(.A1(new_n315_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(new_n302_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n311_), .A2(KEYINPUT86), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n312_), .A2(KEYINPUT85), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n312_), .A2(KEYINPUT85), .ZN(new_n330_));
  OR3_X1    g129(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT86), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .A4(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n324_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT4), .ZN(new_n334_));
  AND4_X1   g133(.A1(new_n330_), .A2(new_n328_), .A3(new_n329_), .A4(new_n331_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n308_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n299_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(new_n299_), .A3(new_n324_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n298_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT4), .B1(new_n335_), .B2(new_n336_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(KEYINPUT4), .B2(new_n333_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n341_), .B(new_n297_), .C1(new_n345_), .C2(new_n299_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G183gat), .ZN(new_n348_));
  INV_X1    g147(.A(G190gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT23), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT83), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(G183gat), .A3(G190gat), .ZN(new_n354_));
  OAI211_X1 g153(.A(KEYINPUT83), .B(KEYINPUT23), .C1(new_n348_), .C2(new_n349_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(G183gat), .B2(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(G176gat), .ZN(new_n359_));
  OR2_X1    g158(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n362_), .A2(KEYINPUT95), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT95), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n359_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n357_), .A2(new_n358_), .A3(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n350_), .A2(new_n354_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT25), .B(G183gat), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT26), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G190gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n370_), .A2(G190gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n368_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G169gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n359_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n378_), .A2(KEYINPUT24), .A3(new_n358_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(KEYINPUT24), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n367_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G197gat), .B(G204gat), .Z(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT21), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G197gat), .B(G204gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT21), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G211gat), .ZN(new_n389_));
  INV_X1    g188(.A(G218gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G211gat), .A2(G218gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT92), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT92), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n395_), .A3(new_n392_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n385_), .A2(new_n388_), .A3(new_n394_), .A4(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n399_));
  OAI211_X1 g198(.A(KEYINPUT21), .B(new_n384_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n383_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT19), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n397_), .A2(new_n400_), .ZN(new_n406_));
  XOR2_X1   g205(.A(KEYINPUT81), .B(G190gat), .Z(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT26), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n373_), .A2(new_n408_), .A3(KEYINPUT82), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT81), .B(G190gat), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n411_), .A2(new_n370_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n410_), .B1(new_n412_), .B2(new_n372_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n409_), .A2(new_n413_), .A3(new_n356_), .A4(new_n381_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n359_), .B1(new_n415_), .B2(KEYINPUT22), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G169gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n362_), .A2(new_n415_), .A3(new_n359_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n411_), .A2(G183gat), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n417_), .B(new_n418_), .C1(new_n368_), .C2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n406_), .A2(new_n414_), .A3(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n402_), .A2(KEYINPUT20), .A3(new_n405_), .A4(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT98), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n414_), .A2(new_n420_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n425_), .B2(new_n401_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n406_), .A2(new_n367_), .A3(new_n382_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n404_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n421_), .A2(KEYINPUT20), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT98), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n405_), .A4(new_n402_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n423_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT18), .B(G64gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G92gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G8gat), .B(G36gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  AND2_X1   g236(.A1(new_n437_), .A2(KEYINPUT32), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n421_), .A2(KEYINPUT20), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n406_), .B1(new_n367_), .B2(new_n382_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n404_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n426_), .A2(new_n405_), .A3(new_n427_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT96), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT96), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n426_), .A2(new_n445_), .A3(new_n405_), .A4(new_n427_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n347_), .B(new_n439_), .C1(new_n448_), .C2(new_n438_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n437_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n437_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n444_), .A2(new_n451_), .A3(new_n446_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n299_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n337_), .A2(new_n453_), .A3(new_n324_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n298_), .B(new_n454_), .C1(new_n345_), .C2(new_n453_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n346_), .B(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n449_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G78gat), .B(G106gat), .Z(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n401_), .B1(new_n327_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(G228gat), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n406_), .B1(KEYINPUT29), .B2(new_n336_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(new_n467_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n461_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT93), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n463_), .A2(new_n468_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n467_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n460_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G22gat), .B(G50gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n327_), .A2(new_n462_), .A3(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n478_), .B1(new_n336_), .B2(KEYINPUT29), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(KEYINPUT93), .B(new_n461_), .C1(new_n469_), .C2(new_n471_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n477_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n472_), .A2(new_n485_), .A3(new_n476_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT94), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n472_), .A2(new_n485_), .A3(KEYINPUT94), .A4(new_n476_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n488_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n459_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n450_), .A2(KEYINPUT99), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT27), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n496_), .B1(new_n433_), .B2(new_n451_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n451_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT99), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n347_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n488_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n452_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n496_), .B1(new_n504_), .B2(new_n498_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n494_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G227gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(G15gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(G43gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G71gat), .B(G99gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n414_), .A2(new_n515_), .A3(new_n420_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n514_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n518_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n520_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n512_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n513_), .B1(new_n520_), .B2(new_n516_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n511_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n522_), .A2(KEYINPUT87), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT88), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT88), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n522_), .A2(KEYINPUT87), .A3(new_n528_), .A4(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n522_), .A2(new_n525_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n332_), .B(KEYINPUT31), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n527_), .A2(new_n533_), .A3(new_n534_), .A4(new_n529_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n501_), .A2(new_n493_), .A3(new_n505_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n347_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n507_), .A2(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G169gat), .B(G197gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(G141gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT79), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(G113gat), .ZN(new_n546_));
  AND2_X1   g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G29gat), .B(G36gat), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(G43gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(G43gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(G50gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(G50gat), .A3(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT76), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G15gat), .B(G22gat), .ZN(new_n558_));
  INV_X1    g357(.A(G1gat), .ZN(new_n559_));
  INV_X1    g358(.A(G8gat), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT14), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G1gat), .B(G8gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT76), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n557_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n565_), .B1(new_n557_), .B2(new_n566_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n547_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n547_), .B(KEYINPUT77), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT15), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n549_), .A2(G50gat), .A3(new_n550_), .ZN(new_n573_));
  AOI21_X1  g372(.A(G50gat), .B1(new_n549_), .B2(new_n550_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT15), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n567_), .B(new_n571_), .C1(new_n578_), .C2(new_n565_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n570_), .A2(KEYINPUT78), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT80), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n546_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n570_), .A2(new_n579_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT78), .B1(new_n546_), .B2(new_n581_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT100), .B1(new_n542_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT34), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT35), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n255_), .A2(new_n555_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n255_), .A2(new_n577_), .A3(KEYINPUT71), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT71), .B1(new_n255_), .B2(new_n577_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n592_), .B(new_n594_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n590_), .A2(new_n591_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n255_), .A2(new_n577_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT71), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n593_), .B1(new_n603_), .B2(new_n595_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n599_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n592_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(G134gat), .ZN(new_n609_));
  INV_X1    g408(.A(G162gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n600_), .A2(new_n606_), .A3(new_n607_), .A4(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(KEYINPUT36), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n600_), .B2(new_n606_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT72), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  AOI211_X1 g416(.A(KEYINPUT72), .B(new_n614_), .C1(new_n600_), .C2(new_n606_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT37), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n598_), .A2(new_n599_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n605_), .B1(new_n604_), .B2(new_n592_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT73), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT73), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n600_), .A2(new_n606_), .A3(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(new_n613_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT37), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n612_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n619_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G231gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n564_), .B(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(new_n231_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT16), .B(G183gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(new_n389_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT17), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n637_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n632_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n632_), .B(KEYINPUT74), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n638_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT75), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT75), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n629_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n540_), .A2(new_n541_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT27), .B1(new_n450_), .B2(new_n452_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n498_), .A2(new_n499_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT99), .B(new_n451_), .C1(new_n444_), .C2(new_n446_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n651_), .B1(new_n654_), .B2(new_n497_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n493_), .A2(new_n347_), .ZN(new_n656_));
  AOI22_X1  g455(.A1(new_n655_), .A2(new_n656_), .B1(new_n459_), .B2(new_n493_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n650_), .B1(new_n657_), .B2(new_n538_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659_));
  INV_X1    g458(.A(new_n586_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  AND4_X1   g460(.A1(new_n292_), .A2(new_n587_), .A3(new_n649_), .A4(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n559_), .A3(new_n347_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT38), .Z(new_n664_));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n658_), .A2(new_n292_), .A3(new_n660_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n625_), .A2(new_n612_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n648_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n670_), .A2(KEYINPUT101), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(KEYINPUT101), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n559_), .B1(new_n673_), .B2(new_n347_), .ZN(new_n674_));
  OR3_X1    g473(.A1(new_n664_), .A2(new_n665_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n665_), .B1(new_n664_), .B2(new_n674_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1324gat));
  INV_X1    g476(.A(new_n655_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n560_), .B1(new_n670_), .B2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n662_), .A2(new_n560_), .A3(new_n678_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT40), .ZN(G1325gat));
  NAND3_X1  g484(.A1(new_n662_), .A2(new_n509_), .A3(new_n538_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT104), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n673_), .A2(new_n538_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n688_), .B2(G15gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(G1326gat));
  AOI21_X1  g490(.A(new_n493_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n692_));
  INV_X1    g491(.A(G22gat), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n692_), .A2(KEYINPUT105), .A3(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT105), .B1(new_n692_), .B2(new_n693_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n662_), .A2(new_n693_), .A3(new_n503_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n694_), .A2(KEYINPUT42), .A3(new_n695_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(G1327gat));
  AND2_X1   g500(.A1(new_n648_), .A2(new_n667_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n587_), .A2(new_n661_), .A3(new_n292_), .A4(new_n702_), .ZN(new_n703_));
  OR3_X1    g502(.A1(new_n703_), .A2(G29gat), .A3(new_n502_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n542_), .B2(new_n628_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n658_), .A2(new_n706_), .A3(new_n629_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n292_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n709_), .A2(new_n647_), .A3(new_n586_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n708_), .A2(KEYINPUT44), .A3(new_n710_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n347_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n716_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT106), .B1(new_n716_), .B2(G29gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n704_), .B1(new_n717_), .B2(new_n718_), .ZN(G1328gat));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n703_), .A2(G36gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n678_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n723_));
  NOR4_X1   g522(.A1(new_n703_), .A2(KEYINPUT107), .A3(G36gat), .A4(new_n655_), .ZN(new_n724_));
  OR3_X1    g523(.A1(new_n722_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n723_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n713_), .A2(new_n678_), .A3(new_n714_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G36gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n726_), .A3(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n725_), .A2(new_n726_), .A3(KEYINPUT46), .A4(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1329gat));
  XOR2_X1   g532(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(G43gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n703_), .B2(new_n539_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(KEYINPUT108), .B(new_n736_), .C1(new_n703_), .C2(new_n539_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n713_), .A2(G43gat), .A3(new_n538_), .A4(new_n714_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n742_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n735_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n746_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(new_n734_), .A3(new_n744_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1330gat));
  NOR2_X1   g549(.A1(new_n493_), .A2(new_n552_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n703_), .A2(new_n493_), .ZN(new_n752_));
  AOI22_X1  g551(.A1(new_n715_), .A2(new_n751_), .B1(new_n552_), .B2(new_n752_), .ZN(G1331gat));
  NAND2_X1  g552(.A1(new_n649_), .A2(new_n709_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n658_), .B1(new_n754_), .B2(KEYINPUT111), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n660_), .B(new_n755_), .C1(KEYINPUT111), .C2(new_n754_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G57gat), .B1(new_n756_), .B2(new_n347_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n542_), .A2(new_n292_), .A3(new_n660_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n668_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(new_n502_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n757_), .B1(G57gat), .B2(new_n760_), .ZN(G1332gat));
  INV_X1    g560(.A(G64gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n756_), .A2(new_n762_), .A3(new_n678_), .ZN(new_n763_));
  OAI21_X1  g562(.A(G64gat), .B1(new_n759_), .B2(new_n655_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT48), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n756_), .A2(new_n767_), .A3(new_n538_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G71gat), .B1(new_n759_), .B2(new_n539_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT49), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1334gat));
  NOR2_X1   g570(.A1(new_n493_), .A2(G78gat), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT112), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n756_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G78gat), .B1(new_n759_), .B2(new_n493_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT50), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1335gat));
  AND2_X1   g576(.A1(new_n758_), .A2(new_n702_), .ZN(new_n778_));
  AOI21_X1  g577(.A(G85gat), .B1(new_n778_), .B2(new_n347_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n292_), .A2(new_n647_), .A3(new_n660_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n708_), .A2(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n347_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n779_), .B1(new_n782_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g582(.A(G92gat), .B1(new_n778_), .B2(new_n678_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n655_), .A2(new_n207_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n781_), .B2(new_n785_), .ZN(G1337gat));
  AOI21_X1  g585(.A(new_n237_), .B1(new_n781_), .B2(new_n538_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n539_), .A2(new_n215_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n778_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1338gat));
  NOR3_X1   g590(.A1(new_n542_), .A2(KEYINPUT43), .A3(new_n628_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n706_), .B1(new_n658_), .B2(new_n629_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n503_), .B(new_n780_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT114), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n708_), .A2(new_n796_), .A3(new_n503_), .A4(new_n780_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(G106gat), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT115), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n795_), .A2(new_n800_), .A3(G106gat), .A4(new_n797_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(KEYINPUT52), .A3(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n778_), .A2(new_n238_), .A3(new_n503_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n798_), .A2(KEYINPUT115), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT53), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n802_), .A2(new_n808_), .A3(new_n803_), .A4(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(G1339gat));
  AOI21_X1  g609(.A(KEYINPUT55), .B1(new_n263_), .B2(new_n271_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n259_), .A2(new_n260_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n250_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n275_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n262_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n283_), .B1(new_n811_), .B2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n290_), .B1(new_n817_), .B2(KEYINPUT56), .ZN(new_n818_));
  INV_X1    g617(.A(new_n546_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n570_), .A2(new_n579_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n571_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n568_), .A2(new_n821_), .A3(new_n569_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n567_), .B1(new_n578_), .B2(new_n565_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n567_), .B(KEYINPUT118), .C1(new_n578_), .C2(new_n565_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n822_), .B1(new_n827_), .B2(new_n821_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n820_), .B1(new_n828_), .B2(new_n819_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n283_), .C1(new_n811_), .C2(new_n816_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n818_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n818_), .A2(KEYINPUT58), .A3(new_n830_), .A4(new_n832_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n629_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n831_), .A2(KEYINPUT117), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n817_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n838_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n283_), .B(new_n840_), .C1(new_n811_), .C2(new_n816_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n839_), .A2(new_n287_), .A3(new_n660_), .A4(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n829_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n667_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT57), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n841_), .A2(new_n287_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n586_), .B1(new_n817_), .B2(new_n838_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n843_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n847_), .B1(new_n850_), .B2(new_n667_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n837_), .A2(new_n846_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n648_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n628_), .A2(new_n647_), .A3(new_n292_), .A4(new_n586_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n855_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n540_), .A2(new_n347_), .A3(new_n538_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n859_), .A2(KEYINPUT120), .A3(new_n860_), .A4(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n852_), .A2(new_n648_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n860_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n863_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(G113gat), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT121), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871_));
  OAI21_X1  g670(.A(G113gat), .B1(new_n586_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n855_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n854_), .B(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n845_), .B2(KEYINPUT57), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT119), .B(new_n847_), .C1(new_n850_), .C2(new_n667_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n876_), .A2(new_n846_), .A3(new_n837_), .A4(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n874_), .B1(new_n878_), .B2(new_n648_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT59), .B1(new_n879_), .B2(new_n861_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n868_), .A2(new_n870_), .A3(new_n872_), .A4(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n861_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n869_), .B1(new_n883_), .B2(new_n586_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n881_), .A2(new_n884_), .ZN(G1340gat));
  INV_X1    g684(.A(G120gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n292_), .B2(KEYINPUT60), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n882_), .B(new_n887_), .C1(KEYINPUT60), .C2(new_n886_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n868_), .A2(new_n709_), .A3(new_n880_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n886_), .ZN(G1341gat));
  NAND4_X1  g689(.A1(new_n868_), .A2(G127gat), .A3(new_n647_), .A4(new_n880_), .ZN(new_n891_));
  INV_X1    g690(.A(G127gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n883_), .B2(new_n648_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT122), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n891_), .A2(new_n896_), .A3(new_n893_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1342gat));
  NAND2_X1  g697(.A1(new_n882_), .A2(new_n667_), .ZN(new_n899_));
  INV_X1    g698(.A(G134gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n901_), .A2(KEYINPUT123), .ZN(new_n902_));
  AND4_X1   g701(.A1(G134gat), .A2(new_n868_), .A3(new_n629_), .A4(new_n880_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n901_), .A2(KEYINPUT123), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(G1343gat));
  NAND2_X1  g704(.A1(new_n878_), .A2(new_n648_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n858_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n539_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n502_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n678_), .A2(new_n493_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n909_), .A2(new_n660_), .A3(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g711(.A1(new_n909_), .A2(new_n709_), .A3(new_n910_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g713(.A1(new_n909_), .A2(new_n647_), .A3(new_n910_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT61), .B(G155gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1346gat));
  AND3_X1   g716(.A1(new_n909_), .A2(G162gat), .A3(new_n910_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n909_), .A2(new_n667_), .A3(new_n910_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n918_), .A2(new_n629_), .B1(new_n919_), .B2(new_n610_), .ZN(G1347gat));
  NAND2_X1  g719(.A1(new_n678_), .A2(new_n541_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n865_), .A2(new_n503_), .A3(new_n921_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n922_), .A2(new_n660_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  OR3_X1    g723(.A1(new_n923_), .A2(new_n924_), .A3(new_n377_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n923_), .B1(new_n365_), .B2(new_n363_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n924_), .B1(new_n923_), .B2(new_n377_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(G1348gat));
  AOI21_X1  g727(.A(G176gat), .B1(new_n922_), .B2(new_n709_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n907_), .A2(KEYINPUT124), .A3(new_n493_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n931_), .B1(new_n879_), .B2(new_n503_), .ZN(new_n932_));
  AOI211_X1 g731(.A(new_n359_), .B(new_n292_), .C1(new_n930_), .C2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n921_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n929_), .B1(new_n933_), .B2(new_n934_), .ZN(G1349gat));
  NOR2_X1   g734(.A1(new_n648_), .A2(new_n369_), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n922_), .A2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n930_), .A2(new_n932_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n921_), .A2(new_n648_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n940_), .ZN(new_n942_));
  AOI211_X1 g741(.A(KEYINPUT125), .B(new_n942_), .C1(new_n930_), .C2(new_n932_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n941_), .A2(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n937_), .B1(new_n944_), .B2(new_n348_), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n667_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n946_));
  XOR2_X1   g745(.A(new_n946_), .B(KEYINPUT126), .Z(new_n947_));
  NAND2_X1  g746(.A1(new_n922_), .A2(new_n947_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n922_), .A2(new_n629_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(new_n349_), .ZN(G1351gat));
  NAND4_X1  g749(.A1(new_n907_), .A2(new_n656_), .A3(new_n678_), .A4(new_n539_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n660_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g753(.A1(new_n952_), .A2(new_n709_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g755(.A1(new_n951_), .A2(new_n648_), .ZN(new_n957_));
  XOR2_X1   g756(.A(KEYINPUT63), .B(G211gat), .Z(new_n958_));
  AND3_X1   g757(.A1(new_n957_), .A2(KEYINPUT127), .A3(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n958_), .ZN(new_n960_));
  OR2_X1    g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  OAI21_X1  g760(.A(KEYINPUT127), .B1(new_n957_), .B2(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n959_), .B1(new_n960_), .B2(new_n962_), .ZN(G1354gat));
  NOR3_X1   g762(.A1(new_n951_), .A2(new_n390_), .A3(new_n628_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n952_), .A2(new_n667_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n964_), .B1(new_n390_), .B2(new_n965_), .ZN(G1355gat));
endmodule


