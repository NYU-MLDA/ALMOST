//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n929_, new_n930_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(G204gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT5), .B(G176gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  XNOR2_X1  g005(.A(G57gat), .B(G64gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT11), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(KEYINPUT11), .ZN(new_n209_));
  XOR2_X1   g008(.A(G71gat), .B(G78gat), .Z(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n209_), .A2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT65), .B1(new_n214_), .B2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT10), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT10), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(G99gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n215_), .A2(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  NOR3_X1   g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT6), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(G85gat), .A3(G92gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n228_), .A2(new_n234_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n224_), .A2(KEYINPUT66), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT66), .B1(new_n224_), .B2(new_n235_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT7), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(new_n216_), .A3(new_n222_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n240_), .A2(new_n231_), .A3(new_n233_), .A4(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n225_), .A2(new_n226_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT8), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(KEYINPUT67), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n242_), .B(new_n243_), .C1(KEYINPUT67), .C2(new_n245_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n213_), .B1(new_n238_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT12), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G230gat), .A2(G233gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT64), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n238_), .A2(new_n249_), .A3(new_n213_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n221_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n257_));
  AOI211_X1 g056(.A(KEYINPUT65), .B(G106gat), .C1(new_n217_), .C2(new_n219_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n235_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n224_), .A2(KEYINPUT66), .A3(new_n235_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n249_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n213_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n251_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n252_), .A2(new_n255_), .A3(new_n256_), .A4(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n263_), .A2(new_n264_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n264_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT68), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n271_), .B1(new_n273_), .B2(KEYINPUT12), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n274_), .A2(KEYINPUT69), .A3(new_n255_), .A4(new_n267_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n255_), .B1(new_n256_), .B2(new_n272_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n206_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n206_), .ZN(new_n280_));
  AOI211_X1 g079(.A(new_n277_), .B(new_n280_), .C1(new_n270_), .C2(new_n275_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT13), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT70), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G229gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G43gat), .B(G50gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT71), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G29gat), .B(G36gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n291_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n293_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G15gat), .B(G22gat), .ZN(new_n301_));
  INV_X1    g100(.A(G1gat), .ZN(new_n302_));
  INV_X1    g101(.A(G8gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT14), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G1gat), .B(G8gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  NAND2_X1  g106(.A1(new_n300_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n299_), .B(KEYINPUT15), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n290_), .B(new_n308_), .C1(new_n309_), .C2(new_n307_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n299_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n290_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G113gat), .B(G141gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G169gat), .B(G197gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n310_), .A2(new_n315_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n310_), .A2(new_n315_), .A3(KEYINPUT75), .A4(new_n321_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n320_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n289_), .A2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G71gat), .B(G99gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT78), .B(G15gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G227gat), .A2(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(G43gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n331_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT25), .B(G183gat), .ZN(new_n336_));
  INV_X1    g135(.A(G190gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT26), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G190gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(KEYINPUT76), .A3(KEYINPUT26), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n336_), .A2(new_n340_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT23), .ZN(new_n346_));
  INV_X1    g145(.A(G169gat), .ZN(new_n347_));
  INV_X1    g146(.A(G176gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(KEYINPUT24), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT24), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n346_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G183gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n337_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n346_), .A2(new_n356_), .B1(G169gat), .B2(G176gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n358_), .A2(new_n347_), .A3(KEYINPUT22), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT22), .B1(new_n358_), .B2(new_n347_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n348_), .A3(new_n360_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n344_), .A2(new_n354_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT30), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(KEYINPUT79), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(KEYINPUT79), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n335_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n365_), .B2(new_n335_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT80), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G127gat), .B(G134gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G113gat), .B(G120gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n371_), .B(KEYINPUT31), .Z(new_n372_));
  NOR2_X1   g171(.A1(new_n368_), .A2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n368_), .A2(new_n372_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n367_), .A2(KEYINPUT80), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n371_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(KEYINPUT81), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(KEYINPUT3), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n379_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(new_n385_));
  NOR2_X1   g184(.A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(new_n386_));
  OAI211_X1 g185(.A(G141gat), .B(G148gat), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(KEYINPUT3), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n388_), .A2(new_n378_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n384_), .A2(new_n387_), .A3(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G155gat), .B(G162gat), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G155gat), .ZN(new_n395_));
  INV_X1    g194(.A(G162gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT1), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(G155gat), .B2(G162gat), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n395_), .A2(new_n396_), .A3(KEYINPUT1), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n379_), .B(new_n389_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n394_), .A2(KEYINPUT83), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT83), .B1(new_n394_), .B2(new_n400_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n377_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n394_), .A2(new_n400_), .A3(new_n371_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(KEYINPUT4), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n406_), .B(new_n377_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT96), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413_));
  INV_X1    g212(.A(G85gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT0), .B(G57gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n405_), .A2(KEYINPUT96), .A3(new_n407_), .A4(new_n409_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n403_), .A2(new_n404_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(new_n409_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n412_), .A2(new_n418_), .A3(new_n419_), .A4(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n418_), .B1(new_n425_), .B2(new_n419_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G22gat), .B(G50gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n401_), .A2(new_n402_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n394_), .A2(new_n400_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n394_), .A2(KEYINPUT83), .A3(new_n400_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n434_), .A3(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n431_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n430_), .B1(new_n435_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n433_), .A2(new_n434_), .A3(new_n432_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n431_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n429_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT88), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n434_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT87), .B1(new_n203_), .B2(G197gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n451_));
  INV_X1    g250(.A(G197gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(G204gat), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n450_), .A2(new_n453_), .B1(G197gat), .B2(new_n203_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT21), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT86), .B1(new_n452_), .B2(G204gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(G204gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n203_), .A2(G197gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(KEYINPUT86), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT21), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G211gat), .B(G218gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n456_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n454_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n463_), .A2(new_n455_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(KEYINPUT85), .A2(G233gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(KEYINPUT85), .A2(G233gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(G228gat), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n448_), .B1(new_n449_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT29), .B1(new_n401_), .B2(new_n402_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n473_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(KEYINPUT88), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n436_), .A2(KEYINPUT29), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n472_), .B1(new_n479_), .B2(new_n468_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n447_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n447_), .ZN(new_n483_));
  AOI211_X1 g282(.A(new_n480_), .B(new_n483_), .C1(new_n474_), .C2(new_n477_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n446_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n446_), .B(KEYINPUT90), .C1(new_n482_), .C2(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n449_), .A2(new_n448_), .A3(new_n473_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT88), .B1(new_n475_), .B2(new_n476_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n481_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n483_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n442_), .A2(new_n445_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n478_), .A2(new_n481_), .A3(new_n447_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n493_), .A2(new_n494_), .A3(KEYINPUT89), .A4(new_n495_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n489_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G226gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT19), .ZN(new_n503_));
  INV_X1    g302(.A(new_n463_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n504_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n505_), .A2(new_n462_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n352_), .A2(KEYINPUT92), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n352_), .A2(KEYINPUT92), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n347_), .B(new_n348_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n509_), .A2(new_n346_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n342_), .A2(new_n338_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n342_), .B2(new_n338_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n336_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT93), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n350_), .A3(new_n349_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n510_), .A2(new_n515_), .A3(new_n516_), .A4(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n509_), .A2(new_n518_), .A3(new_n346_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n336_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n342_), .A2(new_n338_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT91), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n523_), .B2(new_n512_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT93), .B1(new_n520_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G169gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n348_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n357_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n506_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n354_), .A2(new_n344_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n357_), .A2(new_n361_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT20), .B1(new_n533_), .B2(new_n468_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n503_), .B1(new_n530_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n503_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT20), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n533_), .B2(new_n468_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n526_), .A2(new_n529_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n538_), .B1(new_n539_), .B2(new_n468_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n535_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G8gat), .B(G36gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  XNOR2_X1  g343(.A(G64gat), .B(G92gat), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n544_), .A2(new_n545_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n541_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n548_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n535_), .A2(new_n550_), .A3(new_n540_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(KEYINPUT95), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT27), .ZN(new_n553_));
  INV_X1    g352(.A(new_n541_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(new_n550_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT103), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n552_), .A2(new_n556_), .A3(KEYINPUT103), .A4(new_n553_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT101), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n529_), .B1(new_n524_), .B2(new_n520_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n468_), .B1(new_n562_), .B2(KEYINPUT98), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n529_), .B(new_n564_), .C1(new_n524_), .C2(new_n520_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT20), .B1(new_n362_), .B2(new_n506_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n503_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n567_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT99), .B1(new_n572_), .B2(new_n536_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n534_), .B1(new_n539_), .B2(new_n468_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n536_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n561_), .B1(new_n576_), .B2(new_n548_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n551_), .A2(KEYINPUT102), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT102), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n535_), .A2(new_n579_), .A3(new_n550_), .A4(new_n540_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(KEYINPUT27), .A3(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n577_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n576_), .A2(new_n561_), .A3(new_n548_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n559_), .A2(new_n560_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n376_), .A2(new_n428_), .A3(new_n501_), .A4(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT32), .B1(new_n546_), .B2(new_n547_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(KEYINPUT97), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n576_), .A2(new_n587_), .B1(new_n554_), .B2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT100), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n423_), .A2(KEYINPUT33), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT33), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n425_), .A2(new_n593_), .A3(new_n418_), .A4(new_n419_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n417_), .B1(new_n420_), .B2(new_n408_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n407_), .A2(new_n408_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n405_), .B2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n552_), .B2(new_n556_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n589_), .B(new_n601_), .C1(new_n424_), .C2(new_n426_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n591_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n427_), .B1(new_n489_), .B2(new_n500_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n603_), .A2(new_n501_), .B1(new_n604_), .B2(new_n584_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n585_), .B1(new_n605_), .B2(new_n376_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n328_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT34), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT35), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT15), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n299_), .B(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n263_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n238_), .A2(new_n300_), .A3(new_n249_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT72), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n615_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n610_), .B(KEYINPUT35), .Z(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI22_X1  g419(.A1(new_n616_), .A2(new_n617_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(new_n617_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  NAND4_X1  g426(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .A4(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n624_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n627_), .A2(new_n624_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n623_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n629_), .B(new_n630_), .C1(new_n631_), .C2(new_n621_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n628_), .A2(KEYINPUT37), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT37), .B1(new_n628_), .B2(new_n632_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n307_), .B(new_n213_), .Z(new_n637_));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(KEYINPUT74), .ZN(new_n640_));
  XOR2_X1   g439(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n641_));
  XNOR2_X1  g440(.A(G127gat), .B(G155gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(G183gat), .B(G211gat), .Z(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT17), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n640_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n645_), .A2(KEYINPUT17), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n639_), .A2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n650_), .B1(new_n640_), .B2(new_n646_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n636_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n608_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n427_), .A2(new_n302_), .ZN(new_n656_));
  OR3_X1    g455(.A1(new_n654_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n628_), .A2(new_n632_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n652_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n608_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n428_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n655_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n657_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT104), .ZN(G1324gat));
  NAND2_X1  g464(.A1(new_n322_), .A2(new_n323_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n666_), .A2(new_n325_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n288_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n584_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n606_), .A4(new_n660_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G8gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT39), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n608_), .A2(new_n303_), .A3(new_n669_), .A4(new_n653_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1325gat));
  INV_X1    g475(.A(new_n376_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G15gat), .B1(new_n661_), .B2(new_n677_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(KEYINPUT41), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT41), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n654_), .A2(G15gat), .A3(new_n677_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(G1326gat));
  OR3_X1    g481(.A1(new_n654_), .A2(G22gat), .A3(new_n501_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G22gat), .B1(new_n661_), .B2(new_n501_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(KEYINPUT42), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(KEYINPUT42), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(G1327gat));
  INV_X1    g486(.A(new_n652_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(new_n658_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n608_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(G29gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n427_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n606_), .B2(new_n636_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n604_), .A2(new_n584_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n489_), .A2(new_n500_), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n590_), .A2(KEYINPUT100), .B1(new_n595_), .B2(new_n599_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n602_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n677_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n635_), .B1(new_n702_), .B2(new_n585_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT107), .B(new_n697_), .C1(new_n703_), .C2(new_n693_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n695_), .B1(new_n607_), .B2(new_n635_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n696_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n328_), .A2(new_n688_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(KEYINPUT44), .A3(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT44), .B1(new_n706_), .B2(new_n707_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n428_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n692_), .B1(new_n710_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n608_), .A2(new_n712_), .A3(new_n669_), .A4(new_n689_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT45), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n708_), .A2(new_n709_), .A3(new_n584_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n712_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n714_), .B(KEYINPUT46), .C1(new_n715_), .C2(new_n712_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1329gat));
  INV_X1    g519(.A(new_n709_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n706_), .A2(KEYINPUT44), .A3(new_n707_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n721_), .A2(G43gat), .A3(new_n376_), .A4(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n690_), .A2(new_n376_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n333_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT47), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n723_), .A2(new_n728_), .A3(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1330gat));
  INV_X1    g529(.A(G50gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n690_), .A2(new_n731_), .A3(new_n699_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n721_), .A2(new_n699_), .A3(new_n722_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT108), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G50gat), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n733_), .A2(KEYINPUT108), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1331gat));
  NOR3_X1   g536(.A1(new_n289_), .A2(new_n607_), .A3(new_n327_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n660_), .ZN(new_n739_));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n428_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n288_), .A2(new_n653_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n742_), .A2(KEYINPUT109), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n607_), .A2(new_n327_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(KEYINPUT109), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n746_), .A2(new_n428_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n741_), .B1(new_n747_), .B2(new_n740_), .ZN(G1332gat));
  OR3_X1    g547(.A1(new_n746_), .A2(G64gat), .A3(new_n584_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G64gat), .B1(new_n739_), .B2(new_n584_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(KEYINPUT48), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(KEYINPUT48), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n751_), .B2(new_n752_), .ZN(G1333gat));
  OR3_X1    g552(.A1(new_n746_), .A2(G71gat), .A3(new_n677_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G71gat), .B1(new_n739_), .B2(new_n677_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT49), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(KEYINPUT49), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n756_), .B2(new_n757_), .ZN(G1334gat));
  OR3_X1    g557(.A1(new_n746_), .A2(G78gat), .A3(new_n501_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G78gat), .B1(new_n739_), .B2(new_n501_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(KEYINPUT50), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(KEYINPUT50), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(G1335gat));
  AND2_X1   g562(.A1(new_n738_), .A2(new_n689_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G85gat), .B1(new_n764_), .B2(new_n427_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n289_), .A2(new_n327_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n706_), .A2(new_n652_), .A3(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n428_), .A2(new_n414_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n765_), .B1(new_n767_), .B2(new_n768_), .ZN(G1336gat));
  AOI21_X1  g568(.A(G92gat), .B1(new_n764_), .B2(new_n669_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n669_), .A2(G92gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n767_), .B2(new_n771_), .ZN(G1337gat));
  AOI21_X1  g571(.A(new_n216_), .B1(new_n767_), .B2(new_n376_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n764_), .A2(new_n220_), .A3(new_n376_), .ZN(new_n774_));
  OR3_X1    g573(.A1(new_n773_), .A2(new_n774_), .A3(KEYINPUT51), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT51), .B1(new_n773_), .B2(new_n774_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n764_), .A2(new_n222_), .A3(new_n699_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n706_), .A2(new_n699_), .A3(new_n652_), .A4(new_n766_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(G106gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(G106gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n778_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  NAND3_X1  g586(.A1(new_n653_), .A2(new_n667_), .A3(new_n284_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT54), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n314_), .B(new_n308_), .C1(new_n309_), .C2(new_n307_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n321_), .B1(new_n313_), .B2(new_n290_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n792_), .A2(KEYINPUT114), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(KEYINPUT114), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n324_), .A2(new_n326_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n282_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT113), .B1(new_n268_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n256_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n251_), .B(KEYINPUT12), .C1(new_n263_), .C2(new_n264_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(KEYINPUT55), .A4(new_n255_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n254_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT112), .B(new_n254_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n798_), .A2(new_n803_), .A3(new_n806_), .A4(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n270_), .B2(new_n275_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n280_), .B1(new_n808_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT56), .B(new_n280_), .C1(new_n808_), .C2(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n281_), .A2(new_n667_), .A3(KEYINPUT110), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n276_), .A2(new_n278_), .A3(new_n206_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n327_), .B2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n796_), .B1(new_n816_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT57), .B1(new_n822_), .B2(new_n659_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT110), .B1(new_n281_), .B2(new_n667_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n327_), .A2(new_n819_), .A3(new_n818_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n824_), .B(new_n658_), .C1(new_n828_), .C2(new_n796_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n795_), .A2(new_n281_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n816_), .A2(KEYINPUT58), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT69), .B1(new_n801_), .B2(new_n255_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n268_), .A2(new_n269_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n809_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n806_), .A2(new_n807_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n803_), .A4(new_n798_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT56), .B1(new_n836_), .B2(new_n280_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n815_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n635_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n823_), .A2(new_n829_), .B1(new_n831_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n652_), .B1(new_n842_), .B2(KEYINPUT115), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n823_), .A2(new_n829_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n831_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n844_), .A2(KEYINPUT115), .A3(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n789_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n376_), .A2(new_n501_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n848_), .A2(new_n428_), .A3(new_n669_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n327_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n842_), .A2(new_n688_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n789_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n850_), .B2(KEYINPUT59), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n667_), .A2(KEYINPUT116), .ZN(new_n858_));
  MUX2_X1   g657(.A(KEYINPUT116), .B(new_n858_), .S(G113gat), .Z(new_n859_));
  AOI21_X1  g658(.A(new_n852_), .B1(new_n857_), .B2(new_n859_), .ZN(G1340gat));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n861_), .A3(new_n288_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G120gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n857_), .B2(new_n288_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n865_));
  AOI21_X1  g664(.A(G120gat), .B1(new_n288_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n865_), .B2(G120gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT117), .B1(new_n851_), .B2(new_n867_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n851_), .A2(KEYINPUT117), .A3(new_n867_), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n863_), .A2(new_n864_), .B1(new_n868_), .B2(new_n869_), .ZN(G1341gat));
  INV_X1    g669(.A(G127gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n857_), .B2(new_n688_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n850_), .A2(G127gat), .A3(new_n652_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT119), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n873_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876_));
  AOI211_X1 g675(.A(new_n652_), .B(new_n856_), .C1(new_n850_), .C2(KEYINPUT59), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n875_), .B(new_n876_), .C1(new_n877_), .C2(new_n871_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n878_), .ZN(G1342gat));
  AOI21_X1  g678(.A(G134gat), .B1(new_n851_), .B2(new_n659_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n636_), .A2(G134gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n857_), .B2(new_n881_), .ZN(G1343gat));
  NOR4_X1   g681(.A1(new_n669_), .A2(new_n376_), .A3(new_n501_), .A4(new_n428_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n847_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT120), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n847_), .A2(new_n886_), .A3(new_n883_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n667_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(G141gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1344gat));
  AOI21_X1  g689(.A(new_n289_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT121), .B(G148gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1345gat));
  NAND2_X1  g692(.A1(new_n885_), .A2(new_n887_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n894_), .A2(new_n688_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n894_), .B2(new_n688_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1346gat));
  AOI21_X1  g697(.A(G162gat), .B1(new_n894_), .B2(new_n659_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n635_), .A2(new_n396_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n894_), .B2(new_n900_), .ZN(G1347gat));
  NAND2_X1  g700(.A1(new_n855_), .A2(new_n789_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n848_), .A2(new_n427_), .A3(new_n584_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n347_), .B1(new_n904_), .B2(new_n327_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n905_), .A2(KEYINPUT62), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(KEYINPUT62), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n904_), .A2(new_n327_), .A3(new_n527_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n904_), .B2(new_n288_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n288_), .A2(G176gat), .A3(new_n903_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n847_), .B2(new_n911_), .ZN(G1349gat));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n904_), .A2(new_n913_), .A3(new_n521_), .A4(new_n688_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n902_), .A2(new_n688_), .A3(new_n903_), .ZN(new_n915_));
  AOI21_X1  g714(.A(KEYINPUT122), .B1(new_n915_), .B2(new_n355_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n336_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n914_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT123), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n914_), .B(new_n920_), .C1(new_n916_), .C2(new_n917_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1350gat));
  OAI211_X1 g721(.A(new_n904_), .B(new_n659_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n904_), .A2(new_n636_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(G190gat), .ZN(new_n926_));
  AOI211_X1 g725(.A(KEYINPUT124), .B(new_n337_), .C1(new_n904_), .C2(new_n636_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n923_), .B1(new_n926_), .B2(new_n927_), .ZN(G1351gat));
  AND4_X1   g727(.A1(new_n604_), .A2(new_n847_), .A3(new_n669_), .A4(new_n677_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n327_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n288_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g732(.A(new_n652_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT125), .ZN(new_n935_));
  OR2_X1    g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n929_), .A2(new_n935_), .B1(KEYINPUT126), .B2(new_n936_), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n936_), .A2(KEYINPUT126), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n937_), .B(new_n938_), .ZN(G1354gat));
  AOI21_X1  g738(.A(G218gat), .B1(new_n929_), .B2(new_n659_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n636_), .A2(G218gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT127), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n929_), .B2(new_n942_), .ZN(G1355gat));
endmodule


