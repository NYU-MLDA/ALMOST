//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT6), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT65), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT7), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G85gat), .B(G92gat), .Z(new_n209_));
  INV_X1    g008(.A(KEYINPUT8), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(new_n204_), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n212_), .A2(new_n209_), .ZN(new_n213_));
  OAI22_X1  g012(.A1(new_n208_), .A2(new_n211_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT10), .B(G99gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G106gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  OR3_X1    g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT9), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n209_), .A2(KEYINPUT9), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n205_), .A2(new_n217_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n214_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G43gat), .B(G50gat), .Z(new_n224_));
  XNOR2_X1  g023(.A(G29gat), .B(G36gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n202_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n214_), .A2(KEYINPUT73), .A3(new_n222_), .A4(new_n228_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G232gat), .A2(G233gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT68), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT34), .ZN(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n235_));
  OR2_X1    g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n230_), .A2(new_n231_), .A3(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n228_), .B(KEYINPUT15), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n223_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n234_), .A2(new_n235_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT70), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n237_), .A2(new_n240_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G134gat), .B(G162gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT76), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(G190gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(G218gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT36), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT77), .Z(new_n252_));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n237_), .A2(new_n253_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n230_), .A2(KEYINPUT74), .A3(new_n231_), .A4(new_n236_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(new_n239_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n256_), .A2(KEYINPUT75), .A3(new_n243_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT75), .B1(new_n256_), .B2(new_n243_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n245_), .B(new_n252_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT37), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n243_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT75), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n256_), .A2(KEYINPUT75), .A3(new_n243_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n244_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n249_), .B(KEYINPUT36), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT78), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n259_), .B(new_n260_), .C1(new_n265_), .C2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n245_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n267_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n260_), .B1(new_n272_), .B2(new_n259_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G127gat), .B(G155gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT16), .ZN(new_n276_));
  INV_X1    g075(.A(G183gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G211gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT17), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n280_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G15gat), .B(G22gat), .ZN(new_n284_));
  INV_X1    g083(.A(G1gat), .ZN(new_n285_));
  INV_X1    g084(.A(G8gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT14), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G1gat), .B(G8gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G231gat), .A2(G233gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n290_), .B(new_n291_), .Z(new_n292_));
  XNOR2_X1  g091(.A(G57gat), .B(G64gat), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n293_), .A2(KEYINPUT11), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(KEYINPUT11), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G71gat), .B(G78gat), .ZN(new_n296_));
  OR3_X1    g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n296_), .A3(KEYINPUT11), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n292_), .B(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n282_), .A2(new_n283_), .A3(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n299_), .B(KEYINPUT66), .Z(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(new_n292_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n292_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n281_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n274_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT79), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  OR2_X1    g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT1), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT94), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT95), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(KEYINPUT94), .A3(KEYINPUT1), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .A4(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT96), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(new_n315_), .B2(KEYINPUT1), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n326_), .A2(KEYINPUT96), .A3(G155gat), .A4(G162gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n321_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n319_), .B1(new_n330_), .B2(new_n320_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n314_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT97), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT97), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n334_), .B(new_n314_), .C1(new_n329_), .C2(new_n331_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n322_), .A2(new_n315_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT2), .ZN(new_n338_));
  OAI22_X1  g137(.A1(new_n312_), .A2(KEYINPUT3), .B1(new_n338_), .B2(new_n313_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n312_), .A2(KEYINPUT3), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT98), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n312_), .A2(KEYINPUT98), .A3(KEYINPUT3), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n339_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n313_), .A2(new_n338_), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT99), .Z(new_n346_));
  AOI21_X1  g145(.A(new_n337_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G113gat), .B(G120gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT103), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n351_), .A2(KEYINPUT103), .ZN(new_n353_));
  AND4_X1   g152(.A1(new_n336_), .A2(new_n348_), .A3(new_n352_), .A4(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n347_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n352_), .B1(new_n355_), .B2(new_n353_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n311_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT0), .ZN(new_n359_));
  INV_X1    g158(.A(G57gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(new_n218_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT104), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT4), .B1(new_n354_), .B2(new_n356_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n311_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n351_), .A2(KEYINPUT4), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n355_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n366_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n318_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT95), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n323_), .A3(new_n328_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n334_), .B1(new_n376_), .B2(new_n314_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n335_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n348_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(KEYINPUT103), .A3(new_n351_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n355_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n373_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n382_), .A2(KEYINPUT104), .A3(new_n370_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n365_), .B1(new_n372_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT33), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(KEYINPUT105), .A3(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT104), .B1(new_n382_), .B2(new_n370_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n367_), .A2(new_n366_), .A3(new_n371_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n364_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT105), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT33), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT86), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT86), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(G169gat), .A3(G176gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT23), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G176gat), .ZN(new_n404_));
  INV_X1    g203(.A(G169gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT22), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n407_), .B2(KEYINPUT89), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n409_), .B1(new_n405_), .B2(KEYINPUT22), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT22), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(KEYINPUT90), .A3(G169gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n410_), .B(new_n412_), .C1(new_n413_), .C2(new_n406_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n397_), .B(new_n403_), .C1(new_n408_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT84), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(G190gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n277_), .A2(KEYINPUT82), .A3(KEYINPUT25), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT82), .B1(new_n277_), .B2(KEYINPUT25), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n418_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT83), .B1(new_n277_), .B2(KEYINPUT25), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT25), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(new_n425_), .A3(G183gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n417_), .B1(new_n422_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n421_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n419_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n431_), .A2(KEYINPUT84), .A3(new_n427_), .A4(new_n418_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n405_), .A2(new_n404_), .A3(KEYINPUT85), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(G169gat), .B2(G176gat), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n433_), .A2(new_n435_), .A3(KEYINPUT24), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n397_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n433_), .A2(new_n435_), .A3(KEYINPUT24), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT87), .B1(new_n439_), .B2(new_n396_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n429_), .A2(new_n432_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n398_), .B(KEYINPUT23), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n433_), .A2(new_n435_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n442_), .B(new_n443_), .C1(new_n444_), .C2(KEYINPUT24), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT24), .B1(new_n433_), .B2(new_n435_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n398_), .B(new_n399_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT88), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n416_), .B1(new_n441_), .B2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G197gat), .B(G204gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(G211gat), .B(G218gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(KEYINPUT21), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(KEYINPUT21), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT102), .B1(new_n450_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n429_), .A2(new_n432_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n438_), .A2(new_n440_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n449_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n415_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT102), .ZN(new_n461_));
  INV_X1    g260(.A(new_n455_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n456_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n403_), .A2(KEYINPUT100), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT100), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n400_), .A2(new_n401_), .A3(new_n466_), .A4(new_n402_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n411_), .A2(G169gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n406_), .A2(new_n468_), .A3(new_n404_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n465_), .A2(new_n397_), .A3(new_n467_), .A4(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT101), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n436_), .A2(new_n392_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n447_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n425_), .A2(G183gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n277_), .A2(KEYINPUT25), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n418_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n473_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n406_), .A2(new_n468_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n396_), .B1(new_n480_), .B2(new_n404_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n481_), .A2(KEYINPUT101), .A3(new_n467_), .A4(new_n465_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n472_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n483_), .A2(new_n462_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G226gat), .A2(G233gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT19), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n464_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n450_), .A2(new_n455_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n485_), .B1(new_n483_), .B2(new_n462_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n487_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G8gat), .B(G36gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT18), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G64gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(new_n219_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n489_), .A2(new_n493_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n354_), .A2(new_n356_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n311_), .B1(new_n355_), .B2(new_n369_), .ZN(new_n502_));
  OAI221_X1 g301(.A(new_n362_), .B1(new_n501_), .B2(new_n311_), .C1(new_n382_), .C2(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n386_), .A2(new_n391_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n387_), .A2(new_n388_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n363_), .B1(new_n506_), .B2(new_n357_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n384_), .A2(KEYINPUT106), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT106), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n389_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n507_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n464_), .A2(new_n488_), .B1(new_n492_), .B2(new_n487_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n497_), .A2(KEYINPUT32), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n487_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n490_), .A2(new_n515_), .A3(new_n491_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n455_), .A2(new_n479_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n470_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT20), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n464_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n517_), .B1(new_n522_), .B2(new_n487_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n514_), .B1(new_n523_), .B2(new_n513_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n505_), .B1(new_n511_), .B2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G22gat), .B(G50gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT28), .ZN(new_n527_));
  XOR2_X1   g326(.A(G78gat), .B(G106gat), .Z(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT29), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n462_), .B1(new_n355_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G228gat), .A2(G233gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n533_), .B(new_n462_), .C1(new_n355_), .C2(new_n531_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n379_), .A2(KEYINPUT29), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n535_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n538_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n530_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n536_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n537_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n529_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n525_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT27), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT107), .ZN(new_n550_));
  INV_X1    g349(.A(new_n497_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n515_), .B1(new_n464_), .B2(new_n521_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n550_), .B(new_n551_), .C1(new_n552_), .C2(new_n517_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n548_), .B1(new_n512_), .B2(new_n497_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n520_), .B1(new_n456_), .B2(new_n463_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n516_), .B1(new_n556_), .B2(new_n515_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n550_), .B1(new_n557_), .B2(new_n551_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n549_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(new_n546_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n511_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n547_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n460_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n450_), .A2(KEYINPUT30), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n563_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n566_), .A3(new_n563_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G71gat), .B(G99gat), .Z(new_n570_));
  NAND2_X1  g369(.A1(G227gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G15gat), .B(G43gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n569_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n569_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(new_n567_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n351_), .B(KEYINPUT31), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n579_), .B1(new_n581_), .B2(KEYINPUT92), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n575_), .A2(new_n578_), .A3(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n582_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n541_), .A2(new_n545_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT108), .B1(new_n559_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT108), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT107), .B1(new_n523_), .B2(new_n497_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n546_), .A2(new_n591_), .A3(new_n593_), .A4(new_n549_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n357_), .B1(new_n372_), .B2(new_n383_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n362_), .ZN(new_n597_));
  AOI211_X1 g396(.A(KEYINPUT106), .B(new_n364_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n509_), .B1(new_n506_), .B2(new_n365_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n597_), .B(new_n587_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT109), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT109), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n595_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n562_), .A2(new_n588_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n310_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n223_), .A2(new_n300_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT12), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n214_), .A2(new_n222_), .A3(new_n299_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n303_), .A2(KEYINPUT12), .A3(new_n223_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .A4(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n612_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n611_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n619_));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n621_), .B(new_n622_), .Z(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n614_), .A2(new_n617_), .A3(new_n623_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n628_), .A2(KEYINPUT13), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(KEYINPUT13), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n228_), .B(new_n290_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G229gat), .A2(G233gat), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n229_), .A2(new_n290_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(new_n633_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n238_), .A2(new_n290_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(KEYINPUT81), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G113gat), .B(G141gat), .ZN(new_n640_));
  INV_X1    g439(.A(G197gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT80), .B(G169gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n639_), .B(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n631_), .A2(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n607_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n511_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n285_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n272_), .A2(new_n259_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n606_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n648_), .A3(new_n308_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n511_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n651_), .A2(KEYINPUT110), .A3(new_n652_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT110), .B1(new_n651_), .B2(new_n652_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n653_), .B(new_n658_), .C1(new_n659_), .C2(new_n660_), .ZN(G1324gat));
  INV_X1    g460(.A(KEYINPUT40), .ZN(new_n662_));
  INV_X1    g461(.A(new_n559_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G8gat), .B1(new_n657_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT39), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT111), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n607_), .A2(new_n286_), .A3(new_n648_), .A4(new_n559_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n666_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n662_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n665_), .A2(new_n667_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT111), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(KEYINPUT40), .A3(new_n668_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n674_), .ZN(G1325gat));
  OAI21_X1  g474(.A(G15gat), .B1(new_n657_), .B2(new_n588_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT41), .Z(new_n677_));
  INV_X1    g476(.A(G15gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n649_), .A2(new_n678_), .A3(new_n587_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1326gat));
  INV_X1    g479(.A(G22gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n649_), .A2(new_n681_), .A3(new_n589_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G22gat), .B1(new_n657_), .B2(new_n546_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT42), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1327gat));
  NOR3_X1   g484(.A1(new_n606_), .A2(new_n654_), .A3(new_n308_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(new_n648_), .ZN(new_n687_));
  INV_X1    g486(.A(G29gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n650_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT114), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n270_), .A2(new_n273_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n595_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n604_), .B1(new_n595_), .B2(new_n601_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n587_), .B1(new_n547_), .B2(new_n561_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n691_), .B(new_n692_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT112), .ZN(new_n698_));
  AOI22_X1  g497(.A1(new_n525_), .A2(new_n546_), .B1(new_n511_), .B2(new_n560_), .ZN(new_n699_));
  OAI22_X1  g498(.A1(new_n699_), .A2(new_n587_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT112), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n691_), .A4(new_n692_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n606_), .B2(new_n274_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n698_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(new_n648_), .A3(new_n307_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT113), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n704_), .A2(KEYINPUT113), .A3(new_n648_), .A4(new_n307_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n704_), .A2(KEYINPUT44), .A3(new_n648_), .A4(new_n307_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n650_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n690_), .B1(new_n713_), .B2(G29gat), .ZN(new_n714_));
  AOI211_X1 g513(.A(KEYINPUT114), .B(new_n688_), .C1(new_n710_), .C2(new_n712_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n689_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  NOR2_X1   g515(.A1(new_n663_), .A2(G36gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n686_), .A2(new_n648_), .A3(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT115), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT45), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n711_), .A2(new_n559_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n710_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(G36gat), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n720_), .B(KEYINPUT46), .C1(new_n722_), .C2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n719_), .B(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n723_), .B1(new_n710_), .B2(new_n721_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n724_), .A2(new_n729_), .ZN(G1329gat));
  INV_X1    g529(.A(G43gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n711_), .A2(new_n587_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n710_), .B2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n687_), .A2(new_n731_), .A3(new_n587_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT47), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT44), .B1(new_n705_), .B2(new_n706_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n732_), .B1(new_n739_), .B2(new_n709_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n738_), .B(new_n735_), .C1(new_n740_), .C2(new_n731_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1330gat));
  AOI21_X1  g541(.A(G50gat), .B1(new_n687_), .B2(new_n589_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n711_), .A2(G50gat), .A3(new_n589_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n710_), .B2(new_n744_), .ZN(G1331gat));
  INV_X1    g544(.A(new_n631_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(new_n646_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n656_), .A2(new_n308_), .A3(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n511_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n607_), .A2(new_n747_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n650_), .A2(new_n360_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(G1332gat));
  OAI21_X1  g551(.A(G64gat), .B1(new_n748_), .B2(new_n663_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT48), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n663_), .A2(G64gat), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT116), .Z(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n750_), .B2(new_n756_), .ZN(G1333gat));
  OAI21_X1  g556(.A(G71gat), .B1(new_n748_), .B2(new_n588_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT49), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n588_), .A2(G71gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n750_), .B2(new_n760_), .ZN(G1334gat));
  OAI21_X1  g560(.A(G78gat), .B1(new_n748_), .B2(new_n546_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT50), .ZN(new_n763_));
  INV_X1    g562(.A(G78gat), .ZN(new_n764_));
  INV_X1    g563(.A(new_n747_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n765_), .A2(new_n546_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n607_), .A2(new_n764_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n763_), .A2(new_n767_), .ZN(G1335gat));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n704_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n704_), .A2(new_n769_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n770_), .A2(new_n307_), .A3(new_n747_), .A4(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n511_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n686_), .A2(new_n747_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n218_), .A3(new_n650_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1336gat));
  OAI21_X1  g576(.A(G92gat), .B1(new_n772_), .B2(new_n663_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n219_), .A3(new_n559_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1337gat));
  OAI21_X1  g579(.A(G99gat), .B1(new_n772_), .B2(new_n588_), .ZN(new_n781_));
  OR3_X1    g580(.A1(new_n774_), .A2(new_n215_), .A3(new_n588_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT51), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n785_), .A3(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1338gat));
  OR3_X1    g586(.A1(new_n774_), .A2(new_n216_), .A3(new_n546_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n704_), .A2(new_n307_), .A3(new_n766_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(G106gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G106gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g593(.A1(new_n610_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n616_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n614_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n614_), .A2(new_n797_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n614_), .A2(KEYINPUT118), .A3(new_n797_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT56), .B1(new_n803_), .B2(new_n623_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n801_), .A2(new_n802_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n805_), .B(new_n624_), .C1(new_n806_), .C2(new_n798_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n633_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n637_), .A2(new_n635_), .A3(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n632_), .A2(new_n808_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n645_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n638_), .B2(new_n645_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n804_), .A2(new_n807_), .A3(new_n626_), .A4(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n804_), .A2(new_n626_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(KEYINPUT58), .A3(new_n812_), .A4(new_n807_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n692_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n804_), .A2(new_n807_), .A3(new_n626_), .A4(new_n646_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n627_), .A2(new_n812_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n654_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n821_), .B2(new_n654_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n818_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n308_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n818_), .B(KEYINPUT119), .C1(new_n823_), .C2(new_n824_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n631_), .A2(new_n646_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n274_), .A2(new_n308_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT54), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n830_), .A2(KEYINPUT54), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n827_), .A2(new_n828_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n595_), .A2(new_n587_), .A3(new_n650_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n646_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n832_), .A2(new_n831_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n825_), .A2(new_n307_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  INV_X1    g639(.A(new_n834_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n835_), .B2(new_n840_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT120), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n845_), .B(new_n842_), .C1(new_n835_), .C2(new_n840_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n647_), .A2(KEYINPUT121), .ZN(new_n848_));
  MUX2_X1   g647(.A(KEYINPUT121), .B(new_n848_), .S(G113gat), .Z(new_n849_));
  AOI21_X1  g648(.A(new_n836_), .B1(new_n847_), .B2(new_n849_), .ZN(G1340gat));
  NAND2_X1  g649(.A1(new_n825_), .A2(new_n826_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n307_), .A3(new_n828_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n837_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n746_), .A2(G120gat), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n853_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n631_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G120gat), .B1(new_n856_), .B2(new_n843_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(KEYINPUT60), .B2(new_n855_), .ZN(G1341gat));
  AOI21_X1  g657(.A(G127gat), .B1(new_n835_), .B2(new_n308_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n308_), .A2(G127gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT122), .Z(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n847_), .B2(new_n861_), .ZN(G1342gat));
  AOI21_X1  g661(.A(G134gat), .B1(new_n835_), .B2(new_n655_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT123), .B(G134gat), .Z(new_n864_));
  NOR2_X1   g663(.A1(new_n274_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n847_), .B2(new_n865_), .ZN(G1343gat));
  NOR2_X1   g665(.A1(new_n546_), .A2(new_n587_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n868_), .A2(new_n511_), .A3(new_n559_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n853_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n647_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT124), .B(G141gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1344gat));
  INV_X1    g672(.A(new_n870_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n631_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g675(.A1(new_n870_), .A2(new_n307_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT61), .B(G155gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  OR3_X1    g678(.A1(new_n870_), .A2(G162gat), .A3(new_n654_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G162gat), .B1(new_n870_), .B2(new_n274_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1347gat));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n600_), .A2(new_n663_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n839_), .A2(new_n546_), .A3(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n647_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n883_), .B1(new_n886_), .B2(new_n405_), .ZN(new_n887_));
  OAI211_X1 g686(.A(KEYINPUT62), .B(G169gat), .C1(new_n885_), .C2(new_n647_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n480_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(G1348gat));
  NOR2_X1   g689(.A1(new_n833_), .A2(new_n589_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n891_), .A2(G176gat), .A3(new_n631_), .A4(new_n884_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n404_), .B1(new_n885_), .B2(new_n746_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1349gat));
  AOI211_X1 g693(.A(new_n307_), .B(new_n885_), .C1(new_n476_), .C2(new_n477_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n308_), .A3(new_n884_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n277_), .B2(new_n896_), .ZN(G1350gat));
  OAI21_X1  g696(.A(G190gat), .B1(new_n885_), .B2(new_n274_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n655_), .A2(new_n418_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n885_), .B2(new_n899_), .ZN(G1351gat));
  NOR3_X1   g699(.A1(new_n650_), .A2(new_n868_), .A3(new_n663_), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT125), .B1(new_n853_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903_));
  INV_X1    g702(.A(new_n901_), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n903_), .B(new_n904_), .C1(new_n852_), .C2(new_n837_), .ZN(new_n905_));
  OAI211_X1 g704(.A(G197gat), .B(new_n646_), .C1(new_n902_), .C2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT126), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n903_), .B1(new_n833_), .B2(new_n904_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n853_), .A2(KEYINPUT125), .A3(new_n901_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n910_), .A2(new_n911_), .A3(G197gat), .A4(new_n646_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n646_), .B1(new_n902_), .B2(new_n905_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n641_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n907_), .A2(new_n912_), .A3(new_n914_), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n910_), .A2(new_n631_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g716(.A(KEYINPUT63), .B(G211gat), .Z(new_n918_));
  OAI211_X1 g717(.A(new_n308_), .B(new_n918_), .C1(new_n902_), .C2(new_n905_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n910_), .A2(KEYINPUT127), .A3(new_n308_), .A4(new_n918_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n308_), .B1(new_n902_), .B2(new_n905_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n921_), .A2(new_n922_), .A3(new_n925_), .ZN(G1354gat));
  INV_X1    g725(.A(G218gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n910_), .A2(new_n927_), .A3(new_n655_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n274_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(G1355gat));
endmodule


