//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  XOR2_X1   g000(.A(KEYINPUT100), .B(KEYINPUT18), .Z(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT22), .B(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT84), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT23), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(G183gat), .B2(G190gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G190gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT83), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT26), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n221_), .A2(KEYINPUT83), .A3(G190gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n220_), .A2(new_n224_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT24), .A3(new_n215_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(KEYINPUT24), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n228_), .A2(new_n217_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n219_), .A2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G197gat), .B(G204gat), .Z(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(KEYINPUT21), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(KEYINPUT21), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n237_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT20), .B1(new_n234_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT95), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n241_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT97), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n211_), .B(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n215_), .B1(new_n247_), .B2(G176gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT98), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n249_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n218_), .B(KEYINPUT99), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT96), .B(KEYINPUT24), .Z(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(new_n230_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n220_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n215_), .A3(new_n230_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .A4(new_n217_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n245_), .B1(new_n253_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n210_), .B1(new_n244_), .B2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n245_), .B1(new_n219_), .B2(new_n233_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT20), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n262_), .A2(new_n263_), .A3(new_n209_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n253_), .A2(new_n245_), .A3(new_n258_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n207_), .B1(new_n261_), .B2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n242_), .B(KEYINPUT95), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(new_n259_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n206_), .B(new_n266_), .C1(new_n270_), .C2(new_n210_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT106), .B(KEYINPUT27), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT27), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n244_), .A2(new_n260_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n267_), .B1(new_n275_), .B2(new_n209_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n274_), .B1(new_n276_), .B2(new_n206_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT104), .B(KEYINPUT20), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n265_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n262_), .B1(new_n279_), .B2(KEYINPUT105), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT105), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n265_), .A2(new_n281_), .A3(new_n278_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n210_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n269_), .A2(new_n259_), .A3(new_n209_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n207_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n272_), .A2(new_n273_), .B1(new_n277_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT2), .ZN(new_n287_));
  INV_X1    g086(.A(G141gat), .ZN(new_n288_));
  INV_X1    g087(.A(G148gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n290_), .A2(new_n292_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G155gat), .B(G162gat), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT89), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G141gat), .B(G148gat), .Z(new_n300_));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(G155gat), .A3(G162gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(G155gat), .B2(G162gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n301_), .B1(G155gat), .B2(G162gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n300_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT88), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n299_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(G120gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT86), .B(G113gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n313_), .A2(KEYINPUT101), .A3(KEYINPUT4), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n308_), .A2(new_n312_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(KEYINPUT4), .A3(new_n313_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G225gat), .A2(G233gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT101), .B1(new_n313_), .B2(KEYINPUT4), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n314_), .A2(new_n316_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n315_), .A2(new_n313_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n317_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G57gat), .B(G85gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G29gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT103), .B(G1gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n323_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n320_), .A2(new_n329_), .A3(new_n322_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n308_), .A2(KEYINPUT29), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G228gat), .A2(G233gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n241_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n245_), .B1(new_n308_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT94), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G78gat), .B(G106gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n341_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n343_), .B(KEYINPUT93), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G22gat), .B(G50gat), .ZN(new_n348_));
  OR3_X1    g147(.A1(new_n308_), .A2(KEYINPUT29), .A3(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n308_), .B2(KEYINPUT29), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n345_), .A2(new_n347_), .A3(new_n352_), .A4(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n340_), .B(new_n346_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT91), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n354_), .A2(new_n357_), .A3(new_n352_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n354_), .B2(new_n352_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n356_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(KEYINPUT85), .B(KEYINPUT30), .Z(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT31), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n234_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G43gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(G71gat), .B(G99gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(new_n312_), .B(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(G15gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n368_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n366_), .B(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n286_), .A2(new_n334_), .A3(new_n362_), .A4(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n276_), .A2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n283_), .A2(new_n284_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n333_), .B(new_n377_), .C1(new_n378_), .C2(new_n376_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT33), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n332_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n332_), .A2(new_n380_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n329_), .B1(new_n321_), .B2(new_n318_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n314_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(new_n318_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n268_), .A2(new_n271_), .A3(new_n382_), .A4(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n379_), .B1(new_n381_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n362_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n333_), .B1(new_n355_), .B2(new_n360_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n286_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n373_), .B(KEYINPUT87), .Z(new_n392_));
  AOI21_X1  g191(.A(new_n375_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G15gat), .B(G22gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(KEYINPUT78), .B(G8gat), .Z(new_n395_));
  INV_X1    g194(.A(KEYINPUT14), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G1gat), .ZN(new_n398_));
  INV_X1    g197(.A(G1gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n394_), .A2(new_n396_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G8gat), .ZN(new_n402_));
  AND2_X1   g201(.A1(G231gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT68), .ZN(new_n405_));
  AND2_X1   g204(.A1(G57gat), .A2(G64gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G57gat), .A2(G64gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G57gat), .ZN(new_n409_));
  INV_X1    g208(.A(G64gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G57gat), .A2(G64gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(KEYINPUT68), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT11), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G71gat), .B(G78gat), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT69), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n408_), .A2(new_n413_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT70), .B1(new_n419_), .B2(new_n414_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n414_), .B1(new_n408_), .B2(new_n413_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT70), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT69), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n415_), .A2(new_n424_), .A3(new_n416_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n418_), .A2(new_n420_), .A3(new_n423_), .A4(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n415_), .A2(new_n424_), .A3(new_n416_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n421_), .A2(new_n422_), .ZN(new_n429_));
  AOI211_X1 g228(.A(KEYINPUT70), .B(new_n414_), .C1(new_n408_), .C2(new_n413_), .ZN(new_n430_));
  OAI22_X1  g229(.A1(new_n427_), .A2(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n404_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G127gat), .B(G155gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G211gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT16), .B(G183gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT17), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n437_), .A2(KEYINPUT79), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n438_), .B2(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n433_), .A2(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n404_), .A2(new_n432_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n404_), .A2(new_n432_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n439_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G43gat), .B(G50gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT74), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G29gat), .B(G36gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT15), .ZN(new_n451_));
  AND3_X1   g250(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G99gat), .ZN(new_n455_));
  INV_X1    g254(.A(G106gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT67), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT7), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n459_), .A2(new_n455_), .A3(new_n456_), .A4(KEYINPUT67), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n454_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G85gat), .B(G92gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT8), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n462_), .A2(KEYINPUT8), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n452_), .A2(new_n453_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT66), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n458_), .A2(new_n460_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n466_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n465_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT9), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(G85gat), .A3(G92gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n462_), .B2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT65), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT65), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n482_), .B(new_n479_), .C1(new_n462_), .C2(new_n478_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n454_), .A2(KEYINPUT66), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n467_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT10), .B(G99gat), .Z(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT64), .B(G106gat), .Z(new_n488_));
  AOI22_X1  g287(.A1(new_n485_), .A2(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n477_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n451_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G232gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT34), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n465_), .A2(new_n476_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n450_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n492_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n495_), .A2(new_n496_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n501_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G134gat), .B(G162gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT75), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G190gat), .B(G218gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT77), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n502_), .A2(new_n503_), .A3(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n502_), .A2(new_n503_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n507_), .B(KEYINPUT36), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n446_), .B(new_n511_), .C1(new_n512_), .C2(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n502_), .A2(new_n503_), .A3(new_n510_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT37), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n393_), .A2(new_n445_), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n450_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n402_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT80), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n402_), .A2(new_n522_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n402_), .A2(KEYINPUT80), .A3(new_n522_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n526_), .A2(G229gat), .A3(G233gat), .A4(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n451_), .A2(new_n402_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT81), .Z(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n523_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G113gat), .B(G141gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G197gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT82), .B(G169gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n533_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n528_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G120gat), .B(G148gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT72), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT71), .ZN(new_n545_));
  XOR2_X1   g344(.A(G176gat), .B(G204gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT5), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n545_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n498_), .A2(new_n426_), .A3(new_n431_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n426_), .A2(new_n431_), .B1(new_n477_), .B2(new_n490_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT12), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n553_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n550_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n432_), .A2(new_n491_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n498_), .A2(new_n426_), .A3(new_n431_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n550_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n549_), .B1(new_n557_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n550_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n558_), .A2(KEYINPUT12), .A3(new_n559_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n564_), .B2(new_n555_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n565_), .A2(new_n560_), .A3(new_n548_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT13), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(KEYINPUT13), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(KEYINPUT73), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT73), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n521_), .A2(new_n542_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n399_), .A3(new_n333_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT38), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n268_), .A2(new_n271_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n381_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n582_), .A2(new_n583_), .A3(new_n382_), .A4(new_n385_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n361_), .B1(new_n584_), .B2(new_n379_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n272_), .A2(new_n273_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n277_), .A2(new_n285_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n389_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n392_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n445_), .B1(new_n589_), .B2(new_n374_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n516_), .A2(new_n517_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n572_), .A2(new_n541_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G1gat), .B1(new_n594_), .B2(new_n334_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n579_), .A2(new_n580_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n581_), .A2(new_n595_), .A3(new_n596_), .ZN(G1324gat));
  OR3_X1    g396(.A1(new_n577_), .A2(new_n286_), .A3(new_n395_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n594_), .A2(new_n286_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(G8gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n599_), .B2(G8gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n598_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(KEYINPUT40), .B(new_n598_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1325gat));
  OAI21_X1  g407(.A(G15gat), .B1(new_n594_), .B2(new_n392_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT107), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT41), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n611_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT108), .ZN(new_n614_));
  INV_X1    g413(.A(new_n392_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n370_), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n577_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n614_), .B1(new_n577_), .B2(new_n616_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n612_), .A2(new_n613_), .A3(new_n617_), .A4(new_n618_), .ZN(G1326gat));
  OR3_X1    g418(.A1(new_n577_), .A2(G22gat), .A3(new_n362_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G22gat), .B1(new_n594_), .B2(new_n362_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n620_), .A2(new_n623_), .A3(new_n624_), .ZN(G1327gat));
  INV_X1    g424(.A(new_n445_), .ZN(new_n626_));
  AOI211_X1 g425(.A(new_n626_), .B(new_n592_), .C1(new_n589_), .C2(new_n374_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n593_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(G29gat), .B1(new_n629_), .B2(new_n333_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n572_), .A2(new_n626_), .A3(new_n541_), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT43), .B(new_n519_), .C1(new_n589_), .C2(new_n374_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n387_), .A2(new_n362_), .B1(new_n389_), .B2(new_n286_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n374_), .B1(new_n634_), .B2(new_n615_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n633_), .B1(new_n635_), .B2(new_n520_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n631_), .B1(new_n632_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n639_), .A2(G29gat), .A3(new_n333_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n631_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT43), .B1(new_n393_), .B2(new_n519_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n633_), .A3(new_n520_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT44), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n630_), .B1(new_n640_), .B2(new_n645_), .ZN(G1328gat));
  INV_X1    g445(.A(KEYINPUT46), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT110), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(KEYINPUT110), .ZN(new_n649_));
  INV_X1    g448(.A(G36gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n286_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(new_n645_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n586_), .A2(new_n587_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n627_), .A2(new_n650_), .A3(new_n653_), .A4(new_n593_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT45), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n648_), .B(new_n649_), .C1(new_n652_), .C2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n644_), .B2(KEYINPUT44), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n637_), .A2(new_n638_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G36gat), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n654_), .B(KEYINPUT45), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n660_), .A2(KEYINPUT110), .A3(new_n647_), .A4(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n657_), .A2(new_n662_), .ZN(G1329gat));
  INV_X1    g462(.A(G43gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n664_), .B1(new_n628_), .B2(new_n392_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n639_), .A2(G43gat), .A3(new_n373_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n659_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g467(.A(G50gat), .B1(new_n629_), .B2(new_n361_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n639_), .A2(G50gat), .A3(new_n361_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(new_n645_), .ZN(G1331gat));
  NOR2_X1   g470(.A1(new_n576_), .A2(new_n542_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n673_), .A2(new_n409_), .A3(new_n334_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n573_), .A2(new_n542_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n521_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n333_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n674_), .B1(new_n677_), .B2(new_n409_), .ZN(G1332gat));
  INV_X1    g477(.A(new_n673_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n410_), .B1(new_n679_), .B2(new_n653_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n676_), .A2(new_n410_), .A3(new_n653_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n681_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT112), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT112), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n682_), .A2(new_n683_), .A3(new_n687_), .A4(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1333gat));
  INV_X1    g488(.A(G71gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n676_), .A2(new_n690_), .A3(new_n615_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n679_), .A2(new_n615_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT49), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(G71gat), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n692_), .B2(G71gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n691_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT113), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT113), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n699_), .B(new_n691_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1334gat));
  OAI21_X1  g500(.A(G78gat), .B1(new_n673_), .B2(new_n362_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT50), .ZN(new_n703_));
  INV_X1    g502(.A(G78gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n676_), .A2(new_n704_), .A3(new_n361_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1335gat));
  INV_X1    g505(.A(KEYINPUT114), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n627_), .A2(new_n707_), .A3(new_n672_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n627_), .B2(new_n672_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n333_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n642_), .A2(new_n643_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT115), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT115), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n642_), .A2(new_n715_), .A3(new_n643_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n675_), .A2(new_n445_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n714_), .A2(new_n716_), .A3(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT116), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n333_), .A2(G85gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n712_), .B1(new_n720_), .B2(new_n721_), .ZN(G1336gat));
  AOI21_X1  g521(.A(G92gat), .B1(new_n711_), .B2(new_n653_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n653_), .A2(G92gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n720_), .B2(new_n724_), .ZN(G1337gat));
  NAND4_X1  g524(.A1(new_n714_), .A2(new_n615_), .A3(new_n716_), .A4(new_n718_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(G99gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n373_), .A2(new_n487_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n710_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT51), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n726_), .A2(G99gat), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n731_), .B(new_n732_), .C1(new_n710_), .C2(new_n728_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1338gat));
  OAI211_X1 g533(.A(new_n361_), .B(new_n488_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n717_), .A2(new_n362_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n632_), .B2(new_n636_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT117), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .A4(G106gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n456_), .B1(new_n713_), .B2(new_n736_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(new_n739_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n739_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n735_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT53), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n735_), .B(new_n746_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1339gat));
  NAND4_X1  g547(.A1(new_n539_), .A2(new_n444_), .A3(new_n441_), .A4(new_n540_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n573_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT118), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(KEYINPUT54), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(KEYINPUT54), .B2(new_n751_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n751_), .B2(KEYINPUT54), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT57), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n526_), .A2(new_n527_), .A3(new_n531_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n529_), .A2(new_n523_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n758_), .B(new_n538_), .C1(new_n759_), .C2(new_n531_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n540_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(new_n567_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT55), .B(new_n550_), .C1(new_n554_), .C2(new_n556_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT120), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT120), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n565_), .A2(new_n765_), .A3(KEYINPUT55), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT119), .B1(new_n565_), .B2(KEYINPUT55), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT119), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n557_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n564_), .A2(new_n555_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n550_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n771_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n548_), .B1(new_n768_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n779_), .A2(KEYINPUT122), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT56), .B(new_n548_), .C1(new_n768_), .C2(new_n775_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT122), .ZN(new_n783_));
  INV_X1    g582(.A(new_n780_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n776_), .A2(new_n777_), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n783_), .A3(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n541_), .A2(new_n566_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n762_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n757_), .B1(new_n788_), .B2(new_n591_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n783_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n784_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n762_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT57), .A3(new_n592_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n761_), .A2(new_n566_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n776_), .A2(new_n779_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n782_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT58), .B1(new_n799_), .B2(KEYINPUT123), .ZN(new_n800_));
  INV_X1    g599(.A(new_n782_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT55), .B1(new_n772_), .B2(new_n550_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n773_), .B1(new_n802_), .B2(new_n769_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n803_), .A2(new_n766_), .A3(new_n767_), .A4(new_n764_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n548_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n796_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT123), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n800_), .A2(new_n809_), .A3(new_n520_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n789_), .A2(new_n795_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n756_), .B1(new_n811_), .B2(new_n445_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n373_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n653_), .A2(new_n361_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n812_), .A2(new_n334_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816_), .B2(new_n542_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n591_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n810_), .B1(new_n819_), .B2(KEYINPUT57), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n788_), .A2(new_n757_), .A3(new_n591_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n445_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n756_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n334_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n818_), .B1(new_n824_), .B2(new_n814_), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n812_), .A2(KEYINPUT59), .A3(new_n334_), .A4(new_n815_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n542_), .A2(G113gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n817_), .B1(new_n827_), .B2(new_n828_), .ZN(G1340gat));
  INV_X1    g628(.A(G120gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n816_), .B(new_n831_), .C1(KEYINPUT60), .C2(new_n830_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n825_), .A2(new_n826_), .A3(new_n576_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n830_), .ZN(G1341gat));
  AOI21_X1  g633(.A(G127gat), .B1(new_n816_), .B2(new_n626_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n626_), .A2(G127gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n827_), .B2(new_n836_), .ZN(G1342gat));
  AOI21_X1  g636(.A(G134gat), .B1(new_n816_), .B2(new_n591_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n520_), .A2(G134gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n827_), .B2(new_n839_), .ZN(G1343gat));
  NOR3_X1   g639(.A1(new_n615_), .A2(new_n653_), .A3(new_n362_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n812_), .A2(new_n334_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n542_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g644(.A(new_n576_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n843_), .B2(new_n626_), .ZN(new_n852_));
  AND4_X1   g651(.A1(new_n851_), .A2(new_n824_), .A3(new_n626_), .A4(new_n841_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n850_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n824_), .A2(new_n626_), .A3(new_n841_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT124), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n843_), .A2(new_n851_), .A3(new_n626_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n849_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n858_), .ZN(G1346gat));
  AOI21_X1  g658(.A(G162gat), .B1(new_n843_), .B2(new_n591_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n520_), .A2(G162gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n843_), .B2(new_n861_), .ZN(G1347gat));
  AOI21_X1  g661(.A(new_n361_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n392_), .A2(new_n333_), .A3(new_n286_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT126), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n864_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n812_), .A2(new_n361_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT126), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n541_), .A2(new_n247_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n864_), .A2(new_n542_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n812_), .A2(new_n361_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(G169gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT62), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n822_), .A2(new_n823_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n873_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n362_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .A4(G169gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n876_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n875_), .B1(new_n863_), .B2(new_n878_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n880_), .B1(new_n884_), .B2(new_n881_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n872_), .B1(new_n883_), .B2(new_n885_), .ZN(G1348gat));
  NOR3_X1   g685(.A1(new_n865_), .A2(new_n212_), .A3(new_n576_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n867_), .A2(new_n870_), .A3(new_n572_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n212_), .ZN(G1349gat));
  AOI21_X1  g688(.A(G183gat), .B1(new_n869_), .B2(new_n626_), .ZN(new_n890_));
  AOI21_X1  g689(.A(KEYINPUT126), .B1(new_n863_), .B2(new_n864_), .ZN(new_n891_));
  NOR4_X1   g690(.A1(new_n812_), .A2(new_n866_), .A3(new_n361_), .A4(new_n868_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n445_), .A2(new_n220_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n890_), .B1(new_n893_), .B2(new_n894_), .ZN(G1350gat));
  NOR3_X1   g694(.A1(new_n891_), .A2(new_n892_), .A3(new_n519_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n867_), .A2(new_n870_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n591_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n898_));
  OAI22_X1  g697(.A1(new_n896_), .A2(new_n225_), .B1(new_n897_), .B2(new_n898_), .ZN(G1351gat));
  NAND3_X1  g698(.A1(new_n392_), .A2(new_n389_), .A3(new_n653_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n812_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n542_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n846_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n904_), .B(new_n905_), .Z(G1353gat));
  AOI21_X1  g705(.A(new_n445_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n901_), .A2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n908_), .B(new_n909_), .Z(G1354gat));
  AOI21_X1  g709(.A(G218gat), .B1(new_n901_), .B2(new_n591_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n520_), .A2(G218gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n901_), .B2(new_n912_), .ZN(G1355gat));
endmodule


