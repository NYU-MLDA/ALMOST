//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  AND3_X1   g003(.A1(KEYINPUT79), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT79), .B1(G183gat), .B2(G190gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n204_), .B1(new_n207_), .B2(new_n203_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT78), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT78), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G169gat), .A3(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n210_), .A2(new_n212_), .A3(new_n215_), .A4(KEYINPUT24), .ZN(new_n216_));
  NOR3_X1   g015(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n208_), .A2(new_n216_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n210_), .A2(new_n212_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(new_n214_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n213_), .A2(KEYINPUT22), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G169gat), .ZN(new_n229_));
  AND4_X1   g028(.A1(new_n224_), .A2(new_n227_), .A3(new_n229_), .A4(new_n214_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n223_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT79), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n202_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT79), .A2(G183gat), .A3(G190gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(KEYINPUT23), .A3(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n203_), .A2(G183gat), .A3(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(G183gat), .ZN(new_n237_));
  INV_X1    g036(.A(G190gat), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n235_), .A2(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n221_), .B1(new_n231_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT30), .ZN(new_n241_));
  XOR2_X1   g040(.A(G71gat), .B(G99gat), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G43gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(G15gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n243_), .B(new_n246_), .Z(new_n247_));
  XNOR2_X1  g046(.A(new_n241_), .B(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n248_), .A2(KEYINPUT81), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(KEYINPUT81), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G113gat), .B(G120gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT31), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(new_n250_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n254_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n248_), .A2(KEYINPUT81), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(G155gat), .A3(G162gat), .ZN(new_n260_));
  INV_X1    g059(.A(G155gat), .ZN(new_n261_));
  INV_X1    g060(.A(G162gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT1), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n262_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n260_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT82), .ZN(new_n266_));
  INV_X1    g065(.A(G141gat), .ZN(new_n267_));
  INV_X1    g066(.A(G148gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n269_), .A2(new_n270_), .B1(G141gat), .B2(G148gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT83), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n265_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n265_), .B2(new_n271_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT86), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT2), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT84), .B(KEYINPUT3), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT85), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n286_));
  NOR2_X1   g085(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n287_));
  OAI211_X1 g086(.A(KEYINPUT85), .B(new_n284_), .C1(new_n286_), .C2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n282_), .B1(new_n285_), .B2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n264_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n276_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n284_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT85), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n281_), .B1(new_n296_), .B2(new_n288_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n292_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n297_), .A2(KEYINPUT86), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n275_), .B1(new_n293_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n253_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n273_), .A2(new_n274_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n290_), .A2(new_n276_), .A3(new_n292_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT86), .B1(new_n297_), .B2(new_n298_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n253_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n302_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G1gat), .B(G29gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT0), .ZN(new_n311_));
  INV_X1    g110(.A(G57gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G85gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI211_X1 g115(.A(new_n301_), .B(new_n303_), .C1(new_n305_), .C2(new_n304_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n304_), .A2(new_n305_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n253_), .B1(new_n318_), .B2(new_n275_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT4), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n300_), .A2(new_n320_), .A3(new_n301_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n308_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n309_), .B(new_n316_), .C1(new_n321_), .C2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n302_), .A2(KEYINPUT4), .A3(new_n307_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(new_n323_), .A3(new_n322_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n316_), .B1(new_n328_), .B2(new_n309_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n258_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT28), .B1(new_n300_), .B2(KEYINPUT29), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n306_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G22gat), .B(G50gat), .Z(new_n337_));
  AND3_X1   g136(.A1(new_n333_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G228gat), .ZN(new_n342_));
  INV_X1    g141(.A(G233gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT88), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n335_), .B1(new_n318_), .B2(new_n275_), .ZN(new_n347_));
  INV_X1    g146(.A(G204gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(G197gat), .ZN(new_n349_));
  INV_X1    g148(.A(G197gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(G204gat), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT87), .B1(new_n348_), .B2(G197gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT21), .ZN(new_n354_));
  INV_X1    g153(.A(G218gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G211gat), .ZN(new_n356_));
  INV_X1    g155(.A(G211gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G218gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n352_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n361_), .A2(KEYINPUT21), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n349_), .A2(new_n351_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n363_), .A2(new_n361_), .A3(KEYINPUT21), .A4(new_n353_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n345_), .B2(new_n344_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n346_), .B1(new_n347_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n346_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n366_), .B(new_n369_), .C1(new_n306_), .C2(new_n335_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n372_), .A2(new_n373_), .A3(KEYINPUT89), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT89), .ZN(new_n375_));
  INV_X1    g174(.A(new_n371_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n300_), .A2(KEYINPUT29), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n369_), .B1(new_n377_), .B2(new_n366_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n370_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n376_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n375_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n341_), .B1(new_n374_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT89), .B1(new_n372_), .B2(new_n373_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(new_n375_), .A3(new_n381_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n340_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT27), .ZN(new_n388_));
  INV_X1    g187(.A(new_n365_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n240_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT19), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n233_), .A2(new_n203_), .A3(new_n234_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n204_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n237_), .A2(new_n238_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n227_), .A2(new_n229_), .A3(new_n214_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n223_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n235_), .A2(new_n236_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n209_), .A2(KEYINPUT24), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT90), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT90), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n209_), .A2(new_n403_), .A3(KEYINPUT24), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n215_), .A3(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n220_), .A2(new_n400_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n365_), .A2(new_n399_), .A3(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n390_), .A2(KEYINPUT20), .A3(new_n393_), .A4(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G8gat), .B(G36gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT18), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G64gat), .B(G92gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n365_), .B(new_n221_), .C1(new_n231_), .C2(new_n239_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT20), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n399_), .A2(new_n406_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n389_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT91), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT91), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n389_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n414_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n408_), .B(new_n412_), .C1(new_n420_), .C2(new_n393_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT20), .ZN(new_n423_));
  INV_X1    g222(.A(new_n239_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n398_), .A2(KEYINPUT80), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n225_), .A2(new_n224_), .A3(new_n214_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n222_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n237_), .A2(KEYINPUT25), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT25), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(G183gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n238_), .A2(KEYINPUT26), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT26), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(G190gat), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .A4(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n217_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n216_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n424_), .A2(new_n427_), .B1(new_n436_), .B2(new_n208_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n423_), .B1(new_n437_), .B2(new_n365_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n415_), .A2(new_n418_), .A3(new_n389_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n418_), .B1(new_n415_), .B2(new_n389_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n392_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n412_), .B1(new_n442_), .B2(new_n408_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n388_), .B1(new_n422_), .B2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n390_), .A2(KEYINPUT20), .A3(new_n392_), .A4(new_n407_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n420_), .B2(new_n392_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n421_), .B(KEYINPUT27), .C1(new_n446_), .C2(new_n412_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n332_), .A2(new_n387_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n386_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n328_), .A2(new_n309_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n315_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n444_), .A2(new_n452_), .A3(new_n447_), .A4(new_n325_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n340_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n450_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n412_), .A2(KEYINPUT32), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n408_), .B(new_n456_), .C1(new_n420_), .C2(new_n393_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n456_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n445_), .B(new_n458_), .C1(new_n420_), .C2(new_n392_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n457_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n460_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n462_), .B(new_n463_), .C1(new_n326_), .C2(new_n329_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n325_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n422_), .A2(new_n443_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n328_), .A2(KEYINPUT33), .A3(new_n309_), .A4(new_n316_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n327_), .A2(new_n308_), .A3(new_n322_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n302_), .A2(new_n307_), .A3(new_n323_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n315_), .A3(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .A4(new_n471_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n386_), .A2(new_n383_), .B1(new_n464_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n258_), .B1(new_n455_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT93), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n464_), .A2(new_n472_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n387_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n383_), .A2(new_n448_), .A3(new_n330_), .A4(new_n386_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n258_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n449_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G71gat), .B(G78gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n483_), .B1(KEYINPUT11), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n487_), .A2(KEYINPUT11), .A3(new_n484_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n485_), .B(KEYINPUT67), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(KEYINPUT11), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT68), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT68), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n488_), .A2(new_n494_), .A3(new_n491_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G85gat), .B(G92gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT9), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT10), .B(G99gat), .Z(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G92gat), .ZN(new_n503_));
  OR3_X1    g302(.A1(new_n314_), .A2(new_n503_), .A3(KEYINPUT9), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT6), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n499_), .A2(new_n502_), .A3(new_n504_), .A4(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT8), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n506_), .B(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n511_));
  INV_X1    g310(.A(G99gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n501_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n508_), .B1(new_n516_), .B2(new_n498_), .ZN(new_n517_));
  AOI211_X1 g316(.A(KEYINPUT8), .B(new_n497_), .C1(new_n515_), .C2(new_n506_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n507_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n496_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n496_), .A2(new_n520_), .ZN(new_n523_));
  OAI211_X1 g322(.A(G230gat), .B(G233gat), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT12), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n525_), .B1(new_n496_), .B2(new_n520_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G230gat), .A2(G233gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n492_), .A2(KEYINPUT69), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT69), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n488_), .A2(new_n529_), .A3(new_n491_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n528_), .A2(new_n519_), .A3(KEYINPUT12), .A4(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n526_), .A2(new_n527_), .A3(new_n521_), .A4(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n524_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G120gat), .B(G148gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT5), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n524_), .A2(new_n532_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT13), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT13), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n538_), .A2(new_n543_), .A3(new_n540_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G29gat), .B(G36gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G43gat), .B(G50gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n548_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n546_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G1gat), .B(G8gat), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT73), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G15gat), .B(G22gat), .ZN(new_n558_));
  INV_X1    g357(.A(G1gat), .ZN(new_n559_));
  INV_X1    g358(.A(G8gat), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT14), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n557_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n554_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n557_), .B(new_n562_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n552_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n564_), .A2(new_n552_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n571_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G169gat), .B(G197gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT77), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n574_), .A2(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n545_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n482_), .A2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n493_), .A2(new_n495_), .ZN(new_n585_));
  AND2_X1   g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n566_), .B(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n496_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G127gat), .B(G155gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n595_), .A2(KEYINPUT17), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(KEYINPUT17), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n588_), .A2(new_n590_), .A3(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT75), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n589_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n528_), .A2(new_n530_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n587_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(new_n603_), .A3(new_n596_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n605_), .B(KEYINPUT76), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n507_), .B(new_n567_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT70), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT35), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT34), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n519_), .A2(new_n554_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n609_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n613_), .A2(new_n610_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n609_), .B(new_n614_), .C1(new_n610_), .C2(new_n613_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT72), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(KEYINPUT72), .A3(new_n618_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT36), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n621_), .A2(new_n622_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT37), .ZN(new_n628_));
  INV_X1    g427(.A(new_n625_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(KEYINPUT36), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n617_), .A2(new_n630_), .A3(new_n618_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n627_), .A2(new_n628_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n626_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT37), .B1(new_n631_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT71), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT71), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n638_), .B(KEYINPUT37), .C1(new_n631_), .C2(new_n635_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n633_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n607_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n584_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n559_), .A3(new_n331_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT38), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT94), .Z(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n645_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n583_), .B(KEYINPUT95), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n627_), .A2(new_n632_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n605_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n449_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n480_), .B1(new_n479_), .B2(new_n258_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n258_), .ZN(new_n655_));
  AOI211_X1 g454(.A(KEYINPUT93), .B(new_n655_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n652_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n330_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n647_), .A2(new_n648_), .A3(new_n659_), .ZN(G1324gat));
  XNOR2_X1  g459(.A(KEYINPUT96), .B(KEYINPUT40), .ZN(new_n661_));
  INV_X1    g460(.A(new_n448_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n652_), .A2(new_n662_), .A3(new_n657_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G8gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT39), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n643_), .A2(new_n560_), .A3(new_n662_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n664_), .A2(KEYINPUT39), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n663_), .B2(G8gat), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n666_), .B(new_n661_), .C1(new_n668_), .C2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n667_), .A2(new_n672_), .ZN(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n658_), .B2(new_n258_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n643_), .A2(new_n245_), .A3(new_n655_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n676_), .A3(new_n677_), .ZN(G1326gat));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n387_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n643_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G22gat), .B1(new_n658_), .B2(new_n387_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n682_), .A2(KEYINPUT42), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(KEYINPUT42), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT97), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT97), .B(new_n681_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1327gat));
  NOR2_X1   g488(.A1(new_n606_), .A2(new_n650_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n584_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT99), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n584_), .A2(new_n693_), .A3(new_n690_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n330_), .A2(G29gat), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT100), .Z(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n482_), .A2(KEYINPUT43), .A3(new_n640_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n657_), .B2(new_n641_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n607_), .B(new_n649_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n482_), .B2(new_n640_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n657_), .A2(new_n700_), .A3(new_n641_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n707_), .A2(KEYINPUT44), .A3(new_n607_), .A4(new_n649_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n331_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT98), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(G29gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n709_), .B2(G29gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n698_), .B1(new_n711_), .B2(new_n712_), .ZN(G1328gat));
  NOR2_X1   g512(.A1(new_n448_), .A2(G36gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n692_), .A2(new_n694_), .A3(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT45), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n704_), .A2(new_n662_), .A3(new_n708_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n717_), .A2(KEYINPUT101), .A3(G36gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT101), .B1(new_n717_), .B2(G36gat), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT46), .B(new_n716_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n715_), .B(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n717_), .A2(G36gat), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n717_), .A2(KEYINPUT101), .A3(G36gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n720_), .B1(new_n727_), .B2(new_n728_), .ZN(G1329gat));
  NAND4_X1  g528(.A1(new_n704_), .A2(G43gat), .A3(new_n655_), .A4(new_n708_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n695_), .A2(new_n655_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G43gat), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g532(.A(G50gat), .B1(new_n695_), .B2(new_n680_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n704_), .A2(G50gat), .A3(new_n680_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n708_), .B2(new_n735_), .ZN(G1331gat));
  INV_X1    g535(.A(new_n582_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n545_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n642_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n482_), .B(new_n741_), .C1(new_n740_), .C2(new_n739_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n312_), .A3(new_n331_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n545_), .A2(new_n582_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n657_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n650_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n607_), .A2(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G57gat), .B1(new_n749_), .B2(new_n330_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n743_), .A2(new_n750_), .ZN(G1332gat));
  INV_X1    g550(.A(G64gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n748_), .B2(new_n662_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT48), .Z(new_n754_));
  NAND3_X1  g553(.A1(new_n742_), .A2(new_n752_), .A3(new_n662_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1333gat));
  INV_X1    g555(.A(G71gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n742_), .A2(new_n757_), .A3(new_n655_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G71gat), .B1(new_n749_), .B2(new_n258_), .ZN(new_n759_));
  XOR2_X1   g558(.A(KEYINPUT104), .B(KEYINPUT49), .Z(new_n760_));
  OR2_X1    g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n760_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(new_n761_), .A3(new_n762_), .ZN(G1334gat));
  INV_X1    g562(.A(G78gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n742_), .A2(new_n764_), .A3(new_n680_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n748_), .B2(new_n680_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n765_), .A2(new_n768_), .ZN(G1335gat));
  AND2_X1   g568(.A1(new_n745_), .A2(new_n690_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(new_n314_), .A3(new_n331_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n607_), .B(new_n744_), .C1(new_n699_), .C2(new_n701_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n772_), .A2(KEYINPUT106), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(KEYINPUT106), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n331_), .A3(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n775_), .B2(new_n314_), .ZN(G1336gat));
  NAND3_X1  g575(.A1(new_n770_), .A2(new_n503_), .A3(new_n662_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n773_), .A2(new_n662_), .A3(new_n774_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n503_), .ZN(G1337gat));
  NAND3_X1  g578(.A1(new_n770_), .A2(new_n500_), .A3(new_n655_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n772_), .A2(new_n258_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n781_), .A2(KEYINPUT107), .A3(G99gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT107), .B1(new_n781_), .B2(G99gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT51), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n786_), .B(new_n780_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1338gat));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n707_), .A2(new_n607_), .A3(new_n680_), .A4(new_n744_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(G106gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(G106gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(G106gat), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT109), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n790_), .A2(new_n791_), .A3(G106gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(KEYINPUT52), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n770_), .A2(new_n501_), .A3(new_n680_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT108), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n794_), .A2(new_n798_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT53), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n794_), .A2(new_n798_), .A3(new_n803_), .A4(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1339gat));
  INV_X1    g604(.A(G113gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n582_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n606_), .A2(new_n640_), .A3(new_n807_), .A4(new_n808_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n809_), .A2(KEYINPUT111), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(KEYINPUT111), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n606_), .A2(new_n640_), .A3(new_n807_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n808_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n573_), .A2(new_n570_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n577_), .C1(new_n570_), .C2(new_n569_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n580_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n541_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n532_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n526_), .A2(new_n521_), .A3(new_n531_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(G230gat), .A3(G233gat), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n821_), .B1(new_n532_), .B2(new_n820_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n537_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT113), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n582_), .A2(new_n540_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT113), .B(new_n537_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT56), .B1(new_n834_), .B2(KEYINPUT114), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n819_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n650_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT57), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(new_n839_), .A3(new_n650_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n818_), .A2(new_n540_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n827_), .A2(new_n829_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT56), .B(new_n537_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n844_), .A2(KEYINPUT58), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n640_), .B1(new_n844_), .B2(KEYINPUT58), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n838_), .A2(new_n840_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n815_), .B1(new_n847_), .B2(new_n651_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n680_), .A2(new_n662_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(new_n655_), .A3(new_n331_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n806_), .B1(new_n852_), .B2(new_n737_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n854_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n846_), .A2(new_n845_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n836_), .A2(new_n839_), .A3(new_n650_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n839_), .B1(new_n836_), .B2(new_n650_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(KEYINPUT116), .A3(new_n607_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT116), .B1(new_n860_), .B2(new_n607_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n815_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n850_), .A2(KEYINPUT59), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n864_), .A2(new_n865_), .B1(KEYINPUT59), .B2(new_n852_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT117), .B(G113gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n737_), .A2(new_n867_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT118), .Z(new_n869_));
  AOI22_X1  g668(.A1(new_n855_), .A2(new_n856_), .B1(new_n866_), .B2(new_n869_), .ZN(G1340gat));
  INV_X1    g669(.A(new_n852_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT119), .B(G120gat), .Z(new_n873_));
  NAND3_X1  g672(.A1(new_n738_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n852_), .A2(KEYINPUT59), .ZN(new_n877_));
  INV_X1    g676(.A(new_n815_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n847_), .B2(new_n606_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n880_), .B2(new_n861_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n865_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n877_), .B(new_n738_), .C1(new_n881_), .C2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n876_), .B1(new_n884_), .B2(new_n873_), .ZN(G1341gat));
  INV_X1    g684(.A(G127gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n871_), .A2(new_n886_), .A3(new_n606_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n877_), .B(new_n651_), .C1(new_n881_), .C2(new_n882_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n889_), .B2(new_n886_), .ZN(G1342gat));
  INV_X1    g689(.A(G134gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n640_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n866_), .A2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n852_), .B2(new_n650_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n895_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n893_), .A2(new_n896_), .A3(new_n897_), .ZN(G1343gat));
  INV_X1    g697(.A(new_n848_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n387_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n655_), .A2(new_n662_), .A3(new_n330_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n900_), .A2(new_n582_), .A3(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g702(.A1(new_n900_), .A2(new_n738_), .A3(new_n901_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT121), .B(G148gat), .Z(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1345gat));
  NAND3_X1  g705(.A1(new_n900_), .A2(new_n606_), .A3(new_n901_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT61), .B(G155gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1346gat));
  NAND2_X1  g708(.A1(new_n900_), .A2(new_n901_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G162gat), .B1(new_n910_), .B2(new_n640_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n746_), .A2(new_n262_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n910_), .B2(new_n912_), .ZN(G1347gat));
  NAND2_X1  g712(.A1(new_n332_), .A2(new_n662_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n680_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n881_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n917_), .A2(new_n582_), .A3(new_n225_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT122), .B1(new_n914_), .B2(new_n737_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n914_), .A2(KEYINPUT122), .A3(new_n737_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n680_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n864_), .A2(new_n920_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n919_), .B1(new_n923_), .B2(G169gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n920_), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n919_), .B(G169gat), .C1(new_n881_), .C2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n918_), .B1(new_n924_), .B2(new_n927_), .ZN(G1348gat));
  NOR2_X1   g727(.A1(new_n899_), .A2(new_n680_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n545_), .A2(new_n214_), .A3(new_n914_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n881_), .A2(new_n545_), .A3(new_n916_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT123), .B1(new_n932_), .B2(G176gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n864_), .A2(new_n738_), .A3(new_n915_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n934_), .A2(new_n935_), .A3(new_n214_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n931_), .B1(new_n933_), .B2(new_n936_), .ZN(G1349gat));
  NOR2_X1   g736(.A1(new_n607_), .A2(new_n914_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n929_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT124), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n848_), .A2(new_n941_), .A3(new_n387_), .A4(new_n938_), .ZN(new_n942_));
  AND2_X1   g741(.A1(new_n942_), .A2(new_n237_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n605_), .A2(new_n218_), .ZN(new_n944_));
  AOI22_X1  g743(.A1(new_n940_), .A2(new_n943_), .B1(new_n917_), .B2(new_n944_), .ZN(G1350gat));
  NAND2_X1  g744(.A1(new_n746_), .A2(new_n219_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(KEYINPUT126), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n917_), .A2(new_n947_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n864_), .A2(new_n641_), .A3(new_n915_), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n949_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(KEYINPUT125), .B1(new_n949_), .B2(G190gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n948_), .B1(new_n950_), .B2(new_n951_), .ZN(G1351gat));
  NOR3_X1   g751(.A1(new_n655_), .A2(new_n448_), .A3(new_n331_), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n848_), .A2(new_n582_), .A3(new_n680_), .A4(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(KEYINPUT127), .B1(new_n954_), .B2(new_n350_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n954_), .A2(new_n350_), .ZN(new_n956_));
  MUX2_X1   g755(.A(new_n955_), .B(KEYINPUT127), .S(new_n956_), .Z(G1352gat));
  NAND3_X1  g756(.A1(new_n900_), .A2(new_n738_), .A3(new_n953_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g758(.A1(new_n900_), .A2(new_n953_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(KEYINPUT63), .B(G211gat), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n960_), .A2(new_n651_), .A3(new_n961_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n900_), .A2(new_n953_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n963_), .A2(new_n605_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n962_), .B1(new_n964_), .B2(new_n965_), .ZN(G1354gat));
  NAND3_X1  g765(.A1(new_n960_), .A2(new_n355_), .A3(new_n746_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G218gat), .B1(new_n963_), .B2(new_n640_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(G1355gat));
endmodule


