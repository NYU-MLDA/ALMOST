//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT75), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT36), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n208_));
  NAND2_X1  g007(.A1(G232gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(KEYINPUT76), .A3(KEYINPUT35), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(KEYINPUT35), .B2(new_n210_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n217_), .A2(new_n219_), .A3(KEYINPUT66), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT66), .B1(new_n217_), .B2(new_n219_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NOR3_X1   g021(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT67), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n226_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n223_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n215_), .B1(new_n222_), .B2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n223_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(new_n227_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n214_), .B1(new_n232_), .B2(new_n213_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n235_));
  INV_X1    g034(.A(G106gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G85gat), .ZN(new_n241_));
  INV_X1    g040(.A(G92gat), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n241_), .A2(new_n242_), .A3(KEYINPUT9), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n244_));
  AND4_X1   g043(.A1(new_n240_), .A2(new_n222_), .A3(new_n243_), .A4(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n234_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G29gat), .B(G36gat), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n247_), .A2(KEYINPUT74), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(KEYINPUT74), .ZN(new_n249_));
  XOR2_X1   g048(.A(G43gat), .B(G50gat), .Z(new_n250_));
  OR3_X1    g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n212_), .B1(new_n246_), .B2(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n251_), .A2(new_n252_), .A3(KEYINPUT15), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT15), .B1(new_n251_), .B2(new_n252_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n225_), .A2(new_n227_), .ZN(new_n261_));
  OR3_X1    g060(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n218_), .B1(G99gat), .B2(G106gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n213_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT8), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n217_), .A2(new_n219_), .A3(KEYINPUT66), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n228_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n215_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n267_), .A2(KEYINPUT70), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n245_), .B1(new_n260_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n255_), .B1(new_n258_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n210_), .A2(KEYINPUT35), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT76), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n255_), .B(new_n279_), .C1(new_n258_), .C2(new_n275_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n207_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n276_), .A2(new_n280_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n205_), .B(KEYINPUT36), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(KEYINPUT77), .B(new_n207_), .C1(new_n281_), .C2(new_n283_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT37), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT78), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n287_), .A2(KEYINPUT78), .A3(new_n282_), .A4(new_n288_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n284_), .A3(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n292_), .B1(KEYINPUT37), .B2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G71gat), .B(G78gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(G57gat), .B(G64gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(KEYINPUT11), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n301_), .A3(KEYINPUT11), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n301_), .B1(new_n299_), .B2(KEYINPUT11), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n300_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT68), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(new_n298_), .A4(new_n302_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G15gat), .B(G22gat), .ZN(new_n311_));
  INV_X1    g110(.A(G1gat), .ZN(new_n312_));
  INV_X1    g111(.A(G8gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT14), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G1gat), .B(G8gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n310_), .B(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G231gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT79), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G127gat), .B(G155gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G183gat), .B(G211gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n320_), .A2(new_n321_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n322_), .A2(KEYINPUT17), .A3(new_n327_), .A4(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n327_), .B(KEYINPUT17), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT81), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n320_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n297_), .A2(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n240_), .A2(new_n222_), .A3(new_n243_), .A4(new_n244_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n229_), .A2(new_n233_), .A3(new_n259_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT70), .B1(new_n267_), .B2(new_n273_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n305_), .A2(new_n309_), .A3(KEYINPUT12), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(KEYINPUT71), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT71), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n275_), .B2(new_n340_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n267_), .A2(new_n273_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n336_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n310_), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT12), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n345_), .A2(new_n336_), .A3(new_n310_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G230gat), .A2(G233gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n352_), .B(KEYINPUT64), .Z(new_n353_));
  NOR2_X1   g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n342_), .A2(new_n344_), .A3(new_n349_), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT72), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n260_), .A2(new_n274_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n340_), .B1(new_n357_), .B2(new_n336_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n348_), .B1(new_n358_), .B2(KEYINPUT71), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n344_), .A4(new_n354_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n310_), .B1(new_n345_), .B2(new_n336_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n353_), .B1(new_n351_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(KEYINPUT69), .B(new_n353_), .C1(new_n351_), .C2(new_n362_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n356_), .A2(new_n361_), .A3(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G120gat), .B(G148gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT5), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G176gat), .B(G204gat), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n370_), .B(new_n371_), .Z(new_n372_));
  NAND2_X1  g171(.A1(new_n368_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n372_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n356_), .A2(new_n361_), .A3(new_n367_), .A4(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT13), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n373_), .A2(KEYINPUT13), .A3(new_n375_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n335_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G43gat), .ZN(new_n383_));
  INV_X1    g182(.A(G71gat), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(G99gat), .ZN(new_n385_));
  INV_X1    g184(.A(G99gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(G71gat), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n383_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n383_), .ZN(new_n390_));
  OR3_X1    g189(.A1(new_n389_), .A2(KEYINPUT31), .A3(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT31), .B1(new_n389_), .B2(new_n390_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT88), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G127gat), .B(G134gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G113gat), .B(G120gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n395_), .A2(new_n396_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n394_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n395_), .A2(new_n396_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(KEYINPUT88), .A3(new_n397_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n393_), .A2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n391_), .A2(new_n402_), .A3(new_n400_), .A4(new_n392_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT26), .B(G190gat), .ZN(new_n407_));
  INV_X1    g206(.A(G183gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT85), .B1(new_n408_), .B2(KEYINPUT25), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT25), .B(G183gat), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n407_), .B(new_n409_), .C1(new_n410_), .C2(KEYINPUT85), .ZN(new_n411_));
  INV_X1    g210(.A(G190gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT23), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT23), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(G183gat), .A3(G190gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G169gat), .ZN(new_n417_));
  INV_X1    g216(.A(G176gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G169gat), .A2(G176gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(KEYINPUT24), .A3(new_n420_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n419_), .A2(KEYINPUT24), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n411_), .A2(new_n416_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n413_), .A2(new_n424_), .A3(new_n415_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n408_), .A2(new_n412_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n414_), .A2(KEYINPUT86), .A3(G183gat), .A4(G190gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G169gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n423_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G15gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n435_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n406_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n405_), .B(new_n404_), .C1(new_n440_), .C2(new_n436_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT89), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n439_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT105), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G226gat), .A2(G233gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT19), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G197gat), .B(G204gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT21), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G218gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G211gat), .ZN(new_n454_));
  INV_X1    g253(.A(G211gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(G218gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT95), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n457_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(G197gat), .A2(G204gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G197gat), .A2(G204gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n451_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT94), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n452_), .B1(new_n460_), .B2(new_n464_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n450_), .A2(new_n451_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT94), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n466_), .B(new_n468_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n465_), .A2(new_n469_), .A3(new_n431_), .A4(new_n423_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(KEYINPUT98), .A3(KEYINPUT20), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n465_), .A2(new_n469_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n425_), .A2(new_n422_), .A3(new_n427_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n410_), .A2(new_n407_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n421_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT99), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(KEYINPUT99), .A3(new_n421_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n473_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n430_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n416_), .A2(new_n426_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT100), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n416_), .A2(KEYINPUT100), .A3(new_n426_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n480_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n472_), .B1(new_n479_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n471_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT98), .B1(new_n470_), .B2(KEYINPUT20), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n449_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G8gat), .B(G36gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G64gat), .B(G92gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n479_), .A2(new_n485_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n472_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n449_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n472_), .A2(new_n432_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n489_), .A2(new_n495_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT27), .ZN(new_n504_));
  OR3_X1    g303(.A1(new_n487_), .A2(new_n449_), .A3(new_n488_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n499_), .A2(new_n501_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n449_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n495_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n447_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n487_), .A2(new_n449_), .A3(new_n488_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n500_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n494_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n512_), .A2(KEYINPUT105), .A3(KEYINPUT27), .A4(new_n503_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G141gat), .A2(G148gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT90), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT90), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G141gat), .A3(G148gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT2), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT92), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n515_), .A2(new_n519_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT3), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(G141gat), .B2(G148gat), .ZN(new_n524_));
  INV_X1    g323(.A(G141gat), .ZN(new_n525_));
  INV_X1    g324(.A(G148gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(KEYINPUT3), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n522_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT92), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n516_), .A2(new_n518_), .A3(new_n529_), .A4(new_n519_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n521_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(G155gat), .A2(G162gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G155gat), .A2(G162gat), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT1), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(G141gat), .B2(G148gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n525_), .A2(new_n526_), .A3(KEYINPUT91), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n534_), .A2(new_n535_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n516_), .A2(new_n518_), .A3(new_n540_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n531_), .A2(new_n534_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n472_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(G228gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(G228gat), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n545_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n544_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n550_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n472_), .B(new_n552_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G78gat), .B(G106gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n551_), .A2(new_n553_), .A3(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(KEYINPUT96), .A3(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G22gat), .B(G50gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n542_), .A2(new_n562_), .A3(new_n543_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n561_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(new_n563_), .A3(new_n560_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT96), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n551_), .A2(new_n553_), .A3(new_n570_), .A4(new_n557_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n559_), .A2(new_n569_), .A3(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n558_), .A2(new_n568_), .A3(new_n566_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n557_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT97), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n566_), .A2(new_n568_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT97), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n576_), .A2(new_n556_), .A3(new_n577_), .A4(new_n558_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n572_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G1gat), .B(G29gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT103), .B(G85gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT0), .B(G57gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  AOI22_X1  g383(.A1(new_n539_), .A2(new_n541_), .B1(new_n401_), .B2(new_n397_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n531_), .A2(new_n534_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT102), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n539_), .A2(new_n541_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n403_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT102), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n585_), .A2(new_n586_), .A3(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n588_), .A2(new_n591_), .A3(KEYINPUT4), .A4(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G225gat), .A2(G233gat), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n586_), .A2(new_n589_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT4), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n588_), .A2(new_n591_), .A3(new_n593_), .A4(new_n595_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n584_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n584_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n599_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n489_), .A2(new_n502_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n494_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n503_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT27), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n606_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n514_), .A2(new_n579_), .A3(new_n611_), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT32), .B(new_n495_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n495_), .A2(KEYINPUT32), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n489_), .A2(new_n614_), .A3(new_n502_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n594_), .A2(new_n598_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(new_n603_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n613_), .B(new_n615_), .C1(new_n617_), .C2(new_n601_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n616_), .B2(new_n603_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n594_), .B(new_n595_), .C1(KEYINPUT4), .C2(new_n591_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n584_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n593_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(new_n596_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n624_), .A2(G225gat), .A3(G233gat), .A4(new_n588_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(new_n622_), .A3(new_n625_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n608_), .A2(new_n620_), .A3(new_n503_), .A4(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n599_), .A2(KEYINPUT33), .A3(new_n600_), .A4(new_n584_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n604_), .A2(KEYINPUT104), .A3(KEYINPUT33), .A4(new_n599_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n618_), .B1(new_n627_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n579_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n446_), .B1(new_n612_), .B2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n446_), .A2(new_n605_), .A3(new_n602_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n579_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n503_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n495_), .B1(new_n489_), .B2(new_n502_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n610_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n638_), .A2(new_n514_), .A3(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n636_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n253_), .A2(new_n317_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT82), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT82), .B1(new_n253_), .B2(new_n317_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n317_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(G229gat), .A2(G233gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n646_), .A2(new_n647_), .B1(new_n317_), .B2(new_n253_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n650_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G113gat), .B(G141gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT83), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G169gat), .B(G197gat), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n657_), .B(new_n658_), .Z(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n655_), .A2(KEYINPUT84), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n651_), .B(new_n660_), .C1(new_n653_), .C2(new_n650_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(KEYINPUT84), .A3(new_n663_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n643_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n382_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n606_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT38), .ZN(new_n671_));
  AOI211_X1 g470(.A(G1gat), .B(new_n669_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OAI22_X1  g472(.A1(new_n668_), .A2(new_n673_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n668_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n675_), .A2(KEYINPUT106), .A3(KEYINPUT38), .A4(new_n672_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n514_), .A2(new_n641_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n638_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n579_), .A2(new_n669_), .A3(new_n641_), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n679_), .A2(new_n514_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n680_), .B2(new_n446_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n334_), .A3(new_n296_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n378_), .A2(new_n665_), .A3(new_n379_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n378_), .A2(KEYINPUT107), .A3(new_n665_), .A4(new_n379_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n682_), .A2(new_n687_), .A3(new_n669_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n674_), .B(new_n676_), .C1(new_n312_), .C2(new_n688_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT108), .Z(G1324gat));
  INV_X1    g489(.A(new_n677_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n675_), .A2(new_n313_), .A3(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n682_), .A2(new_n687_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n691_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n682_), .A2(new_n687_), .A3(new_n677_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n313_), .B1(new_n697_), .B2(KEYINPUT109), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT39), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n696_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n692_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n702_), .B(new_n704_), .ZN(G1325gat));
  NAND2_X1  g504(.A1(new_n693_), .A2(new_n446_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G15gat), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT41), .ZN(new_n708_));
  INV_X1    g507(.A(new_n446_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n668_), .A2(G15gat), .A3(new_n709_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1326gat));
  INV_X1    g510(.A(G22gat), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n579_), .B(KEYINPUT111), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n693_), .B2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT42), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n675_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1327gat));
  INV_X1    g516(.A(KEYINPUT114), .ZN(new_n718_));
  INV_X1    g517(.A(new_n296_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n333_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n381_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n667_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(G29gat), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n606_), .A2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT113), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n685_), .A2(new_n686_), .A3(new_n333_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n643_), .B2(new_n297_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT37), .ZN(new_n732_));
  AND4_X1   g531(.A1(new_n732_), .A2(new_n294_), .A3(new_n295_), .A4(new_n284_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(KEYINPUT37), .B2(new_n291_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n731_), .B(new_n734_), .C1(new_n636_), .C2(new_n642_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n729_), .B1(new_n730_), .B2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n728_), .B1(new_n736_), .B2(KEYINPUT44), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n685_), .A2(new_n686_), .A3(new_n333_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n731_), .B1(new_n681_), .B2(new_n734_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n735_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(KEYINPUT112), .A3(new_n742_), .ZN(new_n743_));
  AOI22_X1  g542(.A1(new_n737_), .A2(new_n743_), .B1(KEYINPUT44), .B2(new_n736_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(new_n606_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n718_), .B(new_n727_), .C1(new_n745_), .C2(new_n724_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n724_), .B1(new_n744_), .B2(new_n606_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n727_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT114), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(G1328gat));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n751_));
  INV_X1    g550(.A(G36gat), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n667_), .A2(new_n721_), .A3(new_n752_), .A4(new_n691_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT115), .B(KEYINPUT45), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n677_), .B1(new_n736_), .B2(KEYINPUT44), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n736_), .A2(new_n728_), .A3(KEYINPUT44), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT112), .B1(new_n741_), .B2(new_n742_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n755_), .B1(new_n759_), .B2(G36gat), .ZN(new_n760_));
  XNOR2_X1  g559(.A(KEYINPUT116), .B(KEYINPUT46), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n751_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(KEYINPUT46), .ZN(new_n763_));
  INV_X1    g562(.A(new_n761_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n737_), .A2(new_n743_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n752_), .B1(new_n765_), .B2(new_n756_), .ZN(new_n766_));
  OAI211_X1 g565(.A(KEYINPUT117), .B(new_n764_), .C1(new_n766_), .C2(new_n755_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n762_), .A2(new_n763_), .A3(new_n767_), .ZN(G1329gat));
  AOI21_X1  g567(.A(G43gat), .B1(new_n723_), .B2(new_n446_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n709_), .A2(new_n383_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n744_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(G1330gat));
  AOI21_X1  g572(.A(G50gat), .B1(new_n723_), .B2(new_n713_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n579_), .A2(G50gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n744_), .B2(new_n775_), .ZN(G1331gat));
  NOR2_X1   g575(.A1(new_n643_), .A2(new_n719_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n380_), .A2(new_n665_), .A3(new_n333_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G57gat), .B1(new_n779_), .B2(new_n669_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n335_), .A2(new_n380_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n643_), .A2(new_n665_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n669_), .A2(G57gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT118), .Z(G1332gat));
  OAI21_X1  g585(.A(G64gat), .B1(new_n779_), .B2(new_n677_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT48), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n677_), .A2(G64gat), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT119), .Z(new_n790_));
  OAI21_X1  g589(.A(new_n788_), .B1(new_n783_), .B2(new_n790_), .ZN(G1333gat));
  OAI21_X1  g590(.A(G71gat), .B1(new_n779_), .B2(new_n709_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT49), .ZN(new_n793_));
  INV_X1    g592(.A(new_n783_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n384_), .A3(new_n446_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1334gat));
  NAND3_X1  g595(.A1(new_n777_), .A2(new_n713_), .A3(new_n778_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(G78gat), .ZN(new_n798_));
  XOR2_X1   g597(.A(KEYINPUT120), .B(KEYINPUT50), .Z(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(G78gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n801_), .A3(new_n713_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1335gat));
  NOR4_X1   g602(.A1(new_n643_), .A2(new_n380_), .A3(new_n665_), .A4(new_n720_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G85gat), .B1(new_n804_), .B2(new_n606_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n730_), .A2(new_n735_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n665_), .A2(new_n334_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n381_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n606_), .A2(G85gat), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT121), .Z(new_n811_));
  AOI21_X1  g610(.A(new_n805_), .B1(new_n809_), .B2(new_n811_), .ZN(G1336gat));
  OAI21_X1  g611(.A(G92gat), .B1(new_n808_), .B2(new_n677_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n804_), .A2(new_n242_), .A3(new_n691_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1337gat));
  OAI21_X1  g614(.A(G99gat), .B1(new_n808_), .B2(new_n709_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n804_), .A2(new_n235_), .A3(new_n237_), .A4(new_n446_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(KEYINPUT122), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n818_), .B(new_n820_), .ZN(G1338gat));
  NAND3_X1  g620(.A1(new_n804_), .A2(new_n236_), .A3(new_n579_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT123), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT52), .B(G106gat), .C1(new_n808_), .C2(new_n634_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n236_), .B1(new_n809_), .B2(new_n579_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n825_), .B(new_n826_), .C1(KEYINPUT52), .C2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(KEYINPUT52), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n823_), .A2(new_n824_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT53), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(G1339gat));
  INV_X1    g631(.A(new_n650_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n659_), .B1(new_n653_), .B2(new_n833_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n834_), .A2(KEYINPUT125), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n648_), .A2(new_n649_), .A3(new_n833_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n834_), .B2(KEYINPUT125), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n835_), .A2(new_n837_), .B1(new_n655_), .B2(new_n660_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n838_), .A2(new_n375_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n355_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n342_), .A2(new_n344_), .A3(new_n349_), .A4(new_n350_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n840_), .A2(KEYINPUT55), .B1(new_n353_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n356_), .A2(new_n843_), .A3(new_n361_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT56), .B1(new_n845_), .B2(new_n372_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT56), .ZN(new_n847_));
  AOI211_X1 g646(.A(new_n847_), .B(new_n374_), .C1(new_n842_), .C2(new_n844_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n839_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n297_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n849_), .A2(new_n850_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n665_), .B(new_n375_), .C1(new_n846_), .C2(new_n848_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n376_), .A2(new_n838_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n719_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(KEYINPUT126), .A2(KEYINPUT57), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n853_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n856_), .A2(new_n858_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n333_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n297_), .A2(new_n380_), .A3(new_n666_), .A4(new_n334_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n579_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n691_), .A2(new_n669_), .A3(new_n709_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(KEYINPUT59), .A3(new_n867_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n851_), .A2(new_n852_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n861_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n334_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n865_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n634_), .B(new_n867_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n666_), .B1(new_n868_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G113gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n665_), .A2(new_n877_), .ZN(new_n878_));
  OAI22_X1  g677(.A1(new_n876_), .A2(new_n877_), .B1(new_n873_), .B2(new_n878_), .ZN(G1340gat));
  AOI21_X1  g678(.A(new_n380_), .B1(new_n868_), .B2(new_n875_), .ZN(new_n880_));
  INV_X1    g679(.A(G120gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n380_), .B2(KEYINPUT60), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(KEYINPUT60), .B2(new_n881_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n880_), .A2(new_n881_), .B1(new_n873_), .B2(new_n883_), .ZN(G1341gat));
  AOI21_X1  g683(.A(new_n333_), .B1(new_n868_), .B2(new_n875_), .ZN(new_n885_));
  INV_X1    g684(.A(G127gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n866_), .A2(new_n334_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n867_), .A2(new_n886_), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n885_), .A2(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1342gat));
  AOI21_X1  g688(.A(new_n297_), .B1(new_n868_), .B2(new_n875_), .ZN(new_n890_));
  INV_X1    g689(.A(G134gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n719_), .A2(new_n891_), .ZN(new_n892_));
  OAI22_X1  g691(.A1(new_n890_), .A2(new_n891_), .B1(new_n873_), .B2(new_n892_), .ZN(G1343gat));
  NAND2_X1  g692(.A1(new_n862_), .A2(new_n865_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n677_), .A2(new_n606_), .A3(new_n579_), .A4(new_n709_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(KEYINPUT127), .Z(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n666_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n525_), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n380_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n526_), .ZN(G1345gat));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n333_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT61), .B(G155gat), .Z(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n897_), .B2(new_n297_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n296_), .A2(G162gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n897_), .B2(new_n906_), .ZN(G1347gat));
  INV_X1    g706(.A(KEYINPUT22), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n677_), .A2(new_n637_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n713_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n894_), .A2(new_n908_), .A3(new_n665_), .A4(new_n911_), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n912_), .A2(KEYINPUT62), .A3(new_n417_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(KEYINPUT62), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n894_), .A2(new_n665_), .A3(new_n911_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n417_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n913_), .B1(new_n914_), .B2(new_n917_), .ZN(G1348gat));
  NAND3_X1  g717(.A1(new_n894_), .A2(new_n381_), .A3(new_n911_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n910_), .A2(new_n380_), .A3(new_n418_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n919_), .A2(new_n418_), .B1(new_n866_), .B2(new_n920_), .ZN(G1349gat));
  NAND2_X1  g720(.A1(new_n894_), .A2(new_n911_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n922_), .A2(new_n333_), .A3(new_n410_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n866_), .A2(new_n334_), .A3(new_n909_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(new_n408_), .ZN(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n922_), .B2(new_n297_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n719_), .A2(new_n407_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n922_), .B2(new_n927_), .ZN(G1351gat));
  NOR4_X1   g727(.A1(new_n677_), .A2(new_n606_), .A3(new_n634_), .A4(new_n446_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n894_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n666_), .ZN(new_n931_));
  INV_X1    g730(.A(G197gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1352gat));
  NOR2_X1   g732(.A1(new_n930_), .A2(new_n380_), .ZN(new_n934_));
  INV_X1    g733(.A(G204gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1353gat));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  AND2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  NOR4_X1   g737(.A1(new_n930_), .A2(new_n333_), .A3(new_n937_), .A4(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n930_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n334_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n939_), .B1(new_n941_), .B2(new_n937_), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n930_), .B2(new_n297_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n719_), .A2(new_n453_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n930_), .B2(new_n944_), .ZN(G1355gat));
endmodule


