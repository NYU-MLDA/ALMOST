//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(G85gat), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  OR3_X1    g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT9), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n205_), .A2(new_n207_), .A3(new_n209_), .A4(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n208_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NOR3_X1   g017(.A1(KEYINPUT64), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT7), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n209_), .A2(KEYINPUT65), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n214_), .B1(new_n222_), .B2(new_n206_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n206_), .A2(new_n214_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n224_), .B1(new_n220_), .B2(new_n209_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n213_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G57gat), .B(G64gat), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n227_), .A2(KEYINPUT11), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(KEYINPUT11), .ZN(new_n229_));
  XOR2_X1   g028(.A(G71gat), .B(G78gat), .Z(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n229_), .A2(new_n230_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n226_), .A2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n233_), .B(new_n213_), .C1(new_n223_), .C2(new_n225_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT12), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT12), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n226_), .A2(new_n238_), .A3(new_n234_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G230gat), .A2(G233gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n235_), .A2(new_n243_), .A3(new_n236_), .ZN(new_n244_));
  OR3_X1    g043(.A1(new_n226_), .A2(new_n243_), .A3(new_n234_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n241_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G120gat), .B(G148gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT5), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G176gat), .B(G204gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n249_), .B(new_n250_), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n242_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(KEYINPUT67), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n253_), .B2(KEYINPUT67), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n256_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n253_), .A2(KEYINPUT67), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT68), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n262_), .B2(new_n255_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n202_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n259_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n262_), .A2(new_n258_), .A3(new_n255_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT13), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n269_), .A2(KEYINPUT69), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(KEYINPUT69), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G1gat), .B(G8gat), .Z(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT73), .B(G8gat), .ZN(new_n275_));
  INV_X1    g074(.A(G1gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT14), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT74), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n279_), .B(KEYINPUT14), .C1(new_n275_), .C2(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G15gat), .B(G22gat), .Z(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n274_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  AOI211_X1 g083(.A(new_n282_), .B(new_n273_), .C1(new_n278_), .C2(new_n280_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G29gat), .B(G36gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G43gat), .B(G50gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT75), .B1(new_n286_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n292_), .B(new_n289_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n286_), .A2(new_n290_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n295_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n298_));
  OAI211_X1 g097(.A(G229gat), .B(G233gat), .C1(new_n297_), .C2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G229gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n289_), .B(KEYINPUT15), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n286_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G113gat), .B(G141gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G169gat), .B(G197gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  NAND3_X1  g105(.A1(new_n299_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT77), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n299_), .A2(new_n303_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n306_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n314_), .A3(new_n307_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G190gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT25), .B(G183gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G190gat), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n321_), .B(new_n322_), .C1(new_n323_), .C2(new_n320_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT23), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(G183gat), .A3(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n330_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n324_), .A2(new_n329_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n325_), .A2(new_n327_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(G183gat), .ZN(new_n338_));
  INV_X1    g137(.A(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n337_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT80), .B1(G183gat), .B2(G190gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n329_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n347_));
  INV_X1    g146(.A(G176gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G169gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(G169gat), .A3(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n343_), .A2(new_n346_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n335_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(G71gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G99gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n355_), .A2(new_n360_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G15gat), .B(G43gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT30), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n365_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n367_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT31), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT31), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n369_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n363_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n375_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G127gat), .B(G134gat), .Z(new_n382_));
  XOR2_X1   g181(.A(G113gat), .B(G120gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  OR3_X1    g183(.A1(new_n380_), .A2(new_n381_), .A3(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n384_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G1gat), .B(G29gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G85gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT0), .B(G57gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n389_), .B(new_n390_), .Z(new_n391_));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(G141gat), .B(G148gat), .Z(new_n393_));
  NAND2_X1  g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT1), .ZN(new_n395_));
  INV_X1    g194(.A(G155gat), .ZN(new_n396_));
  INV_X1    g195(.A(G162gat), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(KEYINPUT83), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(G155gat), .B2(G162gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n393_), .B1(new_n395_), .B2(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n398_), .A2(new_n400_), .A3(new_n394_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n404_));
  INV_X1    g203(.A(G141gat), .ZN(new_n405_));
  INV_X1    g204(.A(G148gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G141gat), .A2(G148gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT2), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n407_), .A2(new_n410_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n403_), .A2(KEYINPUT84), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT84), .B1(new_n403_), .B2(new_n413_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n402_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n384_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n384_), .B(new_n402_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(KEYINPUT4), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n416_), .A2(new_n421_), .A3(new_n417_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n392_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n392_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n391_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n339_), .A2(KEYINPUT26), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n338_), .A2(KEYINPUT25), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT25), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G183gat), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n319_), .A2(new_n429_), .A3(new_n430_), .A4(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n334_), .A2(new_n329_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n323_), .A2(new_n322_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(KEYINPUT87), .A3(new_n334_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G211gat), .B(G218gat), .Z(new_n440_));
  INV_X1    g239(.A(KEYINPUT21), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G197gat), .B(G204gat), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(G204gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(G197gat), .ZN(new_n446_));
  INV_X1    g245(.A(G197gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(G204gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(KEYINPUT21), .B(new_n445_), .C1(new_n449_), .C2(KEYINPUT85), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n442_), .A2(new_n441_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n443_), .A2(new_n450_), .B1(new_n440_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n350_), .A2(KEYINPUT22), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT22), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G169gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT88), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n348_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(new_n341_), .A3(new_n333_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n439_), .A2(new_n452_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G226gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT19), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n442_), .A2(new_n441_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G211gat), .B(G218gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n446_), .A2(new_n448_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n445_), .A2(KEYINPUT21), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n466_), .B(new_n467_), .C1(new_n469_), .C2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n451_), .A2(new_n440_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n355_), .A2(KEYINPUT89), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT89), .B1(new_n355_), .B2(new_n473_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n461_), .B(new_n465_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n452_), .B1(new_n439_), .B2(new_n460_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT20), .B1(new_n355_), .B2(new_n473_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n463_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G8gat), .B(G36gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G64gat), .B(G92gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n476_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(KEYINPUT33), .B(new_n391_), .C1(new_n423_), .C2(new_n425_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n391_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n418_), .A2(new_n424_), .A3(new_n419_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n420_), .A2(new_n422_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n489_), .B(new_n490_), .C1(new_n491_), .C2(new_n424_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n428_), .A2(new_n487_), .A3(new_n488_), .A4(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n484_), .A2(KEYINPUT32), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n476_), .A2(new_n479_), .A3(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n437_), .A2(KEYINPUT87), .A3(new_n334_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT87), .B1(new_n437_), .B2(new_n334_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n460_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n473_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n463_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n329_), .A2(new_n345_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n326_), .A2(new_n328_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(new_n350_), .A3(new_n348_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n333_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n504_), .B1(new_n505_), .B2(new_n331_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n343_), .A2(new_n501_), .B1(new_n507_), .B2(new_n324_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n464_), .B1(new_n508_), .B2(new_n452_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n499_), .A2(new_n500_), .A3(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n471_), .A2(new_n434_), .A3(new_n472_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n341_), .A2(new_n333_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n453_), .A2(new_n455_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT88), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n512_), .B1(new_n516_), .B2(new_n348_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT20), .B1(new_n511_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n508_), .B2(new_n452_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n355_), .A2(KEYINPUT89), .A3(new_n473_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n510_), .B1(new_n522_), .B2(new_n500_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(KEYINPUT32), .A3(new_n484_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n491_), .A2(new_n424_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n425_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n489_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n423_), .A2(new_n391_), .A3(new_n425_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n495_), .B(new_n524_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n493_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G78gat), .B(G106gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G228gat), .A2(G233gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n416_), .A2(KEYINPUT29), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n533_), .B2(new_n473_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n532_), .ZN(new_n535_));
  AOI211_X1 g334(.A(new_n535_), .B(new_n452_), .C1(new_n416_), .C2(KEYINPUT29), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n531_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n416_), .A2(KEYINPUT29), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G22gat), .B(G50gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT28), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n540_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n403_), .A2(new_n413_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT84), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n403_), .A2(KEYINPUT84), .A3(new_n413_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n395_), .A2(new_n401_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n546_), .A2(new_n547_), .B1(new_n548_), .B2(new_n393_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n473_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n535_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n533_), .A2(new_n532_), .A3(new_n473_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n531_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n539_), .A2(new_n543_), .B1(new_n537_), .B2(new_n555_), .ZN(new_n556_));
  AND4_X1   g355(.A1(KEYINPUT86), .A2(new_n537_), .A3(new_n555_), .A4(new_n543_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n530_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n525_), .A2(new_n489_), .A3(new_n526_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n426_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n556_), .A2(new_n561_), .A3(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n476_), .A2(new_n479_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n484_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n476_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT27), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n484_), .B(KEYINPUT91), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT92), .B1(new_n523_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(KEYINPUT27), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n523_), .A2(KEYINPUT92), .A3(new_n568_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n567_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n562_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n387_), .B1(new_n559_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n561_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n387_), .A2(new_n558_), .A3(new_n573_), .A4(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n317_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n226_), .A2(new_n301_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT34), .Z(new_n583_));
  INV_X1    g382(.A(KEYINPUT35), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n581_), .B(new_n585_), .C1(new_n290_), .C2(new_n226_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n583_), .A2(new_n584_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n587_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n593_), .B(KEYINPUT36), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT70), .ZN(new_n597_));
  INV_X1    g396(.A(new_n590_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n588_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT71), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n595_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n589_), .A2(new_n590_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT71), .B1(new_n602_), .B2(new_n597_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT37), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(KEYINPUT72), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT72), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n602_), .A2(new_n606_), .A3(new_n597_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n605_), .A2(new_n607_), .A3(new_n608_), .A4(new_n595_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n604_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n233_), .B(new_n612_), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(new_n286_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G127gat), .B(G155gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT16), .ZN(new_n616_));
  XOR2_X1   g415(.A(G183gat), .B(G211gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n614_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n620_), .B2(new_n614_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n611_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n580_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n272_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n629_), .A2(KEYINPUT93), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(KEYINPUT93), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n561_), .B(KEYINPUT94), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n276_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n264_), .A2(new_n316_), .A3(new_n267_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT95), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT95), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n264_), .A2(new_n316_), .A3(new_n640_), .A4(new_n267_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n605_), .A2(new_n607_), .A3(new_n595_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT96), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n644_), .A2(new_n579_), .A3(new_n624_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n276_), .B1(new_n646_), .B2(new_n561_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT97), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n632_), .A2(KEYINPUT38), .A3(new_n276_), .A4(new_n634_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n637_), .A2(new_n648_), .A3(new_n649_), .ZN(G1324gat));
  INV_X1    g449(.A(new_n573_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n630_), .A2(new_n275_), .A3(new_n651_), .A4(new_n631_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n642_), .A2(new_n651_), .A3(new_n645_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G8gat), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT98), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n654_), .A2(new_n657_), .A3(G8gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n653_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n656_), .A2(new_n653_), .A3(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n652_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n652_), .B(new_n662_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1325gat));
  INV_X1    g465(.A(G15gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n646_), .B2(new_n387_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT41), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n629_), .A2(new_n667_), .A3(new_n387_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1326gat));
  OR3_X1    g470(.A1(new_n628_), .A2(G22gat), .A3(new_n558_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n558_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n646_), .A2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(G22gat), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n676_), .B2(new_n677_), .ZN(G1327gat));
  NAND3_X1  g477(.A1(new_n639_), .A2(new_n641_), .A3(new_n624_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n680_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n558_), .A2(new_n530_), .B1(new_n562_), .B2(new_n573_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT101), .B(new_n577_), .C1(new_n682_), .C2(new_n387_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n681_), .A2(new_n611_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n604_), .A2(new_n687_), .A3(new_n609_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n579_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n577_), .B1(new_n682_), .B2(new_n387_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n611_), .A2(new_n690_), .A3(KEYINPUT103), .A4(new_n687_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n685_), .A2(KEYINPUT102), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n610_), .B1(new_n690_), .B2(new_n680_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n687_), .B1(new_n693_), .B2(new_n683_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n679_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n639_), .A2(new_n641_), .A3(new_n624_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n691_), .A2(new_n689_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n685_), .A2(KEYINPUT102), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT44), .B(new_n700_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n699_), .A2(new_n634_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G29gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n643_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(new_n623_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n269_), .A2(new_n580_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OR3_X1    g509(.A1(new_n710_), .A2(G29gat), .A3(new_n576_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n706_), .A2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT105), .ZN(G1328gat));
  XNOR2_X1  g512(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n704_), .B(new_n651_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G36gat), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT106), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n715_), .A2(new_n718_), .A3(G36gat), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n710_), .A2(G36gat), .A3(new_n573_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n714_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n715_), .A2(new_n718_), .A3(G36gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n718_), .B1(new_n715_), .B2(G36gat), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n723_), .B(new_n714_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n724_), .A2(new_n728_), .ZN(G1329gat));
  NAND2_X1  g528(.A1(new_n699_), .A2(new_n704_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n387_), .A2(G43gat), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n709_), .A2(new_n387_), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n730_), .A2(new_n731_), .B1(G43gat), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n733_), .B(new_n734_), .Z(G1330gat));
  NAND2_X1  g534(.A1(new_n673_), .A2(G50gat), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n710_), .A2(new_n558_), .ZN(new_n737_));
  OAI22_X1  g536(.A1(new_n730_), .A2(new_n736_), .B1(G50gat), .B2(new_n737_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT110), .Z(G1331gat));
  AND2_X1   g538(.A1(new_n270_), .A2(new_n271_), .ZN(new_n740_));
  NOR4_X1   g539(.A1(new_n644_), .A2(new_n579_), .A3(new_n316_), .A4(new_n624_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n576_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n579_), .A2(new_n316_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n744_), .A2(new_n625_), .A3(new_n268_), .ZN(new_n745_));
  INV_X1    g544(.A(G57gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n634_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n743_), .A2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT111), .ZN(G1332gat));
  INV_X1    g548(.A(G64gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n745_), .A2(new_n750_), .A3(new_n651_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G64gat), .B1(new_n742_), .B2(new_n573_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(KEYINPUT48), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(KEYINPUT48), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(G1333gat));
  NAND3_X1  g554(.A1(new_n745_), .A2(new_n357_), .A3(new_n387_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n742_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n387_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G71gat), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT49), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT49), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n756_), .B1(new_n760_), .B2(new_n761_), .ZN(G1334gat));
  INV_X1    g561(.A(G78gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n745_), .A2(new_n763_), .A3(new_n673_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n757_), .A2(new_n673_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G78gat), .ZN(new_n767_));
  AOI211_X1 g566(.A(KEYINPUT50), .B(new_n763_), .C1(new_n757_), .C2(new_n673_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(G1335gat));
  AND2_X1   g568(.A1(new_n744_), .A2(new_n708_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n740_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n210_), .A3(new_n634_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n268_), .A2(new_n317_), .A3(new_n624_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(new_n561_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n773_), .B1(new_n210_), .B2(new_n776_), .ZN(G1336gat));
  NAND3_X1  g576(.A1(new_n772_), .A2(new_n211_), .A3(new_n651_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n775_), .A2(new_n651_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n211_), .B2(new_n779_), .ZN(G1337gat));
  AOI21_X1  g579(.A(new_n359_), .B1(new_n775_), .B2(new_n387_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n387_), .A2(new_n203_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n772_), .B2(new_n782_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g583(.A(new_n204_), .B1(new_n775_), .B2(new_n673_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n785_), .A2(KEYINPUT52), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(KEYINPUT52), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n558_), .A2(G106gat), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n771_), .A2(KEYINPUT112), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n772_), .B2(new_n788_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n786_), .B(new_n787_), .C1(new_n790_), .C2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g593(.A(new_n253_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n310_), .B2(new_n315_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n241_), .B1(new_n240_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n797_), .B2(new_n240_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n246_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT55), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT113), .B1(new_n242_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n800_), .A2(new_n804_), .A3(KEYINPUT55), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n799_), .B(new_n801_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n251_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(KEYINPUT56), .A3(new_n251_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n796_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n294_), .A2(new_n302_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n300_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n814_), .B2(new_n813_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n300_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n312_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n307_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n307_), .A3(KEYINPUT116), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n265_), .A2(new_n266_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT57), .B(new_n707_), .C1(new_n812_), .C2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n796_), .A2(new_n811_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(new_n643_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n826_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n810_), .A2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n806_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n251_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n809_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n795_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n834_), .A2(KEYINPUT58), .A3(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT58), .B1(new_n834_), .B2(new_n835_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n610_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n624_), .B1(new_n830_), .B2(new_n838_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n611_), .A2(new_n316_), .A3(new_n624_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n269_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n841_), .A2(KEYINPUT54), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(KEYINPUT54), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n844_), .ZN(new_n845_));
  AND4_X1   g644(.A1(new_n558_), .A2(new_n634_), .A3(new_n573_), .A4(new_n387_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n316_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(KEYINPUT59), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n847_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n317_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n850_), .B1(new_n854_), .B2(new_n849_), .ZN(G1340gat));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n269_), .B2(KEYINPUT60), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(KEYINPUT60), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(KEYINPUT118), .B2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n848_), .B(new_n859_), .C1(KEYINPUT118), .C2(new_n857_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n272_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n856_), .ZN(G1341gat));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n848_), .A2(new_n863_), .A3(new_n623_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n624_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n863_), .ZN(G1342gat));
  INV_X1    g665(.A(G134gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n848_), .A2(new_n867_), .A3(new_n644_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n610_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1343gat));
  NOR3_X1   g669(.A1(new_n651_), .A2(new_n558_), .A3(new_n387_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n845_), .A2(new_n634_), .A3(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n317_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n405_), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n272_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT119), .B(G148gat), .Z(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1345gat));
  NOR2_X1   g676(.A1(new_n872_), .A2(new_n624_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT61), .B(G155gat), .Z(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  OAI21_X1  g679(.A(G162gat), .B1(new_n872_), .B2(new_n610_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n644_), .A2(new_n397_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n872_), .B2(new_n882_), .ZN(G1347gat));
  OR2_X1    g682(.A1(new_n837_), .A2(new_n610_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n829_), .B(new_n826_), .C1(new_n884_), .C2(new_n836_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n885_), .A2(new_n624_), .B1(new_n843_), .B2(new_n842_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n651_), .A2(new_n633_), .A3(new_n387_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n887_), .A2(KEYINPUT120), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(KEYINPUT120), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n888_), .A2(new_n558_), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT122), .B1(new_n886_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n845_), .A2(new_n893_), .A3(new_n890_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n316_), .A3(new_n516_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n845_), .A2(new_n898_), .A3(new_n316_), .A4(new_n890_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n899_), .A2(G169gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n891_), .B1(new_n839_), .B2(new_n844_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n898_), .B1(new_n901_), .B2(new_n316_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n897_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n899_), .A2(G169gat), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n905_), .A2(KEYINPUT62), .A3(new_n902_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n896_), .B1(new_n904_), .B2(new_n906_), .ZN(G1348gat));
  NAND3_X1  g706(.A1(new_n895_), .A2(new_n348_), .A3(new_n268_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n901_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G176gat), .B1(new_n909_), .B2(new_n272_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1349gat));
  OR2_X1    g710(.A1(new_n624_), .A2(new_n322_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n901_), .A2(new_n914_), .A3(new_n623_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n338_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n901_), .B2(new_n623_), .ZN(new_n917_));
  OAI22_X1  g716(.A1(new_n913_), .A2(KEYINPUT123), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n913_), .A2(KEYINPUT123), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1350gat));
  NAND2_X1  g719(.A1(new_n644_), .A2(new_n323_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT125), .Z(new_n922_));
  NAND2_X1  g721(.A1(new_n895_), .A2(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n610_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n339_), .B2(new_n924_), .ZN(G1351gat));
  NOR4_X1   g724(.A1(new_n558_), .A2(new_n387_), .A3(new_n573_), .A4(new_n561_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n845_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n317_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(new_n447_), .ZN(G1352gat));
  INV_X1    g728(.A(new_n927_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n740_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n444_), .A2(KEYINPUT126), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n444_), .A2(KEYINPUT126), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n934_), .B1(new_n931_), .B2(new_n932_), .ZN(G1353gat));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  NOR4_X1   g736(.A1(new_n927_), .A2(new_n624_), .A3(new_n936_), .A4(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n930_), .A2(new_n623_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n939_), .B2(new_n936_), .ZN(G1354gat));
  AND3_X1   g739(.A1(new_n845_), .A2(new_n644_), .A3(new_n926_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(G218gat), .B1(new_n941_), .B2(new_n942_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n611_), .A2(G218gat), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n943_), .A2(new_n944_), .B1(new_n930_), .B2(new_n945_), .ZN(G1355gat));
endmodule


