//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n206_), .B1(G169gat), .B2(G176gat), .ZN(new_n207_));
  NOR3_X1   g006(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT23), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT79), .B1(new_n214_), .B2(KEYINPUT25), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n213_), .B(new_n215_), .C1(new_n216_), .C2(KEYINPUT79), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n211_), .B1(G183gat), .B2(G190gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(G169gat), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n212_), .A2(new_n217_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G227gat), .A2(G233gat), .ZN(new_n222_));
  INV_X1    g021(.A(G71gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n221_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G15gat), .B(G43gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT80), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT30), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n227_), .B(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n205_), .B1(new_n231_), .B2(KEYINPUT81), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(KEYINPUT81), .B2(new_n231_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n231_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n205_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT97), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G155gat), .A2(G162gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(KEYINPUT1), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(KEYINPUT1), .B2(new_n241_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT83), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n246_), .B(KEYINPUT2), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(KEYINPUT3), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(G141gat), .B2(G148gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT82), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT82), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n249_), .A2(new_n256_), .A3(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n241_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n259_), .A2(new_n240_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n248_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n260_), .ZN(new_n262_));
  AOI211_X1 g061(.A(KEYINPUT83), .B(new_n262_), .C1(new_n255_), .C2(new_n257_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n247_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n204_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n247_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n249_), .A2(new_n256_), .A3(new_n253_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n256_), .B1(new_n249_), .B2(new_n253_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n260_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT83), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n258_), .A2(new_n248_), .A3(new_n260_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n266_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n204_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n265_), .A2(new_n274_), .A3(KEYINPUT4), .ZN(new_n275_));
  OR3_X1    g074(.A1(new_n272_), .A2(KEYINPUT4), .A3(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G225gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT93), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n278_), .B(KEYINPUT94), .Z(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n276_), .A3(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n272_), .B(new_n204_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n278_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G1gat), .B(G29gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n280_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n239_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n280_), .A2(new_n282_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n287_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n280_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(KEYINPUT97), .A3(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G197gat), .B(G204gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT21), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n297_), .A2(KEYINPUT86), .A3(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G211gat), .B(G218gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n298_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n299_), .A2(new_n300_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(KEYINPUT87), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT87), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n302_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n307_), .B1(new_n308_), .B2(new_n304_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n221_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G226gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n308_), .A2(new_n304_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n218_), .A2(new_n220_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n216_), .A2(new_n213_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n209_), .A2(new_n211_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT20), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  OR3_X1    g118(.A1(new_n310_), .A2(new_n313_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n313_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n306_), .A2(new_n309_), .A3(new_n221_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT20), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n323_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT18), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n320_), .A2(new_n326_), .A3(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n310_), .A2(new_n319_), .A3(new_n313_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n330_), .B1(new_n333_), .B2(new_n325_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n313_), .B1(new_n310_), .B2(new_n319_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n322_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n332_), .B(KEYINPUT27), .C1(new_n331_), .C2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n272_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n344_), .B1(new_n272_), .B2(new_n345_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G22gat), .B(G50gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n272_), .A2(new_n345_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT28), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n349_), .B1(new_n353_), .B2(new_n346_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n351_), .A2(new_n354_), .A3(KEYINPUT84), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT84), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n350_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n353_), .A2(new_n346_), .A3(new_n349_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G78gat), .B(G106gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT90), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT89), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n272_), .B2(new_n345_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n264_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n314_), .ZN(new_n368_));
  INV_X1    g167(.A(G228gat), .ZN(new_n369_));
  INV_X1    g168(.A(G233gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT88), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT87), .B1(new_n303_), .B2(new_n305_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n308_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n375_));
  OAI22_X1  g174(.A1(new_n374_), .A2(new_n375_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n270_), .A2(new_n271_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n345_), .B1(new_n377_), .B2(new_n247_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT85), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n376_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT85), .B1(new_n272_), .B2(new_n345_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n373_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n264_), .A2(new_n379_), .A3(KEYINPUT29), .ZN(new_n383_));
  INV_X1    g182(.A(new_n376_), .ZN(new_n384_));
  AND4_X1   g183(.A1(new_n373_), .A2(new_n381_), .A3(new_n383_), .A4(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n372_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n362_), .A2(KEYINPUT90), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n364_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n381_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT88), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n381_), .A2(new_n383_), .A3(new_n384_), .A4(new_n373_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n390_), .A2(new_n391_), .B1(new_n371_), .B2(new_n368_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n387_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n360_), .B1(new_n388_), .B2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n351_), .A2(new_n354_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n362_), .A2(KEYINPUT91), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n396_), .B1(new_n386_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n397_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n392_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n296_), .B(new_n343_), .C1(new_n395_), .C2(new_n401_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n333_), .A2(new_n325_), .A3(KEYINPUT96), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n340_), .A2(new_n404_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n320_), .A2(KEYINPUT96), .A3(new_n326_), .ZN(new_n406_));
  OAI22_X1  g205(.A1(new_n403_), .A2(new_n405_), .B1(new_n406_), .B2(new_n404_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n275_), .A2(new_n278_), .A3(new_n276_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n288_), .B1(new_n281_), .B2(new_n279_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n335_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n294_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n294_), .A2(new_n412_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n408_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n357_), .A2(new_n358_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT84), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n363_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n386_), .A2(new_n387_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n417_), .B1(new_n392_), .B2(new_n399_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n386_), .A2(new_n397_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n416_), .A2(new_n421_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n238_), .B1(new_n402_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n296_), .A2(new_n238_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n421_), .A2(new_n424_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n342_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G29gat), .B(G36gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G43gat), .B(G50gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n431_), .A2(new_n433_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT15), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G15gat), .B(G22gat), .ZN(new_n439_));
  INV_X1    g238(.A(G1gat), .ZN(new_n440_));
  INV_X1    g239(.A(G8gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT14), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G1gat), .B(G8gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n438_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n437_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n447_), .A2(new_n445_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n447_), .B(new_n445_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n449_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G113gat), .B(G141gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G169gat), .B(G197gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n455_), .B(new_n456_), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n450_), .A2(new_n453_), .A3(new_n457_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n430_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n296_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT9), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(G85gat), .A3(G92gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT10), .B(G99gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G85gat), .B(G92gat), .ZN(new_n469_));
  OAI221_X1 g268(.A(new_n467_), .B1(new_n468_), .B2(G106gat), .C1(new_n466_), .C2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT64), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT6), .ZN(new_n474_));
  AND2_X1   g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n472_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n470_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n469_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n481_), .B(new_n482_), .C1(G99gat), .C2(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(G106gat), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n225_), .B(new_n484_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n480_), .B1(new_n478_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT8), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n487_), .B(new_n486_), .C1(new_n476_), .C2(new_n477_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n480_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n479_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G57gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(G64gat), .ZN(new_n496_));
  INV_X1    g295(.A(G64gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(G57gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT67), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT11), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(G57gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(G64gat), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT67), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n223_), .A2(KEYINPUT66), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT66), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G71gat), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n506_), .A2(new_n508_), .A3(G78gat), .ZN(new_n509_));
  AOI21_X1  g308(.A(G78gat), .B1(new_n506_), .B2(new_n508_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n505_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT68), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n499_), .A2(new_n504_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n514_), .B2(KEYINPUT11), .ZN(new_n515_));
  AOI211_X1 g314(.A(KEYINPUT68), .B(new_n500_), .C1(new_n499_), .C2(new_n504_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n512_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n503_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT11), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT68), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n513_), .B(KEYINPUT11), .C1(new_n518_), .C2(new_n519_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n521_), .A2(new_n505_), .A3(new_n511_), .A4(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n465_), .B1(new_n494_), .B2(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(G230gat), .A2(G233gat), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(new_n494_), .B2(new_n524_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n493_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n492_), .B1(new_n491_), .B2(new_n480_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT69), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT69), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n490_), .A2(new_n531_), .A3(new_n493_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n479_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n517_), .A2(new_n523_), .A3(KEYINPUT12), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n525_), .B(new_n527_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n494_), .A2(new_n524_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n494_), .A2(new_n524_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n526_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G120gat), .B(G148gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT5), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G176gat), .B(G204gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n535_), .A2(new_n538_), .A3(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(KEYINPUT71), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT71), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n539_), .A2(new_n548_), .A3(new_n543_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n547_), .A2(KEYINPUT13), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT13), .B1(new_n547_), .B2(new_n549_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT72), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n494_), .A2(new_n437_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n479_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT69), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n531_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n558_), .B1(new_n438_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n438_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT74), .B1(new_n533_), .B2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n563_), .A2(new_n565_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n570_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n573_), .B(new_n557_), .C1(new_n533_), .C2(new_n564_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n562_), .B2(new_n438_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n571_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n574_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT75), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n572_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n583_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT76), .Z(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n572_), .B2(new_n578_), .ZN(new_n589_));
  OR3_X1    g388(.A1(new_n585_), .A2(new_n589_), .A3(KEYINPUT37), .ZN(new_n590_));
  INV_X1    g389(.A(new_n524_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n445_), .B(new_n592_), .Z(new_n593_));
  OR2_X1    g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n593_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(G127gat), .B(G155gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT17), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n596_), .A2(new_n603_), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n594_), .B(new_n595_), .C1(new_n602_), .C2(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n606_), .A2(KEYINPUT78), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(KEYINPUT78), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT37), .B1(new_n585_), .B2(new_n589_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n590_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n556_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n463_), .A2(new_n440_), .A3(new_n464_), .A4(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND4_X1   g414(.A1(new_n461_), .A2(new_n553_), .A3(new_n555_), .A4(new_n609_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT99), .B1(new_n585_), .B2(new_n589_), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n563_), .A2(new_n573_), .B1(new_n565_), .B2(new_n571_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n533_), .A2(new_n564_), .ZN(new_n619_));
  NOR4_X1   g418(.A1(new_n619_), .A2(KEYINPUT74), .A3(new_n558_), .A4(new_n577_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n587_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n572_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n617_), .A2(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n616_), .B(new_n625_), .C1(new_n426_), .C2(new_n429_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n296_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n613_), .A2(new_n614_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n615_), .A2(new_n627_), .A3(new_n628_), .ZN(G1324gat));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631_));
  OAI21_X1  g430(.A(G8gat), .B1(new_n626_), .B2(new_n343_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(KEYINPUT39), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n386_), .A2(new_n387_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n394_), .A3(new_n363_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n635_), .A2(new_n418_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n636_), .A2(new_n343_), .A3(new_n296_), .A4(new_n238_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n342_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n638_));
  AOI22_X1  g437(.A1(new_n638_), .A2(new_n296_), .B1(new_n636_), .B2(new_n416_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n637_), .B1(new_n639_), .B2(new_n238_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n640_), .A2(new_n342_), .A3(new_n625_), .A4(new_n616_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n641_), .A2(KEYINPUT102), .A3(new_n642_), .A4(G8gat), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n633_), .A2(new_n643_), .ZN(new_n644_));
  AOI211_X1 g443(.A(KEYINPUT101), .B(new_n642_), .C1(new_n641_), .C2(G8gat), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n632_), .B2(KEYINPUT39), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n644_), .A2(new_n645_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n463_), .A2(new_n612_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n342_), .A2(new_n441_), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n649_), .A2(KEYINPUT100), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT100), .B1(new_n649_), .B2(new_n650_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n630_), .B1(new_n648_), .B2(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n645_), .A2(new_n647_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT40), .B(new_n653_), .C1(new_n656_), .C2(new_n644_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1325gat));
  NOR3_X1   g457(.A1(new_n649_), .A2(G15gat), .A3(new_n237_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT103), .Z(new_n660_));
  OAI21_X1  g459(.A(G15gat), .B1(new_n626_), .B2(new_n237_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT41), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(KEYINPUT41), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n662_), .A3(new_n663_), .ZN(G1326gat));
  XNOR2_X1  g463(.A(new_n636_), .B(KEYINPUT104), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G22gat), .B1(new_n626_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT42), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(G22gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT105), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n668_), .B1(new_n649_), .B2(new_n670_), .ZN(G1327gat));
  NOR2_X1   g470(.A1(new_n625_), .A2(new_n609_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n556_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n463_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n464_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n556_), .A2(new_n462_), .A3(new_n609_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n590_), .A2(new_n610_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n640_), .B2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n679_), .B(new_n680_), .C1(new_n426_), .C2(new_n429_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT44), .B(new_n678_), .C1(new_n681_), .C2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n678_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n680_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT43), .B1(new_n430_), .B2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n687_), .B2(new_n682_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n689_));
  OAI21_X1  g488(.A(new_n684_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n464_), .A2(G29gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n677_), .B1(new_n691_), .B2(new_n692_), .ZN(G1328gat));
  OAI211_X1 g492(.A(new_n684_), .B(new_n342_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n343_), .A2(G36gat), .ZN(new_n696_));
  OR3_X1    g495(.A1(new_n675_), .A2(KEYINPUT45), .A3(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT45), .B1(new_n675_), .B2(new_n696_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n695_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n695_), .A2(KEYINPUT46), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  NAND2_X1  g503(.A1(new_n238_), .A2(G43gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n675_), .A2(new_n237_), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n690_), .A2(new_n705_), .B1(G43gat), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g507(.A(G50gat), .B1(new_n676_), .B2(new_n665_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n428_), .A2(G50gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n691_), .B2(new_n710_), .ZN(G1331gat));
  OAI21_X1  g510(.A(KEYINPUT107), .B1(new_n430_), .B2(new_n461_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n640_), .A2(new_n713_), .A3(new_n462_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n556_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(new_n611_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n715_), .A2(KEYINPUT108), .A3(new_n717_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(new_n495_), .A3(new_n464_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n625_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n430_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n609_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n461_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n556_), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n296_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n723_), .A2(new_n729_), .ZN(G1332gat));
  NAND2_X1  g529(.A1(new_n342_), .A2(new_n497_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT109), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n722_), .A2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G64gat), .B1(new_n728_), .B2(new_n343_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1333gat));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n237_), .A2(G71gat), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n720_), .A2(new_n721_), .A3(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n725_), .A2(new_n238_), .A3(new_n556_), .A4(new_n727_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT49), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(G71gat), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n740_), .B2(G71gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n737_), .B1(new_n739_), .B2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n720_), .A2(new_n721_), .A3(new_n738_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n747_), .B(KEYINPUT110), .C1(new_n744_), .C2(new_n743_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1334gat));
  NOR2_X1   g548(.A1(new_n666_), .A2(G78gat), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n720_), .A2(new_n721_), .A3(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n725_), .A2(new_n556_), .A3(new_n665_), .A4(new_n727_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(G78gat), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n753_), .B1(new_n752_), .B2(G78gat), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT111), .B1(new_n751_), .B2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n720_), .A2(new_n721_), .A3(new_n750_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n759_), .B(new_n760_), .C1(new_n756_), .C2(new_n755_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n758_), .A2(new_n761_), .ZN(G1335gat));
  NOR3_X1   g561(.A1(new_n716_), .A2(new_n461_), .A3(new_n609_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n687_), .B2(new_n682_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n296_), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n716_), .B(new_n673_), .C1(new_n712_), .C2(new_n714_), .ZN(new_n768_));
  INV_X1    g567(.A(G85gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n464_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(G1336gat));
  AOI21_X1  g570(.A(G92gat), .B1(new_n768_), .B2(new_n342_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n342_), .A2(G92gat), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT112), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n765_), .B2(new_n774_), .ZN(G1337gat));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n237_), .A2(new_n468_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n768_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G99gat), .B1(new_n766_), .B2(new_n237_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n768_), .A2(new_n484_), .A3(new_n428_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  OAI21_X1  g583(.A(G106gat), .B1(new_n784_), .B2(KEYINPUT115), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(KEYINPUT115), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n785_), .B(new_n786_), .C1(new_n765_), .C2(new_n428_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n428_), .B(new_n763_), .C1(new_n681_), .C2(new_n683_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n785_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n788_), .A2(new_n789_), .B1(KEYINPUT115), .B2(new_n784_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n783_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n793_), .B(new_n783_), .C1(new_n787_), .C2(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1339gat));
  NAND4_X1  g594(.A1(new_n636_), .A2(new_n464_), .A3(new_n343_), .A4(new_n238_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT121), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n457_), .B1(new_n451_), .B2(new_n449_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n446_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n460_), .A2(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n547_), .A2(new_n549_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n494_), .A2(new_n524_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n525_), .B(new_n804_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n526_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n535_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n534_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n562_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n810_), .A2(KEYINPUT55), .A3(new_n525_), .A4(new_n527_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n806_), .A2(new_n808_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n543_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n543_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n461_), .A2(new_n546_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n461_), .B2(new_n546_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n803_), .B1(new_n817_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT118), .B1(new_n822_), .B2(new_n724_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n543_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n543_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n821_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n547_), .A2(new_n549_), .A3(new_n802_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n625_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n823_), .A2(new_n824_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n546_), .A2(new_n802_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n835_), .A2(KEYINPUT58), .B1(new_n590_), .B2(new_n610_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n835_), .A2(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n585_), .A2(new_n589_), .A3(KEYINPUT99), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n622_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT57), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n822_), .A2(new_n841_), .A3(KEYINPUT119), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n824_), .B1(new_n617_), .B2(new_n624_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n829_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n838_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n726_), .B1(new_n833_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n462_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n611_), .A2(new_n848_), .A3(KEYINPUT54), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT54), .B1(new_n611_), .B2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(KEYINPUT120), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n822_), .B2(new_n841_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n829_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n854_), .A2(new_n855_), .B1(new_n837_), .B2(new_n836_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n609_), .B1(new_n856_), .B2(new_n832_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n851_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n853_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n798_), .B1(new_n852_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(G113gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n461_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n847_), .A2(new_n851_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n797_), .B1(new_n864_), .B2(KEYINPUT59), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n863_), .B(new_n865_), .C1(new_n864_), .C2(new_n797_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n461_), .B(new_n866_), .C1(new_n860_), .C2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n862_), .B1(new_n869_), .B2(new_n861_), .ZN(G1340gat));
  OAI211_X1 g669(.A(new_n556_), .B(new_n866_), .C1(new_n860_), .C2(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G120gat), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT120), .B1(new_n847_), .B2(new_n851_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n857_), .A2(new_n858_), .A3(new_n853_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n797_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT123), .B1(new_n876_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n716_), .B2(KEYINPUT60), .ZN(new_n878_));
  MUX2_X1   g677(.A(KEYINPUT123), .B(new_n877_), .S(new_n878_), .Z(new_n879_));
  OAI21_X1  g678(.A(new_n872_), .B1(new_n875_), .B2(new_n879_), .ZN(G1341gat));
  INV_X1    g679(.A(G127gat), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n726_), .A2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n866_), .B(new_n882_), .C1(new_n860_), .C2(new_n867_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n609_), .B(new_n797_), .C1(new_n873_), .C2(new_n874_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT124), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n883_), .A2(new_n888_), .A3(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1342gat));
  AOI21_X1  g689(.A(G134gat), .B1(new_n860_), .B2(new_n724_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n875_), .A2(KEYINPUT59), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n892_), .A2(new_n866_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n680_), .A2(G134gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT125), .Z(new_n895_));
  AOI21_X1  g694(.A(new_n891_), .B1(new_n893_), .B2(new_n895_), .ZN(G1343gat));
  AOI21_X1  g695(.A(new_n238_), .B1(new_n852_), .B2(new_n859_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n638_), .A2(new_n464_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n897_), .A2(new_n461_), .A3(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g700(.A1(new_n897_), .A2(new_n556_), .A3(new_n899_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g702(.A1(new_n897_), .A2(new_n609_), .A3(new_n899_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1346gat));
  NAND3_X1  g705(.A1(new_n897_), .A2(new_n680_), .A3(new_n899_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G162gat), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n625_), .A2(G162gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n897_), .A2(new_n899_), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1347gat));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n427_), .A2(new_n343_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n863_), .A2(new_n666_), .A3(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n462_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT22), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n912_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G169gat), .ZN(new_n918_));
  INV_X1    g717(.A(G169gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(new_n915_), .B2(new_n912_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n918_), .B1(new_n917_), .B2(new_n920_), .ZN(G1348gat));
  AOI21_X1  g720(.A(new_n428_), .B1(new_n852_), .B2(new_n859_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n913_), .ZN(new_n923_));
  INV_X1    g722(.A(G176gat), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n716_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n665_), .B1(new_n847_), .B2(new_n851_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(new_n556_), .A3(new_n913_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n922_), .A2(new_n925_), .B1(new_n927_), .B2(new_n924_), .ZN(G1349gat));
  NOR2_X1   g727(.A1(new_n923_), .A2(new_n726_), .ZN(new_n929_));
  AOI21_X1  g728(.A(G183gat), .B1(new_n922_), .B2(new_n929_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n923_), .A2(new_n216_), .A3(new_n726_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n926_), .B2(new_n931_), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n914_), .B2(new_n686_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n926_), .A2(new_n213_), .A3(new_n724_), .A4(new_n913_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT126), .ZN(G1351gat));
  NOR3_X1   g735(.A1(new_n636_), .A2(new_n464_), .A3(new_n343_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n897_), .A2(new_n461_), .A3(new_n937_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g738(.A1(new_n897_), .A2(new_n937_), .ZN(new_n940_));
  INV_X1    g739(.A(G204gat), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n940_), .B(new_n556_), .C1(KEYINPUT127), .C2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n897_), .A2(new_n937_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n943_), .A2(new_n716_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(KEYINPUT127), .B(G204gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n942_), .B1(new_n944_), .B2(new_n945_), .ZN(G1353gat));
  XOR2_X1   g745(.A(KEYINPUT63), .B(G211gat), .Z(new_n947_));
  NAND3_X1  g746(.A1(new_n940_), .A2(new_n609_), .A3(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n949_), .B1(new_n943_), .B2(new_n726_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n948_), .A2(new_n950_), .ZN(G1354gat));
  OAI21_X1  g750(.A(G218gat), .B1(new_n943_), .B2(new_n686_), .ZN(new_n952_));
  OR2_X1    g751(.A1(new_n625_), .A2(G218gat), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n943_), .B2(new_n953_), .ZN(G1355gat));
endmodule


