//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n997_, new_n998_, new_n999_, new_n1001_, new_n1002_,
    new_n1004_, new_n1005_, new_n1006_, new_n1008_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1025_, new_n1026_, new_n1027_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n203_));
  OR2_X1    g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(KEYINPUT93), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT93), .ZN(new_n207_));
  AND2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n206_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT92), .ZN(new_n212_));
  INV_X1    g011(.A(G141gat), .ZN(new_n213_));
  INV_X1    g012(.A(G148gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT3), .ZN(new_n216_));
  AND3_X1   g015(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n212_), .A3(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n216_), .A2(new_n219_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n208_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n205_), .A2(KEYINPUT1), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n204_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(new_n220_), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n211_), .A2(new_n223_), .B1(new_n227_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n203_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n203_), .A3(new_n232_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n202_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n235_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n202_), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n238_), .A2(new_n233_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n241_), .A3(KEYINPUT99), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT99), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT97), .ZN(new_n245_));
  NAND2_X1  g044(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(KEYINPUT94), .A2(G233gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(G228gat), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n249_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n250_));
  INV_X1    g049(.A(G197gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G204gat), .ZN(new_n252_));
  INV_X1    g051(.A(G204gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G197gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT21), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT96), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n252_), .A2(new_n254_), .A3(KEYINPUT95), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT21), .B1(new_n252_), .B2(KEYINPUT95), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n253_), .A2(G197gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT95), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n258_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n252_), .A2(new_n254_), .A3(KEYINPUT95), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(KEYINPUT96), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n257_), .B1(new_n255_), .B2(KEYINPUT21), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n259_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n245_), .B1(new_n250_), .B2(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n266_), .A2(KEYINPUT96), .A3(new_n267_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT96), .B1(new_n266_), .B2(new_n267_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n271_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n259_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n206_), .A2(new_n210_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT2), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n228_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n221_), .B1(new_n220_), .B2(new_n212_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n279_), .B1(new_n222_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n227_), .A2(new_n230_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT29), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n278_), .A2(new_n289_), .A3(KEYINPUT97), .A4(new_n249_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n273_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT98), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n293_));
  OAI211_X1 g092(.A(KEYINPUT98), .B(KEYINPUT29), .C1(new_n286_), .C2(new_n288_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(new_n278_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n249_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G78gat), .B(G106gat), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n291_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n291_), .B2(new_n297_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n242_), .B(new_n244_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n291_), .A2(new_n297_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n298_), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n236_), .A2(new_n240_), .A3(new_n243_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n291_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G113gat), .B(G120gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n211_), .A2(new_n223_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n309_), .B(new_n310_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n314_), .A3(new_n287_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(KEYINPUT4), .A3(new_n315_), .ZN(new_n316_));
  OR3_X1    g115(.A1(new_n231_), .A2(KEYINPUT4), .A3(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n318_), .B(KEYINPUT102), .Z(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n312_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G85gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT0), .B(G57gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT105), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(KEYINPUT105), .A3(new_n326_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n326_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n320_), .A2(new_n321_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT19), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT101), .ZN(new_n336_));
  OR2_X1    g135(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n337_));
  NAND2_X1  g136(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT86), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n343_));
  NOR2_X1   g142(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n341_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT86), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n341_), .A2(KEYINPUT23), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n342_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G183gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT25), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G183gat), .ZN(new_n353_));
  INV_X1    g152(.A(G190gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT26), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT26), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G190gat), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n351_), .A2(new_n353_), .A3(new_n355_), .A4(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G169gat), .ZN(new_n359_));
  INV_X1    g158(.A(G176gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(KEYINPUT24), .A3(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT24), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n358_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n337_), .A2(new_n369_), .A3(new_n338_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT88), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT23), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n341_), .A2(KEYINPUT88), .A3(KEYINPUT23), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n370_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n350_), .A2(new_n354_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n360_), .A2(KEYINPUT87), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G176gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n359_), .A2(KEYINPUT22), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G169gat), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n378_), .A2(new_n380_), .A3(new_n381_), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n362_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n349_), .A2(new_n368_), .B1(new_n377_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n336_), .B1(new_n272_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n377_), .A2(new_n386_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT25), .B(G183gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT26), .B(G190gat), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n390_), .A2(new_n391_), .B1(new_n365_), .B2(new_n364_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n348_), .B1(new_n345_), .B2(KEYINPUT86), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n340_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n363_), .B(new_n392_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n389_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n278_), .A2(new_n396_), .A3(KEYINPUT101), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n388_), .A2(KEYINPUT20), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n385_), .B1(new_n349_), .B2(new_n376_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n370_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(new_n367_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT104), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n368_), .A2(new_n375_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT104), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n369_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n347_), .B1(new_n405_), .B2(new_n340_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n406_), .A2(new_n346_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n403_), .B(new_n404_), .C1(new_n407_), .C2(new_n385_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n402_), .A2(new_n408_), .A3(new_n272_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n335_), .B1(new_n398_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n272_), .B2(new_n387_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT100), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n400_), .B2(new_n367_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n392_), .A2(new_n375_), .A3(KEYINPUT100), .A4(new_n363_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n278_), .B1(new_n416_), .B2(new_n399_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n335_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n412_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n410_), .A2(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G8gat), .B(G36gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT18), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT32), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n421_), .A2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n270_), .B1(new_n263_), .B2(new_n268_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n367_), .B1(new_n346_), .B2(new_n406_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n385_), .B1(new_n376_), .B2(new_n375_), .ZN(new_n431_));
  OAI22_X1  g230(.A1(new_n429_), .A2(new_n259_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n411_), .B1(new_n432_), .B2(new_n336_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n399_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n434_), .A2(new_n272_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n433_), .A2(new_n418_), .A3(new_n397_), .A4(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n412_), .A2(new_n417_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n335_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n436_), .A2(new_n438_), .A3(KEYINPUT103), .A4(new_n426_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n426_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT103), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n333_), .A2(new_n428_), .A3(new_n439_), .A4(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n312_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n326_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT33), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n332_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n320_), .A2(new_n321_), .A3(new_n331_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT33), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n436_), .A2(new_n438_), .A3(new_n425_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n425_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n308_), .B1(new_n443_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT27), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n436_), .A2(new_n438_), .A3(new_n425_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n402_), .A2(new_n408_), .A3(new_n272_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n433_), .A2(new_n460_), .A3(new_n397_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n419_), .B1(new_n461_), .B2(new_n335_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n459_), .B(KEYINPUT27), .C1(new_n462_), .C2(new_n425_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n458_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n449_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n302_), .A2(new_n465_), .A3(new_n307_), .A4(new_n330_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468_));
  INV_X1    g267(.A(G15gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G71gat), .B(G99gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n389_), .A2(new_n395_), .A3(new_n471_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n473_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n470_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT90), .B(G43gat), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n430_), .A2(new_n431_), .A3(new_n472_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n471_), .B1(new_n389_), .B2(new_n395_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n474_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n470_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n473_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n480_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT91), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n480_), .B1(new_n479_), .B2(new_n486_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT31), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n479_), .A2(new_n486_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n480_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT31), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n493_), .A2(KEYINPUT91), .A3(new_n494_), .A4(new_n487_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n490_), .A2(new_n311_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n311_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n497_));
  OAI22_X1  g296(.A1(new_n456_), .A2(new_n467_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT106), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n490_), .A2(new_n495_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n314_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n490_), .A2(new_n311_), .A3(new_n495_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n504_), .B(KEYINPUT106), .C1(new_n456_), .C2(new_n467_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n496_), .A2(new_n497_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT107), .ZN(new_n508_));
  INV_X1    g307(.A(new_n333_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n302_), .A2(new_n307_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n510_), .A2(new_n458_), .A3(new_n463_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .A4(new_n511_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n502_), .A2(new_n509_), .A3(new_n503_), .A4(new_n511_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT107), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n506_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT7), .ZN(new_n517_));
  INV_X1    g316(.A(G99gat), .ZN(new_n518_));
  INV_X1    g317(.A(G106gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n520_), .A2(new_n523_), .A3(new_n524_), .A4(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(G85gat), .ZN(new_n527_));
  INV_X1    g326(.A(G92gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT65), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT8), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G85gat), .A2(G92gat), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n529_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n526_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT8), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(KEYINPUT65), .A3(new_n535_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n526_), .B(new_n533_), .C1(new_n530_), .C2(KEYINPUT8), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n523_), .A2(new_n524_), .ZN(new_n538_));
  OR2_X1    g337(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n519_), .A3(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n532_), .A2(KEYINPUT9), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n529_), .A2(KEYINPUT9), .A3(new_n532_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n538_), .A2(new_n541_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n536_), .A2(new_n537_), .A3(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G29gat), .B(G36gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT72), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n548_), .A2(KEYINPUT72), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n547_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n548_), .A2(KEYINPUT72), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(new_n549_), .A3(new_n546_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n552_), .A2(KEYINPUT15), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT15), .B1(new_n552_), .B2(new_n554_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n545_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n536_), .A2(new_n537_), .A3(new_n544_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n552_), .A2(new_n554_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n557_), .B2(KEYINPUT73), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n565_), .A2(KEYINPUT35), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n562_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n566_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT15), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n559_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n552_), .A2(KEYINPUT15), .A3(new_n554_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n558_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT73), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n570_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n557_), .A2(new_n561_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT74), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT36), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n569_), .A2(new_n578_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT77), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT77), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n569_), .A2(new_n578_), .A3(new_n586_), .A4(new_n583_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT75), .ZN(new_n590_));
  INV_X1    g389(.A(new_n568_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n577_), .B1(new_n576_), .B2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n562_), .A2(new_n567_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n590_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n585_), .A2(new_n587_), .A3(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n516_), .A2(KEYINPUT109), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT109), .B1(new_n516_), .B2(new_n595_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT66), .ZN(new_n599_));
  INV_X1    g398(.A(G64gat), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(G57gat), .ZN(new_n601_));
  INV_X1    g400(.A(G57gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(G64gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT11), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G71gat), .B(G78gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n599_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT11), .B1(new_n601_), .B2(new_n603_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n610_), .A2(KEYINPUT66), .A3(new_n607_), .ZN(new_n611_));
  OAI22_X1  g410(.A1(new_n609_), .A2(new_n611_), .B1(new_n605_), .B2(new_n604_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(new_n599_), .A3(new_n608_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT66), .B1(new_n610_), .B2(new_n607_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n604_), .A2(new_n605_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(new_n545_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT64), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n616_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n615_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n545_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n624_), .A2(KEYINPUT68), .A3(KEYINPUT12), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT12), .B1(new_n624_), .B2(KEYINPUT68), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n621_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT67), .B1(new_n617_), .B2(new_n545_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT67), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n558_), .A2(new_n629_), .A3(new_n616_), .A4(new_n612_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(new_n630_), .A3(new_n624_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n620_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(G120gat), .B(G148gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT70), .B1(new_n633_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT70), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n627_), .A2(new_n632_), .A3(new_n641_), .A4(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n633_), .A2(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT13), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n643_), .A2(new_n644_), .A3(KEYINPUT13), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G113gat), .B(G141gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G169gat), .B(G197gat), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n650_), .B(new_n651_), .Z(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G1gat), .B(G8gat), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT14), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT78), .B(G1gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(G8gat), .ZN(new_n658_));
  XOR2_X1   g457(.A(G15gat), .B(G22gat), .Z(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT79), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n658_), .A2(KEYINPUT79), .A3(new_n659_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n655_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n657_), .A2(G8gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n659_), .B1(new_n664_), .B2(KEYINPUT14), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT79), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n660_), .A3(new_n654_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n663_), .A2(new_n560_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(G229gat), .A2(G233gat), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n661_), .A2(new_n662_), .A3(new_n655_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n654_), .B1(new_n667_), .B2(new_n660_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n555_), .A2(new_n556_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n669_), .B(new_n670_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n670_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n671_), .A2(new_n672_), .A3(new_n559_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n560_), .B1(new_n663_), .B2(new_n668_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT83), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n559_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n669_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(KEYINPUT83), .A3(new_n677_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n676_), .B1(new_n682_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n653_), .B1(new_n686_), .B2(KEYINPUT84), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT83), .B1(new_n684_), .B2(new_n677_), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n681_), .B(new_n670_), .C1(new_n683_), .C2(new_n669_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n675_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT84), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n652_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n687_), .A2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n649_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(G231gat), .A2(G233gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n617_), .B(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(new_n673_), .ZN(new_n697_));
  XOR2_X1   g496(.A(G127gat), .B(G155gat), .Z(new_n698_));
  XNOR2_X1  g497(.A(G183gat), .B(G211gat), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT17), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n697_), .B1(KEYINPUT82), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n702_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT17), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n705_), .B(new_n708_), .C1(KEYINPUT81), .C2(new_n703_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n706_), .B1(KEYINPUT81), .B2(new_n707_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n697_), .A2(KEYINPUT82), .A3(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n694_), .A2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT108), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n598_), .A2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G1gat), .B1(new_n716_), .B2(new_n509_), .ZN(new_n717_));
  AOI22_X1  g516(.A1(new_n500_), .A2(new_n505_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT76), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n594_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT76), .B(new_n590_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n584_), .A2(KEYINPUT37), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT37), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n722_), .A2(new_n723_), .B1(new_n595_), .B2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n713_), .A2(new_n725_), .A3(new_n647_), .A4(new_n648_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n718_), .A2(new_n693_), .A3(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n509_), .A2(new_n657_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT38), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n717_), .A2(new_n730_), .ZN(G1324gat));
  INV_X1    g530(.A(G8gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n727_), .A2(new_n732_), .A3(new_n464_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n715_), .B(new_n464_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT39), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(G8gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n734_), .B2(G8gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT40), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT40), .B(new_n733_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1325gat));
  OAI21_X1  g541(.A(G15gat), .B1(new_n716_), .B2(new_n504_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT41), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT41), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n745_), .B(G15gat), .C1(new_n716_), .C2(new_n504_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n727_), .A2(new_n469_), .A3(new_n507_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT110), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n744_), .A2(new_n746_), .A3(new_n748_), .ZN(G1326gat));
  INV_X1    g548(.A(G22gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n727_), .A2(new_n750_), .A3(new_n308_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n598_), .A2(new_n308_), .A3(new_n715_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G22gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G22gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(G1327gat));
  NAND2_X1  g555(.A1(new_n694_), .A2(new_n712_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n718_), .B2(new_n725_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n759_));
  INV_X1    g558(.A(new_n725_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n516_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n757_), .B1(new_n758_), .B2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(G29gat), .B(new_n333_), .C1(new_n762_), .C2(KEYINPUT44), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n764_), .B(new_n757_), .C1(new_n758_), .C2(new_n761_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n718_), .A2(new_n693_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n649_), .A2(new_n713_), .A3(new_n595_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(new_n509_), .ZN(new_n769_));
  OAI22_X1  g568(.A1(new_n763_), .A2(new_n765_), .B1(G29gat), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT111), .ZN(G1328gat));
  OAI21_X1  g570(.A(new_n464_), .B1(new_n762_), .B2(KEYINPUT44), .ZN(new_n772_));
  OAI21_X1  g571(.A(G36gat), .B1(new_n772_), .B2(new_n765_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n464_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(G36gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n766_), .A2(new_n767_), .A3(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT45), .ZN(new_n777_));
  XNOR2_X1  g576(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n773_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1329gat));
  INV_X1    g580(.A(new_n693_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n516_), .A2(new_n507_), .A3(new_n782_), .A4(new_n767_), .ZN(new_n783_));
  INV_X1    g582(.A(G43gat), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(G43gat), .B(new_n507_), .C1(new_n762_), .C2(KEYINPUT44), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n765_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT47), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n787_), .B(new_n791_), .C1(new_n765_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1330gat));
  INV_X1    g592(.A(new_n768_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G50gat), .B1(new_n794_), .B2(new_n308_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n762_), .A2(KEYINPUT44), .ZN(new_n796_));
  INV_X1    g595(.A(G50gat), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n510_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n765_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(G1331gat));
  INV_X1    g599(.A(new_n649_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(new_n782_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n713_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT114), .B(new_n804_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n509_), .A2(new_n602_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n810_), .A2(KEYINPUT115), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(KEYINPUT115), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n516_), .A2(new_n802_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n760_), .A2(new_n712_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G57gat), .B1(new_n816_), .B2(new_n333_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n811_), .A2(new_n812_), .A3(new_n817_), .ZN(G1332gat));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n600_), .A3(new_n464_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n807_), .A2(new_n464_), .A3(new_n808_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT48), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n820_), .A2(new_n821_), .A3(G64gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n820_), .B2(G64gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n819_), .B1(new_n822_), .B2(new_n823_), .ZN(G1333gat));
  OR3_X1    g623(.A1(new_n815_), .A2(G71gat), .A3(new_n504_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n807_), .A2(new_n507_), .A3(new_n808_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n826_), .A2(new_n827_), .A3(G71gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n826_), .B2(G71gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n828_), .B2(new_n829_), .ZN(G1334gat));
  OR3_X1    g629(.A1(new_n815_), .A2(G78gat), .A3(new_n510_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n807_), .A2(new_n308_), .A3(new_n808_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(G78gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(G78gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(G1335gat));
  AOI21_X1  g635(.A(new_n759_), .B1(new_n516_), .B2(new_n760_), .ZN(new_n837_));
  AOI211_X1 g636(.A(KEYINPUT43), .B(new_n725_), .C1(new_n506_), .C2(new_n515_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT116), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n758_), .A2(new_n761_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n802_), .A2(new_n712_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n839_), .A2(new_n841_), .A3(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(G85gat), .B1(new_n844_), .B2(new_n509_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n595_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n813_), .A2(new_n846_), .A3(new_n712_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n527_), .A3(new_n333_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(G1336gat));
  OAI21_X1  g648(.A(G92gat), .B1(new_n844_), .B2(new_n774_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n528_), .A3(new_n464_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1337gat));
  OAI21_X1  g651(.A(G99gat), .B1(new_n844_), .B2(new_n504_), .ZN(new_n853_));
  OR2_X1    g652(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n507_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n847_), .A2(new_n855_), .B1(KEYINPUT117), .B2(KEYINPUT51), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n853_), .A2(new_n854_), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n854_), .B1(new_n853_), .B2(new_n856_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1338gat));
  NAND2_X1  g658(.A1(new_n843_), .A2(new_n308_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n758_), .B2(new_n761_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT118), .B1(new_n861_), .B2(new_n519_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n842_), .A2(new_n510_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(G106gat), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n862_), .A2(new_n866_), .A3(KEYINPUT52), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT118), .B(new_n868_), .C1(new_n861_), .C2(new_n519_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n847_), .A2(new_n519_), .A3(new_n308_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT53), .B1(new_n867_), .B2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n862_), .A2(new_n866_), .A3(KEYINPUT52), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n870_), .A4(new_n869_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(G1339gat));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n684_), .A2(new_n670_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n669_), .B(new_n677_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n653_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n690_), .A2(new_n652_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n643_), .A2(new_n644_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n625_), .A2(new_n626_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n628_), .A2(new_n630_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n620_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT55), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n627_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n621_), .B(KEYINPUT55), .C1(new_n625_), .C2(new_n626_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n639_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(KEYINPUT56), .A3(new_n639_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n643_), .A2(new_n687_), .A3(new_n692_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n883_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n877_), .B1(new_n897_), .B2(new_n846_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n882_), .A2(new_n881_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n890_), .A2(KEYINPUT56), .A3(new_n639_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n890_), .B2(new_n639_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n643_), .B(new_n899_), .C1(new_n900_), .C2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n895_), .A2(KEYINPUT58), .A3(new_n643_), .A4(new_n899_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(new_n905_), .A3(new_n760_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n643_), .A2(new_n687_), .A3(new_n692_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n908_));
  OAI211_X1 g707(.A(KEYINPUT57), .B(new_n595_), .C1(new_n908_), .C2(new_n883_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n898_), .A2(new_n906_), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n712_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n814_), .A2(new_n913_), .A3(new_n801_), .A4(new_n693_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT54), .B1(new_n726_), .B2(new_n782_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n911_), .A2(new_n912_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n912_), .B1(new_n911_), .B2(new_n916_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n507_), .A2(new_n333_), .A3(new_n511_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(G113gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n921_), .A2(new_n922_), .A3(new_n782_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n924_));
  INV_X1    g723(.A(new_n909_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n898_), .A2(new_n906_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n595_), .B1(new_n908_), .B2(new_n883_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n725_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n929_), .A2(new_n877_), .B1(new_n930_), .B2(new_n905_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT121), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n713_), .B1(new_n928_), .B2(new_n932_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n914_), .A2(new_n915_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n920_), .B(KEYINPUT120), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n924_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n919_), .A2(KEYINPUT59), .A3(new_n920_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n693_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n923_), .B1(new_n939_), .B2(new_n922_), .ZN(G1340gat));
  INV_X1    g739(.A(G120gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n941_), .B1(new_n801_), .B2(KEYINPUT60), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n921_), .B(new_n942_), .C1(KEYINPUT60), .C2(new_n941_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n801_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n944_), .B2(new_n941_), .ZN(G1341gat));
  INV_X1    g744(.A(G127gat), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n921_), .A2(new_n946_), .A3(new_n713_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n712_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n946_), .ZN(G1342gat));
  INV_X1    g748(.A(G134gat), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n921_), .A2(new_n950_), .A3(new_n846_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n725_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n952_), .B2(new_n950_), .ZN(G1343gat));
  AOI21_X1  g752(.A(new_n713_), .B1(new_n931_), .B2(new_n909_), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT119), .B1(new_n954_), .B2(new_n934_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n911_), .A2(new_n912_), .A3(new_n916_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n464_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n957_));
  NAND4_X1  g756(.A1(new_n955_), .A2(new_n504_), .A3(new_n956_), .A4(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n958_), .A2(new_n693_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(new_n213_), .ZN(G1344gat));
  NOR2_X1   g759(.A1(new_n958_), .A2(new_n801_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(new_n214_), .ZN(G1345gat));
  NOR3_X1   g761(.A1(new_n917_), .A2(new_n918_), .A3(new_n507_), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n963_), .A2(KEYINPUT122), .A3(new_n713_), .A4(new_n957_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n965_), .B1(new_n958_), .B2(new_n712_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(KEYINPUT61), .B(G155gat), .ZN(new_n967_));
  AND3_X1   g766(.A1(new_n964_), .A2(new_n966_), .A3(new_n967_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n967_), .B1(new_n964_), .B2(new_n966_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1346gat));
  OAI21_X1  g769(.A(G162gat), .B1(new_n958_), .B2(new_n725_), .ZN(new_n971_));
  OR2_X1    g770(.A1(new_n595_), .A2(G162gat), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n958_), .B2(new_n972_), .ZN(G1347gat));
  NAND3_X1  g772(.A1(new_n507_), .A2(new_n509_), .A3(new_n464_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n974_), .A2(new_n308_), .ZN(new_n975_));
  OAI211_X1 g774(.A(new_n782_), .B(new_n975_), .C1(new_n933_), .C2(new_n934_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n976_), .A2(KEYINPUT123), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n909_), .B1(new_n931_), .B2(KEYINPUT121), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n926_), .A2(new_n927_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n712_), .B1(new_n978_), .B2(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n980_), .A2(new_n916_), .ZN(new_n981_));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n982_));
  NAND4_X1  g781(.A1(new_n981_), .A2(new_n982_), .A3(new_n782_), .A4(new_n975_), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n977_), .A2(new_n983_), .A3(G169gat), .ZN(new_n984_));
  XNOR2_X1  g783(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(new_n986_));
  AND2_X1   g785(.A1(new_n981_), .A2(new_n975_), .ZN(new_n987_));
  NAND4_X1  g786(.A1(new_n987_), .A2(new_n381_), .A3(new_n383_), .A4(new_n782_), .ZN(new_n988_));
  INV_X1    g787(.A(new_n985_), .ZN(new_n989_));
  NAND4_X1  g788(.A1(new_n977_), .A2(new_n983_), .A3(G169gat), .A4(new_n989_), .ZN(new_n990_));
  NAND3_X1  g789(.A1(new_n986_), .A2(new_n988_), .A3(new_n990_), .ZN(G1348gat));
  NAND2_X1  g790(.A1(new_n987_), .A2(new_n649_), .ZN(new_n992_));
  AND2_X1   g791(.A1(new_n378_), .A2(new_n380_), .ZN(new_n993_));
  NOR3_X1   g792(.A1(new_n917_), .A2(new_n918_), .A3(new_n308_), .ZN(new_n994_));
  NOR3_X1   g793(.A1(new_n974_), .A2(new_n801_), .A3(new_n360_), .ZN(new_n995_));
  AOI22_X1  g794(.A1(new_n992_), .A2(new_n993_), .B1(new_n994_), .B2(new_n995_), .ZN(G1349gat));
  NOR2_X1   g795(.A1(new_n974_), .A2(new_n712_), .ZN(new_n997_));
  AOI21_X1  g796(.A(G183gat), .B1(new_n994_), .B2(new_n997_), .ZN(new_n998_));
  NOR2_X1   g797(.A1(new_n712_), .A2(new_n390_), .ZN(new_n999_));
  AOI21_X1  g798(.A(new_n998_), .B1(new_n987_), .B2(new_n999_), .ZN(G1350gat));
  NAND3_X1  g799(.A1(new_n987_), .A2(new_n391_), .A3(new_n846_), .ZN(new_n1001_));
  AND2_X1   g800(.A1(new_n987_), .A2(new_n760_), .ZN(new_n1002_));
  OAI21_X1  g801(.A(new_n1001_), .B1(new_n1002_), .B2(new_n354_), .ZN(G1351gat));
  NOR2_X1   g802(.A1(new_n774_), .A2(new_n466_), .ZN(new_n1004_));
  NAND4_X1  g803(.A1(new_n955_), .A2(new_n504_), .A3(new_n956_), .A4(new_n1004_), .ZN(new_n1005_));
  NOR2_X1   g804(.A1(new_n1005_), .A2(new_n693_), .ZN(new_n1006_));
  XNOR2_X1  g805(.A(new_n1006_), .B(new_n251_), .ZN(G1352gat));
  NOR2_X1   g806(.A1(new_n1005_), .A2(new_n801_), .ZN(new_n1008_));
  XNOR2_X1  g807(.A(new_n1008_), .B(new_n253_), .ZN(G1353gat));
  NOR2_X1   g808(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1010_));
  INV_X1    g809(.A(new_n1010_), .ZN(new_n1011_));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n1012_));
  INV_X1    g811(.A(new_n1005_), .ZN(new_n1013_));
  NAND2_X1  g812(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1014_));
  NAND2_X1  g813(.A1(new_n713_), .A2(new_n1014_), .ZN(new_n1015_));
  XNOR2_X1  g814(.A(new_n1015_), .B(KEYINPUT125), .ZN(new_n1016_));
  INV_X1    g815(.A(new_n1016_), .ZN(new_n1017_));
  AOI21_X1  g816(.A(new_n1012_), .B1(new_n1013_), .B2(new_n1017_), .ZN(new_n1018_));
  NOR3_X1   g817(.A1(new_n1005_), .A2(KEYINPUT126), .A3(new_n1016_), .ZN(new_n1019_));
  OAI21_X1  g818(.A(new_n1011_), .B1(new_n1018_), .B2(new_n1019_), .ZN(new_n1020_));
  NAND3_X1  g819(.A1(new_n1013_), .A2(new_n1012_), .A3(new_n1017_), .ZN(new_n1021_));
  OAI21_X1  g820(.A(KEYINPUT126), .B1(new_n1005_), .B2(new_n1016_), .ZN(new_n1022_));
  NAND3_X1  g821(.A1(new_n1021_), .A2(new_n1010_), .A3(new_n1022_), .ZN(new_n1023_));
  NAND2_X1  g822(.A1(new_n1020_), .A2(new_n1023_), .ZN(G1354gat));
  XNOR2_X1  g823(.A(KEYINPUT127), .B(G218gat), .ZN(new_n1025_));
  NOR3_X1   g824(.A1(new_n1005_), .A2(new_n725_), .A3(new_n1025_), .ZN(new_n1026_));
  NAND2_X1  g825(.A1(new_n1013_), .A2(new_n846_), .ZN(new_n1027_));
  AOI21_X1  g826(.A(new_n1026_), .B1(new_n1027_), .B2(new_n1025_), .ZN(G1355gat));
endmodule


