//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_;
  INV_X1    g000(.A(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT7), .ZN(new_n205_));
  OAI211_X1 g004(.A(new_n202_), .B(new_n203_), .C1(new_n204_), .C2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(KEYINPUT64), .B2(KEYINPUT7), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n204_), .A2(new_n205_), .A3(new_n202_), .A4(new_n203_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n207_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n211_), .A2(KEYINPUT8), .A3(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(new_n203_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n218_));
  INV_X1    g017(.A(G85gat), .ZN(new_n219_));
  INV_X1    g018(.A(G92gat), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT9), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n217_), .A2(new_n218_), .A3(new_n210_), .A4(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n215_), .A2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT8), .B1(new_n211_), .B2(new_n214_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G57gat), .B(G64gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT11), .ZN(new_n227_));
  XOR2_X1   g026(.A(G71gat), .B(G78gat), .Z(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n227_), .A2(new_n228_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n226_), .A2(KEYINPUT11), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n225_), .B(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G230gat), .A2(G233gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n232_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n223_), .A2(new_n232_), .A3(new_n224_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT12), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT66), .B1(new_n223_), .B2(new_n224_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n211_), .A2(new_n214_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT8), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n215_), .A4(new_n222_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n240_), .A2(new_n245_), .A3(KEYINPUT12), .A4(new_n232_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n246_), .A3(new_n234_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n235_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G120gat), .B(G148gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT5), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n250_), .B(KEYINPUT67), .Z(new_n251_));
  XOR2_X1   g050(.A(G176gat), .B(G204gat), .Z(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n235_), .A2(new_n247_), .A3(new_n253_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT13), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(KEYINPUT13), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G15gat), .B(G22gat), .ZN(new_n262_));
  INV_X1    g061(.A(G1gat), .ZN(new_n263_));
  INV_X1    g062(.A(G8gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT14), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G1gat), .B(G8gat), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n267_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G29gat), .B(G36gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(G43gat), .B(G50gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G43gat), .B(G50gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(G29gat), .B(G36gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n270_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(new_n269_), .A3(new_n268_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G229gat), .A2(G233gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT15), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n277_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n270_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n280_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n283_), .B1(new_n287_), .B2(new_n282_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G113gat), .B(G141gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G169gat), .B(G197gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n288_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n261_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G22gat), .B(G50gat), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G211gat), .B(G218gat), .Z(new_n298_));
  INV_X1    g097(.A(G197gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G204gat), .ZN(new_n300_));
  INV_X1    g099(.A(G204gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G197gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT21), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT85), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT85), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n300_), .A2(new_n302_), .A3(new_n306_), .A4(new_n303_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n298_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT83), .B1(new_n301_), .B2(G197gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT83), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(new_n299_), .A3(G204gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n311_), .A3(new_n302_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT21), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n313_), .B1(new_n312_), .B2(KEYINPUT21), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n308_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n300_), .A2(new_n302_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n298_), .A2(KEYINPUT21), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G141gat), .ZN(new_n320_));
  INV_X1    g119(.A(G148gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325_));
  OR2_X1    g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329_));
  INV_X1    g128(.A(new_n325_), .ZN(new_n330_));
  OAI22_X1  g129(.A1(new_n328_), .A2(new_n329_), .B1(KEYINPUT1), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n325_), .A2(KEYINPUT77), .A3(new_n327_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n324_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT79), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n323_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(new_n323_), .B2(new_n336_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n340_), .A2(new_n320_), .A3(new_n321_), .A4(KEYINPUT78), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342_));
  OAI22_X1  g141(.A1(new_n342_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n334_), .B1(new_n339_), .B2(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n341_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n323_), .A2(new_n336_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT79), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n323_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(KEYINPUT80), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n330_), .A2(new_n326_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n333_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n319_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT81), .B(G233gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G228gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT82), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT86), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n361_), .B1(new_n319_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n363_), .ZN(new_n364_));
  OAI221_X1 g163(.A(new_n319_), .B1(new_n362_), .B2(new_n361_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n297_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n365_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n366_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n296_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n356_), .A2(new_n357_), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n375_), .B(KEYINPUT28), .Z(new_n376_));
  AND3_X1   g175(.A1(new_n370_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G127gat), .B(G134gat), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n380_), .A2(KEYINPUT76), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(KEYINPUT76), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G113gat), .B(G120gat), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G183gat), .ZN(new_n388_));
  INV_X1    g187(.A(G190gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT23), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(G183gat), .A3(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT74), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(KEYINPUT74), .A2(G169gat), .A3(G176gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT22), .B(G169gat), .ZN(new_n402_));
  INV_X1    g201(.A(G176gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n395_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n388_), .A2(KEYINPUT25), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT25), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G183gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n389_), .A2(KEYINPUT26), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT26), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G190gat), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n409_), .A2(new_n411_), .A3(new_n412_), .A4(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT75), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n408_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n416_), .B1(new_n408_), .B2(new_n415_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n405_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(KEYINPUT30), .B(new_n405_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G71gat), .B(G99gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G43gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G15gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n428_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n426_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT31), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n424_), .A2(new_n431_), .A3(new_n425_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n387_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n386_), .A3(new_n436_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n379_), .A2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n439_), .A2(new_n441_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT0), .ZN(new_n448_));
  INV_X1    g247(.A(G57gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(G85gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT4), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n339_), .A2(new_n345_), .A3(new_n334_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT80), .B1(new_n347_), .B2(new_n351_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n355_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n457_));
  INV_X1    g256(.A(new_n333_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n354_), .B1(new_n346_), .B2(new_n352_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT91), .B1(new_n460_), .B2(new_n333_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n461_), .A3(new_n387_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n386_), .B(KEYINPUT91), .C1(new_n460_), .C2(new_n333_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n453_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n387_), .B(new_n453_), .C1(new_n460_), .C2(new_n333_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G225gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n452_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n462_), .A2(new_n463_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n466_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n473_), .B(new_n451_), .C1(new_n464_), .C2(new_n468_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT96), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT96), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n471_), .A2(new_n477_), .A3(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n318_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n312_), .A2(KEYINPUT21), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT84), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT21), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n480_), .B1(new_n484_), .B2(new_n308_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n486_));
  INV_X1    g285(.A(G169gat), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n487_), .A2(KEYINPUT22), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(KEYINPUT22), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n486_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n402_), .A2(KEYINPUT88), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n403_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n400_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n407_), .A2(new_n396_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n419_), .A2(new_n415_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n485_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n319_), .A2(new_n422_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT20), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G226gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT20), .B1(new_n319_), .B2(new_n422_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n509_), .B1(new_n485_), .B2(new_n498_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n319_), .A2(KEYINPUT89), .A3(new_n497_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n508_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n512_), .A2(KEYINPUT90), .A3(new_n504_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n515_));
  INV_X1    g314(.A(new_n422_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n516_), .B2(new_n485_), .ZN(new_n517_));
  AOI221_X4 g316(.A(new_n509_), .B1(new_n494_), .B2(new_n496_), .C1(new_n316_), .C2(new_n318_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT89), .B1(new_n319_), .B2(new_n497_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n514_), .B1(new_n520_), .B2(new_n505_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n507_), .B1(new_n513_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G8gat), .B(G36gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT18), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G64gat), .B(G92gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n522_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT90), .B1(new_n512_), .B2(new_n504_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n520_), .A2(new_n514_), .A3(new_n505_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n506_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n526_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT27), .B1(new_n528_), .B2(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT20), .A4(new_n505_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n512_), .B2(new_n505_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT27), .B1(new_n535_), .B2(new_n526_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n536_), .B1(new_n531_), .B2(new_n526_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n479_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n526_), .A2(KEYINPUT32), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n540_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n529_), .A2(new_n530_), .ZN(new_n542_));
  AND4_X1   g341(.A1(KEYINPUT95), .A2(new_n542_), .A3(new_n507_), .A4(new_n539_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT95), .B1(new_n531_), .B2(new_n539_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n541_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT33), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n474_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(new_n474_), .B2(new_n546_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n464_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n468_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n470_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n554_), .A2(KEYINPUT92), .A3(KEYINPUT33), .A4(new_n451_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n474_), .A2(KEYINPUT93), .A3(new_n546_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n549_), .A2(new_n551_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n451_), .B1(new_n472_), .B2(new_n467_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n559_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n552_), .A2(new_n466_), .A3(new_n465_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(new_n532_), .A3(new_n528_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n545_), .B1(new_n557_), .B2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n379_), .A2(new_n444_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n446_), .A2(new_n538_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n295_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n270_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n232_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT72), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT71), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT69), .B(KEYINPUT16), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT70), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n576_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n572_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n572_), .A2(new_n581_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n580_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n582_), .B(new_n583_), .C1(new_n571_), .C2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT73), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT34), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n225_), .A2(new_n279_), .B1(new_n592_), .B2(new_n591_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n240_), .A2(new_n285_), .A3(new_n245_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n594_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT68), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT68), .A4(new_n594_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(G190gat), .B(G218gat), .Z(new_n603_));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT36), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n605_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AOI211_X1 g410(.A(new_n597_), .B(new_n611_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n588_), .B1(new_n608_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n602_), .A2(new_n610_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n614_), .B(KEYINPUT37), .C1(new_n602_), .C2(new_n607_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n587_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n568_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT97), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n479_), .B(KEYINPUT98), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n263_), .A3(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT38), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n295_), .A2(new_n587_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n608_), .A2(new_n612_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n567_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n478_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n477_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n628_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n623_), .A2(new_n632_), .ZN(G1324gat));
  NAND2_X1  g432(.A1(new_n528_), .A2(new_n532_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT27), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n537_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n619_), .A2(new_n264_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n639_));
  OAI21_X1  g438(.A(G8gat), .B1(new_n628_), .B2(new_n636_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n639_), .B1(new_n640_), .B2(KEYINPUT39), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(KEYINPUT39), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n640_), .A2(new_n639_), .A3(KEYINPUT39), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n638_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(G1325gat));
  OAI21_X1  g446(.A(G15gat), .B1(new_n628_), .B2(new_n442_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(KEYINPUT41), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(KEYINPUT41), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n618_), .A2(G15gat), .A3(new_n442_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(G1326gat));
  INV_X1    g451(.A(G22gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n627_), .B2(new_n379_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT42), .Z(new_n655_));
  NAND2_X1  g454(.A1(new_n379_), .A2(new_n653_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n618_), .B2(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT101), .Z(G1327gat));
  INV_X1    g457(.A(new_n587_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n625_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n568_), .A2(new_n661_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n662_), .A2(G29gat), .A3(new_n631_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n294_), .A2(new_n587_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666_));
  INV_X1    g465(.A(new_n616_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n565_), .A2(new_n566_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n377_), .A2(new_n378_), .A3(new_n444_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n376_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n368_), .A2(new_n369_), .A3(new_n297_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n296_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n370_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n442_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n636_), .B(new_n631_), .C1(new_n669_), .C2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n667_), .B1(new_n668_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n666_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n678_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AOI211_X1 g480(.A(KEYINPUT43), .B(new_n667_), .C1(new_n668_), .C2(new_n676_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n666_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n665_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n664_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  NOR4_X1   g486(.A1(new_n567_), .A2(KEYINPUT102), .A3(KEYINPUT43), .A4(new_n667_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n680_), .B2(new_n679_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT104), .B(new_n685_), .C1(new_n689_), .C2(new_n665_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n665_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n567_), .B2(new_n667_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n682_), .B1(new_n693_), .B2(new_n666_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT44), .B(new_n692_), .C1(new_n694_), .C2(new_n688_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n684_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n691_), .A2(new_n699_), .A3(new_n621_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n700_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT106), .B1(new_n700_), .B2(G29gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n663_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(new_n662_), .ZN(new_n704_));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n637_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT45), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n636_), .B1(new_n687_), .B2(new_n690_), .ZN(new_n708_));
  AOI211_X1 g507(.A(KEYINPUT107), .B(new_n705_), .C1(new_n708_), .C2(new_n699_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n691_), .A2(new_n699_), .A3(new_n637_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(G36gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n709_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI211_X1 g514(.A(KEYINPUT46), .B(new_n707_), .C1(new_n709_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND4_X1  g516(.A1(new_n691_), .A2(new_n699_), .A3(G43gat), .A4(new_n444_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT108), .B(G43gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n662_), .B2(new_n442_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n704_), .B2(new_n379_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n691_), .A2(G50gat), .A3(new_n379_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n699_), .ZN(G1331gat));
  NAND4_X1  g525(.A1(new_n626_), .A2(new_n659_), .A3(new_n293_), .A4(new_n261_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT110), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n631_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n567_), .A2(new_n292_), .A3(new_n260_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n617_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n449_), .A3(new_n621_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1332gat));
  INV_X1    g534(.A(G64gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n728_), .B2(new_n637_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT48), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(new_n736_), .A3(new_n637_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1333gat));
  OAI21_X1  g539(.A(G71gat), .B1(new_n729_), .B2(new_n442_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT49), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n442_), .A2(G71gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n732_), .B2(new_n743_), .ZN(G1334gat));
  INV_X1    g543(.A(G78gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n728_), .B2(new_n379_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT50), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n733_), .A2(new_n745_), .A3(new_n379_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n731_), .A2(new_n661_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n219_), .B1(new_n750_), .B2(new_n620_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT111), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n689_), .A2(KEYINPUT112), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n689_), .A2(KEYINPUT112), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n659_), .A2(new_n292_), .A3(new_n260_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n631_), .A2(new_n219_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n752_), .B1(new_n757_), .B2(new_n758_), .ZN(G1336gat));
  INV_X1    g558(.A(new_n750_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G92gat), .B1(new_n760_), .B2(new_n637_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n636_), .A2(new_n220_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT113), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n757_), .B2(new_n763_), .ZN(G1337gat));
  OAI21_X1  g563(.A(G99gat), .B1(new_n756_), .B2(new_n442_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n760_), .A2(new_n216_), .A3(new_n444_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g567(.A1(new_n755_), .A2(new_n379_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G106gat), .B1(new_n689_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT52), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n760_), .A2(new_n203_), .A3(new_n379_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g573(.A1(new_n621_), .A2(new_n636_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(new_n445_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n288_), .A2(new_n291_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n281_), .A2(new_n282_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n291_), .C1(new_n287_), .C2(new_n282_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n256_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(KEYINPUT115), .A3(new_n256_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n247_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n239_), .A2(new_n246_), .A3(KEYINPUT55), .A4(new_n234_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n239_), .A2(new_n246_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n788_), .B(new_n789_), .C1(new_n234_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n254_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(KEYINPUT56), .A3(new_n254_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n786_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT116), .B(new_n616_), .C1(new_n797_), .C2(KEYINPUT58), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT58), .B1(new_n786_), .B2(new_n796_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n667_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n797_), .A2(KEYINPUT58), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n798_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n791_), .B2(new_n254_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n806_), .A2(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n256_), .A2(new_n292_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n806_), .B2(KEYINPUT56), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n257_), .A2(new_n781_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n804_), .B(new_n660_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n807_), .A2(new_n809_), .B1(new_n257_), .B2(new_n781_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT57), .B1(new_n813_), .B2(new_n625_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n803_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n803_), .B2(new_n815_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n587_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n617_), .A2(new_n293_), .A3(new_n260_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n777_), .B1(new_n819_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n659_), .B1(new_n803_), .B2(new_n815_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n822_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n776_), .A2(new_n825_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n827_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n830_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n832_), .B(KEYINPUT118), .C1(new_n822_), .C2(new_n828_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT119), .B1(new_n826_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n833_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n836_), .B(new_n837_), .C1(new_n825_), .C2(new_n824_), .ZN(new_n838_));
  INV_X1    g637(.A(G113gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n293_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n835_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n824_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n839_), .B1(new_n842_), .B2(new_n293_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n841_), .A2(KEYINPUT120), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT120), .B1(new_n841_), .B2(new_n843_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1340gat));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT60), .B1(new_n261_), .B2(new_n847_), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n842_), .A2(KEYINPUT60), .A3(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n842_), .A2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n842_), .A2(KEYINPUT59), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n261_), .A3(new_n836_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n851_), .A2(KEYINPUT121), .A3(new_n261_), .A4(new_n836_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n850_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n849_), .B1(new_n856_), .B2(new_n847_), .ZN(G1341gat));
  NAND3_X1  g656(.A1(new_n835_), .A2(new_n838_), .A3(new_n659_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G127gat), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n587_), .A2(G127gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n842_), .B2(new_n860_), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n667_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n835_), .A2(new_n838_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n824_), .A2(new_n625_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT122), .B1(new_n865_), .B2(new_n862_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  AOI211_X1 g666(.A(new_n867_), .B(G134gat), .C1(new_n824_), .C2(new_n625_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n864_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT123), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n864_), .A2(new_n869_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1343gat));
  AOI21_X1  g673(.A(new_n443_), .B1(new_n819_), .B2(new_n823_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n775_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n293_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n320_), .ZN(G1344gat));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n260_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n321_), .ZN(G1345gat));
  NOR2_X1   g680(.A1(new_n877_), .A2(new_n587_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT61), .B(G155gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  NAND3_X1  g683(.A1(new_n875_), .A2(new_n625_), .A3(new_n876_), .ZN(new_n885_));
  INV_X1    g684(.A(G162gat), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n885_), .A2(KEYINPUT124), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT124), .B1(new_n885_), .B2(new_n886_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n877_), .A2(new_n886_), .A3(new_n667_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(G1347gat));
  NAND3_X1  g689(.A1(new_n620_), .A2(new_n444_), .A3(new_n637_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n829_), .A2(new_n379_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n292_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT125), .Z(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G169gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n896_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n894_), .A2(G169gat), .A3(new_n898_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n892_), .A2(new_n490_), .A3(new_n491_), .A4(new_n292_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n897_), .A2(new_n899_), .A3(new_n900_), .ZN(G1348gat));
  AOI21_X1  g700(.A(G176gat), .B1(new_n892_), .B2(new_n261_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n819_), .A2(new_n823_), .ZN(new_n903_));
  NOR4_X1   g702(.A1(new_n891_), .A2(new_n403_), .A3(new_n379_), .A4(new_n260_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(G1349gat));
  NAND2_X1  g704(.A1(new_n892_), .A2(new_n659_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n388_), .B2(new_n906_), .ZN(G1350gat));
  NAND4_X1  g707(.A1(new_n892_), .A2(new_n625_), .A3(new_n412_), .A4(new_n414_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n892_), .A2(new_n616_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n911_), .B2(new_n389_), .ZN(G1351gat));
  NAND3_X1  g711(.A1(new_n875_), .A2(new_n631_), .A3(new_n637_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n293_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n299_), .ZN(G1352gat));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n260_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n301_), .A2(KEYINPUT127), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n916_), .B(new_n917_), .Z(G1353gat));
  NOR2_X1   g717(.A1(new_n913_), .A2(new_n587_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n922_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  OAI21_X1  g722(.A(G218gat), .B1(new_n913_), .B2(new_n667_), .ZN(new_n924_));
  OR2_X1    g723(.A1(new_n660_), .A2(G218gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n913_), .B2(new_n925_), .ZN(G1355gat));
endmodule


