//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT92), .Z(new_n203_));
  XOR2_X1   g002(.A(G155gat), .B(G162gat), .Z(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n205_));
  INV_X1    g004(.A(G141gat), .ZN(new_n206_));
  INV_X1    g005(.A(G148gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  OAI22_X1  g007(.A1(KEYINPUT84), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT85), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n208_), .B(new_n209_), .C1(new_n211_), .C2(KEYINPUT2), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n211_), .A2(KEYINPUT2), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n204_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n204_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n206_), .A2(new_n207_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n216_), .A2(new_n210_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G113gat), .B(G120gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT4), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n224_), .A2(KEYINPUT90), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n223_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(KEYINPUT90), .A3(new_n223_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n225_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT91), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n226_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AOI211_X1 g032(.A(KEYINPUT91), .B(new_n225_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n203_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n230_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(new_n203_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G1gat), .B(G29gat), .Z(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT93), .B(G85gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G57gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n238_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(G183gat), .A3(G190gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT83), .ZN(new_n248_));
  INV_X1    g047(.A(G183gat), .ZN(new_n249_));
  INV_X1    g048(.A(G190gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT23), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n248_), .B(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(G183gat), .B1(KEYINPUT80), .B2(G190gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(KEYINPUT80), .B2(G190gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G169gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT26), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(new_n250_), .B2(KEYINPUT81), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT81), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n261_), .A2(KEYINPUT80), .A3(KEYINPUT26), .A4(G190gat), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n260_), .B(new_n262_), .C1(KEYINPUT80), .C2(G190gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT25), .B(G183gat), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(KEYINPUT24), .A3(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT82), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n251_), .A2(new_n247_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n266_), .A2(KEYINPUT24), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(KEYINPUT82), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .A4(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n258_), .B1(new_n265_), .B2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G71gat), .B(G99gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G43gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n274_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(new_n223_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G227gat), .A2(G233gat), .ZN(new_n279_));
  INV_X1    g078(.A(G15gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT30), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT31), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n278_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288_));
  OR3_X1    g087(.A1(new_n287_), .A2(KEYINPUT86), .A3(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT86), .B1(new_n287_), .B2(new_n288_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n286_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n287_), .A2(new_n288_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(new_n220_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G228gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G78gat), .B(G106gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(KEYINPUT87), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n298_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n220_), .A2(new_n295_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT28), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G22gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G50gat), .ZN(new_n306_));
  INV_X1    g105(.A(G22gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n304_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G50gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n306_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT88), .B1(new_n298_), .B2(new_n300_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n302_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n306_), .A2(new_n310_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n312_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n314_), .A2(new_n301_), .A3(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n284_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n311_), .A2(new_n302_), .A3(new_n312_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n284_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n301_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n245_), .B1(new_n317_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G8gat), .B(G36gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT18), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G64gat), .B(G92gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT97), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G226gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT19), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n274_), .A2(new_n294_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT26), .B(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n264_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n268_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT89), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(new_n252_), .A3(new_n271_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n270_), .B1(G183gat), .B2(G190gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n257_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT95), .ZN(new_n343_));
  INV_X1    g142(.A(new_n294_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT95), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(new_n345_), .A3(new_n341_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n343_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT20), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n333_), .B1(new_n348_), .B2(KEYINPUT96), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT96), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n350_), .A3(KEYINPUT20), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n331_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n342_), .A2(new_n294_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(KEYINPUT20), .C1(new_n294_), .C2(new_n274_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(new_n330_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n328_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n342_), .A2(new_n294_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n332_), .A2(KEYINPUT20), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n331_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n354_), .B2(new_n331_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n356_), .A2(KEYINPUT98), .B1(new_n360_), .B2(new_n327_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT98), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n362_), .B(new_n328_), .C1(new_n352_), .C2(new_n355_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n323_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n327_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n360_), .B(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n323_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n322_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n313_), .A2(new_n316_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n370_), .A2(new_n284_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n244_), .B1(new_n236_), .B2(new_n203_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n231_), .A2(new_n232_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n234_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n226_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n372_), .B1(new_n375_), .B2(new_n203_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n243_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n366_), .B(new_n376_), .C1(new_n377_), .C2(KEYINPUT33), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(KEYINPUT33), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(KEYINPUT94), .A3(KEYINPUT33), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n378_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n238_), .A2(new_n244_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(new_n377_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n327_), .A2(KEYINPUT32), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n360_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n352_), .A2(new_n355_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n386_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n371_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n369_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT13), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G85gat), .B(G92gat), .ZN(new_n394_));
  INV_X1    g193(.A(G92gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n394_), .B1(KEYINPUT9), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(KEYINPUT9), .B2(new_n394_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT65), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n396_), .B(KEYINPUT65), .C1(KEYINPUT9), .C2(new_n394_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G99gat), .A2(G106gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT6), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(G99gat), .A3(G106gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(KEYINPUT10), .B(G99gat), .Z(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT64), .B(G106gat), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n401_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G57gat), .B(G64gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G71gat), .B(G78gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(KEYINPUT11), .ZN(new_n414_));
  XOR2_X1   g213(.A(G71gat), .B(G78gat), .Z(new_n415_));
  INV_X1    g214(.A(G64gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G57gat), .ZN(new_n417_));
  INV_X1    g216(.A(G57gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G64gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n419_), .A3(KEYINPUT11), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n412_), .A2(KEYINPUT11), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n414_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT68), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT7), .ZN(new_n426_));
  INV_X1    g225(.A(G99gat), .ZN(new_n427_));
  INV_X1    g226(.A(G106gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  AOI211_X1 g230(.A(KEYINPUT8), .B(new_n394_), .C1(new_n431_), .C2(new_n406_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT8), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n404_), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n402_), .A2(KEYINPUT6), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT66), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT66), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n403_), .A2(new_n405_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n439_), .A3(new_n431_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n394_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n434_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT67), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n433_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n438_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n429_), .A2(new_n430_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n394_), .B1(new_n447_), .B2(new_n439_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n448_), .A2(KEYINPUT67), .A3(new_n434_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n411_), .B(new_n425_), .C1(new_n444_), .C2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT69), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n403_), .A2(new_n405_), .A3(new_n438_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n453_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT8), .B1(new_n454_), .B2(new_n394_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT67), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n442_), .A2(new_n443_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n433_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n458_), .A2(KEYINPUT69), .A3(new_n425_), .A4(new_n411_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n411_), .B1(new_n444_), .B2(new_n449_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n425_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n452_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G230gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT12), .ZN(new_n467_));
  INV_X1    g266(.A(new_n410_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n432_), .B1(new_n455_), .B2(KEYINPUT67), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n469_), .B1(new_n470_), .B2(new_n457_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n467_), .B1(new_n471_), .B2(new_n425_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n423_), .A2(new_n467_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n460_), .A2(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n472_), .A2(new_n464_), .A3(new_n475_), .A4(new_n450_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n466_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G120gat), .B(G148gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(G176gat), .B(G204gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n482_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n466_), .A2(new_n476_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n393_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(KEYINPUT13), .A3(new_n486_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT71), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n488_), .A2(KEYINPUT71), .A3(new_n489_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G1gat), .A2(G8gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n280_), .A2(G22gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n307_), .A2(G15gat), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT74), .ZN(new_n502_));
  AND2_X1   g301(.A1(G1gat), .A2(G8gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(G1gat), .A2(G8gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT75), .B1(new_n503_), .B2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(G1gat), .A2(G8gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT75), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n497_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n501_), .A2(new_n505_), .A3(new_n507_), .A4(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n505_), .A2(new_n498_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n507_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G36gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G29gat), .ZN(new_n518_));
  INV_X1    g317(.A(G29gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(G36gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n309_), .A2(G43gat), .ZN(new_n522_));
  INV_X1    g321(.A(G43gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(G50gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n518_), .A2(new_n520_), .A3(new_n522_), .A4(new_n524_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n526_), .A2(new_n527_), .A3(KEYINPUT76), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT76), .B1(new_n526_), .B2(new_n527_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT77), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n516_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n533_));
  INV_X1    g332(.A(new_n527_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n518_), .A2(new_n520_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n526_), .A2(new_n527_), .A3(KEYINPUT76), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n536_), .A2(new_n511_), .A3(new_n537_), .A4(new_n515_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT77), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n532_), .A2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n537_), .A2(new_n536_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT78), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT78), .ZN(new_n544_));
  AOI211_X1 g343(.A(new_n544_), .B(new_n541_), .C1(new_n532_), .C2(new_n539_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n496_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G169gat), .B(G197gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(KEYINPUT79), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n516_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n526_), .A2(new_n527_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT15), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n540_), .A2(new_n495_), .A3(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n546_), .A2(new_n551_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n551_), .B1(new_n546_), .B2(new_n556_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n494_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n471_), .A2(new_n553_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n460_), .A2(new_n554_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT34), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT35), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n562_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n566_), .A2(new_n567_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G190gat), .B(G218gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT72), .ZN(new_n573_));
  XOR2_X1   g372(.A(G134gat), .B(G162gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT36), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n570_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n562_), .A2(new_n578_), .A3(new_n563_), .A4(new_n568_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n571_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n575_), .B(new_n576_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n571_), .B2(new_n579_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n580_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n516_), .B(new_n592_), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(new_n423_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596_));
  XOR2_X1   g395(.A(G127gat), .B(G155gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT16), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n595_), .A2(new_n596_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n594_), .A2(new_n423_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n594_), .A2(new_n461_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n593_), .A2(new_n425_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n600_), .B(KEYINPUT17), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n591_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n392_), .A2(new_n561_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n611_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n614_), .A2(G1gat), .A3(new_n385_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT38), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n584_), .A2(new_n608_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n392_), .A2(new_n561_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n392_), .A2(KEYINPUT100), .A3(new_n561_), .A4(new_n618_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n385_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n624_), .A2(new_n625_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n617_), .B1(new_n626_), .B2(new_n627_), .ZN(G1324gat));
  INV_X1    g427(.A(new_n614_), .ZN(new_n629_));
  INV_X1    g428(.A(G8gat), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n364_), .A2(new_n368_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n364_), .A2(new_n368_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n619_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n636_));
  OAI21_X1  g435(.A(G8gat), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n636_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n639_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n632_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n632_), .A2(KEYINPUT40), .A3(new_n640_), .A4(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1325gat));
  NAND3_X1  g445(.A1(new_n629_), .A2(new_n280_), .A3(new_n284_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n319_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n280_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(KEYINPUT41), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n648_), .A2(new_n651_), .A3(new_n280_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n647_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT103), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n655_), .B(new_n647_), .C1(new_n650_), .C2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1326gat));
  NAND3_X1  g456(.A1(new_n629_), .A2(new_n307_), .A3(new_n370_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n370_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G22gat), .B1(new_n623_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n660_), .A2(new_n662_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n658_), .B1(new_n663_), .B2(new_n664_), .ZN(G1327gat));
  INV_X1    g464(.A(new_n608_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(new_n588_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n392_), .A2(new_n561_), .A3(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n668_), .A2(G29gat), .A3(new_n385_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n494_), .A2(new_n560_), .A3(new_n666_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n392_), .B2(new_n591_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n586_), .A2(new_n590_), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT43), .B(new_n673_), .C1(new_n369_), .C2(new_n391_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n670_), .B(KEYINPUT44), .C1(new_n672_), .C2(new_n674_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n245_), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n669_), .B1(new_n679_), .B2(G29gat), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT105), .ZN(G1328gat));
  INV_X1    g480(.A(new_n668_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n633_), .A2(KEYINPUT106), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n364_), .A2(KEYINPUT106), .A3(new_n368_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n685_), .A3(new_n517_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n687_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n682_), .A2(new_n685_), .A3(new_n517_), .A4(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n677_), .A2(new_n631_), .A3(new_n678_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(G36gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n693_), .B(new_n695_), .ZN(G1329gat));
  NOR2_X1   g495(.A1(new_n319_), .A2(new_n523_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n677_), .A2(new_n678_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT109), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n677_), .A2(new_n700_), .A3(new_n678_), .A4(new_n697_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n523_), .B1(new_n668_), .B2(new_n319_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT47), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n699_), .A2(new_n705_), .A3(new_n701_), .A4(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1330gat));
  AOI21_X1  g506(.A(G50gat), .B1(new_n682_), .B2(new_n370_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n677_), .A2(new_n678_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n659_), .A2(new_n309_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n709_), .B2(new_n710_), .ZN(G1331gat));
  NAND2_X1  g510(.A1(new_n494_), .A2(new_n560_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n369_), .B2(new_n391_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(new_n609_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(new_n418_), .A3(new_n245_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n618_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n385_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1332gat));
  NAND3_X1  g517(.A1(new_n685_), .A2(KEYINPUT110), .A3(new_n416_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n683_), .A2(new_n684_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(G64gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(new_n714_), .A3(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n685_), .A2(new_n618_), .A3(new_n713_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(G64gat), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n724_), .B2(G64gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n723_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(G1333gat));
  OAI21_X1  g530(.A(G71gat), .B1(new_n716_), .B2(new_n319_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT49), .ZN(new_n733_));
  INV_X1    g532(.A(G71gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n714_), .A2(new_n734_), .A3(new_n284_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n714_), .A2(new_n737_), .A3(new_n370_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G78gat), .B1(new_n716_), .B2(new_n659_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(KEYINPUT50), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(KEYINPUT50), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n738_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT112), .Z(G1335gat));
  AND2_X1   g542(.A1(new_n713_), .A2(new_n667_), .ZN(new_n744_));
  INV_X1    g543(.A(G85gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n245_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n672_), .A2(new_n674_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n666_), .A3(new_n712_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(new_n245_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n749_), .B2(new_n745_), .ZN(G1336gat));
  AOI21_X1  g549(.A(G92gat), .B1(new_n744_), .B2(new_n631_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(KEYINPUT113), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n752_), .A2(KEYINPUT113), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n721_), .A2(new_n395_), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n753_), .B(new_n754_), .C1(new_n748_), .C2(new_n755_), .ZN(G1337gat));
  NAND4_X1  g555(.A1(new_n713_), .A2(new_n408_), .A3(new_n284_), .A4(new_n667_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT115), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n712_), .A2(new_n666_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n284_), .B(new_n759_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G99gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G99gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n758_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g564(.A(new_n370_), .B(new_n759_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G106gat), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT52), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(new_n769_), .A3(G106gat), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n744_), .A2(new_n409_), .A3(new_n370_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1339gat));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778_));
  INV_X1    g577(.A(new_n560_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n490_), .A2(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n609_), .A2(new_n778_), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n778_), .B1(new_n609_), .B2(new_n780_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n549_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n543_), .A2(new_n545_), .A3(new_n496_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n495_), .B1(new_n540_), .B2(new_n555_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n546_), .A2(new_n549_), .A3(new_n556_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n486_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n450_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT12), .B1(new_n460_), .B2(new_n461_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n465_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n465_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(KEYINPUT55), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  NOR4_X1   g596(.A1(new_n792_), .A2(new_n793_), .A3(new_n797_), .A4(new_n465_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n482_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT117), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n791_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n795_), .A2(KEYINPUT55), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n476_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n798_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n485_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n801_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n790_), .B1(new_n802_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT57), .B1(new_n809_), .B2(new_n584_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n790_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n477_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n546_), .A2(new_n556_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n550_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n812_), .A2(new_n485_), .B1(new_n814_), .B2(new_n557_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n799_), .A2(new_n801_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n811_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n588_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n486_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n486_), .A2(new_n787_), .A3(KEYINPUT118), .A4(new_n788_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n799_), .A2(KEYINPUT56), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n806_), .A2(new_n800_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n673_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n825_), .A2(new_n827_), .A3(new_n826_), .A4(KEYINPUT58), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n810_), .A2(new_n820_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n608_), .B1(new_n832_), .B2(KEYINPUT119), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n828_), .A2(new_n829_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n591_), .A3(new_n831_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n809_), .A2(KEYINPUT57), .A3(new_n584_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n819_), .B1(new_n818_), .B2(new_n588_), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT119), .B(new_n835_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n783_), .B1(new_n833_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n608_), .A3(new_n838_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(KEYINPUT120), .A3(new_n783_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n631_), .A2(new_n385_), .A3(new_n317_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n842_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(G113gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n850_), .A3(new_n779_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n783_), .B1(new_n666_), .B2(new_n832_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n852_), .A2(new_n853_), .A3(new_n848_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n842_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n560_), .B(new_n854_), .C1(new_n855_), .C2(KEYINPUT59), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n851_), .B1(new_n856_), .B2(new_n850_), .ZN(G1340gat));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858_));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(KEYINPUT60), .ZN(new_n860_));
  INV_X1    g659(.A(new_n494_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n861_), .A2(KEYINPUT60), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n862_), .B2(new_n859_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n858_), .B1(new_n849_), .B2(new_n863_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n849_), .A2(new_n858_), .A3(new_n863_), .ZN(new_n865_));
  AOI211_X1 g664(.A(new_n861_), .B(new_n854_), .C1(new_n855_), .C2(KEYINPUT59), .ZN(new_n866_));
  OAI22_X1  g665(.A1(new_n864_), .A2(new_n865_), .B1(new_n866_), .B2(new_n859_), .ZN(G1341gat));
  NAND2_X1  g666(.A1(new_n666_), .A2(G127gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT122), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI211_X1 g669(.A(new_n854_), .B(new_n870_), .C1(new_n855_), .C2(KEYINPUT59), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n842_), .A2(new_n666_), .A3(new_n847_), .A4(new_n848_), .ZN(new_n872_));
  INV_X1    g671(.A(G127gat), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT123), .B1(new_n871_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n854_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n877_), .B(new_n869_), .C1(new_n849_), .C2(new_n853_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n879_), .A3(new_n874_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n880_), .ZN(G1342gat));
  INV_X1    g680(.A(G134gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n849_), .A2(new_n882_), .A3(new_n584_), .ZN(new_n883_));
  AOI211_X1 g682(.A(new_n673_), .B(new_n854_), .C1(new_n855_), .C2(KEYINPUT59), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n882_), .ZN(G1343gat));
  NOR2_X1   g684(.A1(new_n840_), .A2(new_n841_), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT120), .B1(new_n846_), .B2(new_n783_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n321_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n888_), .A2(new_n245_), .A3(new_n889_), .A4(new_n721_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G141gat), .B1(new_n890_), .B2(new_n560_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n842_), .A2(new_n847_), .ZN(new_n892_));
  NOR4_X1   g691(.A1(new_n892_), .A2(new_n385_), .A3(new_n321_), .A4(new_n685_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(new_n206_), .A3(new_n779_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n891_), .A2(new_n894_), .ZN(G1344gat));
  OAI21_X1  g694(.A(G148gat), .B1(new_n890_), .B2(new_n861_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n207_), .A3(new_n494_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1345gat));
  XNOR2_X1  g697(.A(KEYINPUT61), .B(G155gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n890_), .B2(new_n608_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n899_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n893_), .A2(new_n666_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1346gat));
  NAND2_X1  g702(.A1(new_n893_), .A2(new_n584_), .ZN(new_n904_));
  INV_X1    g703(.A(G162gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n673_), .A2(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT124), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n904_), .A2(new_n905_), .B1(new_n893_), .B2(new_n907_), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n721_), .A2(new_n245_), .A3(new_n317_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n852_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n560_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT22), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n909_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G169gat), .ZN(new_n915_));
  INV_X1    g714(.A(G169gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n912_), .B2(new_n909_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n914_), .B2(new_n917_), .ZN(G1348gat));
  INV_X1    g717(.A(new_n911_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G176gat), .B1(new_n919_), .B2(new_n494_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n892_), .A2(new_n370_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n721_), .A2(new_n245_), .ZN(new_n922_));
  AND4_X1   g721(.A1(G176gat), .A2(new_n922_), .A3(new_n494_), .A4(new_n284_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n920_), .B1(new_n921_), .B2(new_n923_), .ZN(G1349gat));
  NOR3_X1   g723(.A1(new_n911_), .A2(new_n264_), .A3(new_n608_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n921_), .A2(new_n284_), .A3(new_n666_), .A4(new_n922_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n249_), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n911_), .B2(new_n673_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n584_), .A2(new_n334_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n911_), .B2(new_n929_), .ZN(G1351gat));
  NAND4_X1  g729(.A1(new_n842_), .A2(new_n889_), .A3(new_n847_), .A4(new_n922_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n560_), .ZN(new_n932_));
  XOR2_X1   g731(.A(new_n932_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g732(.A1(new_n931_), .A2(new_n861_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1353gat));
  NOR2_X1   g735(.A1(new_n931_), .A2(new_n608_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n937_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938_));
  XNOR2_X1  g737(.A(KEYINPUT63), .B(G211gat), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n931_), .A2(new_n608_), .A3(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1354gat));
  INV_X1    g740(.A(G218gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n942_), .B1(new_n931_), .B2(new_n588_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n673_), .A2(new_n942_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(KEYINPUT126), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n888_), .A2(new_n889_), .A3(new_n922_), .A4(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n943_), .A2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n943_), .A2(new_n946_), .A3(KEYINPUT127), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1355gat));
endmodule


