// Benchmark "c5315" written by ABC on Wed Jul  6 02:18:28 2022

module c5315 ( 
    G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
    G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
    G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
    G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140,
    G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173,
    G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209,
    G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251,
    G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293,
    G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338,
    G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389,
    G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523,
    G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691,
    G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717,
    G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34,
    G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76,
    G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103,
    G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
    G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137,
    G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170,
    G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206,
    G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248,
    G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292,
    G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335,
    G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386,
    G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514,
    G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690,
    G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552,
    G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire new_n320_, new_n322_, new_n332_, new_n340_, new_n342_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n351_, new_n352_, new_n354_,
    new_n355_, new_n357_, new_n358_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1026_, new_n1027_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_;
  BUF_X1    g0000(.A(G141), .Z(G144));
  BUF_X1    g0001(.A(G293), .Z(G298));
  BUF_X1    g0002(.A(G3173), .Z(G973));
  INV_X1    g0003(.A(G545), .ZN(G594));
  INV_X1    g0004(.A(G348), .ZN(G599));
  INV_X1    g0005(.A(G366), .ZN(G600));
  INV_X1    g0006(.A(G552), .ZN(G849));
  INV_X1    g0007(.A(G562), .ZN(G850));
  NOR2_X1   g0008(.A1(G849), .A2(G850), .ZN(G601));
  INV_X1    g0009(.A(G549), .ZN(G602));
  INV_X1    g0010(.A(G545), .ZN(G603));
  INV_X1    g0011(.A(G545), .ZN(G604));
  INV_X1    g0012(.A(G338), .ZN(G611));
  INV_X1    g0013(.A(G358), .ZN(G612));
  AND2_X1   g0014(.A1(G141), .A2(G145), .ZN(G810));
  INV_X1    g0015(.A(G245), .ZN(G848));
  INV_X1    g0016(.A(G559), .ZN(G851));
  AND2_X1   g0017(.A1(G1), .A2(G373), .ZN(G634));
  INV_X1    g0018(.A(G136), .ZN(new_n320_));
  NOR2_X1   g0019(.A1(new_n320_), .A2(G3173), .ZN(G815));
  INV_X1    g0020(.A(G2824), .ZN(new_n322_));
  NAND2_X1  g0021(.A1(new_n322_), .A2(G27), .ZN(G845));
  NAND2_X1  g0022(.A1(G386), .A2(G556), .ZN(G847));
  BUF_X1    g0023(.A(G137), .Z(G926));
  BUF_X1    g0024(.A(G141), .Z(G923));
  BUF_X1    g0025(.A(G1), .Z(G921));
  BUF_X1    g0026(.A(G549), .Z(G892));
  BUF_X1    g0027(.A(G299), .Z(G887));
  INV_X1    g0028(.A(G549), .ZN(G606));
  NAND2_X1  g0029(.A1(G27), .A2(G31), .ZN(G809));
  INV_X1    g0030(.A(G809), .ZN(new_n332_));
  NAND2_X1  g0031(.A1(new_n332_), .A2(G140), .ZN(G656));
  BUF_X1    g0032(.A(G1), .Z(G993));
  BUF_X1    g0033(.A(G1), .Z(G978));
  BUF_X1    g0034(.A(G1), .Z(G949));
  BUF_X1    g0035(.A(G1), .Z(G939));
  BUF_X1    g0036(.A(G299), .Z(G889));
  INV_X1    g0037(.A(G299), .ZN(G593));
  MUX2_X1   g0038(.A(G86), .B(G87), .S(G2358), .Z(new_n340_));
  NAND2_X1  g0039(.A1(new_n340_), .A2(new_n332_), .ZN(G636));
  MUX2_X1   g0040(.A(G88), .B(G34), .S(G2358), .Z(new_n342_));
  NAND2_X1  g0041(.A1(new_n342_), .A2(new_n332_), .ZN(G704));
  NAND2_X1  g0042(.A1(new_n342_), .A2(new_n332_), .ZN(G717));
  NAND3_X1  g0043(.A1(G27), .A2(G31), .A3(G83), .ZN(G820));
  INV_X1    g0044(.A(G141), .ZN(new_n346_));
  NAND3_X1  g0045(.A1(new_n332_), .A2(G25), .A3(G2358), .ZN(new_n347_));
  INV_X1    g0046(.A(G2358), .ZN(new_n348_));
  AOI21_X1  g0047(.A(G809), .B1(G24), .B2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g0048(.A(new_n346_), .B1(new_n347_), .B2(new_n349_), .ZN(G639));
  NAND3_X1  g0049(.A1(new_n332_), .A2(G81), .A3(G2358), .ZN(new_n351_));
  AOI21_X1  g0050(.A(G809), .B1(G26), .B2(new_n348_), .ZN(new_n352_));
  AOI21_X1  g0051(.A(new_n346_), .B1(new_n351_), .B2(new_n352_), .ZN(G673));
  NAND3_X1  g0052(.A1(new_n332_), .A2(G23), .A3(G2358), .ZN(new_n354_));
  AOI21_X1  g0053(.A(G809), .B1(G79), .B2(new_n348_), .ZN(new_n355_));
  AOI21_X1  g0054(.A(new_n346_), .B1(new_n354_), .B2(new_n355_), .ZN(G707));
  NAND3_X1  g0055(.A1(new_n332_), .A2(G80), .A3(G2358), .ZN(new_n357_));
  AOI21_X1  g0056(.A(G809), .B1(G82), .B2(new_n348_), .ZN(new_n358_));
  AOI21_X1  g0057(.A(new_n346_), .B1(new_n357_), .B2(new_n358_), .ZN(G715));
  INV_X1    g0058(.A(G251), .ZN(new_n360_));
  NOR2_X1   g0059(.A1(new_n360_), .A2(G302), .ZN(new_n361_));
  AOI21_X1  g0060(.A(new_n361_), .B1(G248), .B2(G302), .ZN(new_n362_));
  NAND2_X1  g0061(.A1(G242), .A2(G293), .ZN(new_n363_));
  INV_X1    g0062(.A(G254), .ZN(new_n364_));
  OAI21_X1  g0063(.A(new_n363_), .B1(new_n364_), .B2(G293), .ZN(new_n365_));
  NOR2_X1   g0064(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g0065(.A(G479), .B1(G242), .B2(G308), .ZN(new_n367_));
  OAI21_X1  g0066(.A(new_n367_), .B1(new_n364_), .B2(G308), .ZN(new_n368_));
  NAND3_X1  g0067(.A1(G248), .A2(G308), .A3(G479), .ZN(new_n369_));
  INV_X1    g0068(.A(G308), .ZN(new_n370_));
  NAND3_X1  g0069(.A1(new_n370_), .A2(G251), .A3(G479), .ZN(new_n371_));
  NAND3_X1  g0070(.A1(new_n368_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g0071(.A(G490), .B1(G242), .B2(G316), .ZN(new_n373_));
  OAI21_X1  g0072(.A(new_n373_), .B1(new_n364_), .B2(G316), .ZN(new_n374_));
  NAND3_X1  g0073(.A1(G248), .A2(G316), .A3(G490), .ZN(new_n375_));
  INV_X1    g0074(.A(G316), .ZN(new_n376_));
  NAND3_X1  g0075(.A1(new_n376_), .A2(G251), .A3(G490), .ZN(new_n377_));
  NAND3_X1  g0076(.A1(new_n374_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  NAND3_X1  g0077(.A1(new_n366_), .A2(new_n372_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g0078(.A(G3552), .ZN(new_n380_));
  NAND3_X1  g0079(.A1(new_n380_), .A2(G341), .A3(G523), .ZN(new_n381_));
  INV_X1    g0080(.A(G341), .ZN(new_n382_));
  INV_X1    g0081(.A(G3550), .ZN(new_n383_));
  NAND3_X1  g0082(.A1(new_n382_), .A2(new_n383_), .A3(G523), .ZN(new_n384_));
  INV_X1    g0083(.A(G523), .ZN(new_n385_));
  OAI21_X1  g0084(.A(new_n385_), .B1(new_n382_), .B2(G3546), .ZN(new_n386_));
  NOR2_X1   g0085(.A1(G341), .A2(G3548), .ZN(new_n387_));
  OAI211_X1 g0086(.A(new_n381_), .B(new_n384_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g0087(.A1(new_n380_), .A2(G351), .A3(G534), .ZN(new_n389_));
  INV_X1    g0088(.A(G351), .ZN(new_n390_));
  NAND3_X1  g0089(.A1(new_n390_), .A2(new_n383_), .A3(G534), .ZN(new_n391_));
  INV_X1    g0090(.A(G534), .ZN(new_n392_));
  OAI21_X1  g0091(.A(new_n392_), .B1(new_n390_), .B2(G3546), .ZN(new_n393_));
  NOR2_X1   g0092(.A1(G351), .A2(G3548), .ZN(new_n394_));
  OAI211_X1 g0093(.A(new_n389_), .B(new_n391_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g0094(.A1(new_n380_), .A2(G324), .A3(G503), .ZN(new_n396_));
  INV_X1    g0095(.A(G324), .ZN(new_n397_));
  NAND3_X1  g0096(.A1(new_n397_), .A2(new_n383_), .A3(G503), .ZN(new_n398_));
  INV_X1    g0097(.A(G503), .ZN(new_n399_));
  OAI21_X1  g0098(.A(new_n399_), .B1(new_n397_), .B2(G3546), .ZN(new_n400_));
  NOR2_X1   g0099(.A1(G324), .A2(G3548), .ZN(new_n401_));
  OAI211_X1 g0100(.A(new_n396_), .B(new_n398_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n402_));
  INV_X1    g0101(.A(G514), .ZN(new_n403_));
  NAND2_X1  g0102(.A1(new_n403_), .A2(G3546), .ZN(new_n404_));
  OAI21_X1  g0103(.A(new_n404_), .B1(new_n403_), .B2(G3552), .ZN(new_n405_));
  NAND4_X1  g0104(.A1(new_n388_), .A2(new_n395_), .A3(new_n402_), .A4(new_n405_), .ZN(new_n406_));
  NAND2_X1  g0105(.A1(G248), .A2(G361), .ZN(new_n407_));
  OAI21_X1  g0106(.A(new_n407_), .B1(new_n360_), .B2(G361), .ZN(new_n408_));
  INV_X1    g0107(.A(new_n408_), .ZN(new_n409_));
  NOR3_X1   g0108(.A1(new_n379_), .A2(new_n406_), .A3(new_n409_), .ZN(G598));
  NAND3_X1  g0109(.A1(new_n380_), .A2(G218), .A3(G468), .ZN(new_n411_));
  INV_X1    g0110(.A(G218), .ZN(new_n412_));
  NAND2_X1  g0111(.A1(new_n412_), .A2(G468), .ZN(new_n413_));
  INV_X1    g0112(.A(G468), .ZN(new_n414_));
  OAI21_X1  g0113(.A(new_n414_), .B1(new_n412_), .B2(G3546), .ZN(new_n415_));
  NOR2_X1   g0114(.A1(G218), .A2(G3548), .ZN(new_n416_));
  OAI221_X1 g0115(.A(new_n411_), .B1(new_n413_), .B2(G3550), .C1(new_n415_), .C2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g0116(.A1(new_n380_), .A2(G226), .A3(G422), .ZN(new_n418_));
  INV_X1    g0117(.A(G226), .ZN(new_n419_));
  NAND3_X1  g0118(.A1(new_n419_), .A2(new_n383_), .A3(G422), .ZN(new_n420_));
  INV_X1    g0119(.A(G422), .ZN(new_n421_));
  OAI21_X1  g0120(.A(new_n421_), .B1(new_n419_), .B2(G3546), .ZN(new_n422_));
  NOR2_X1   g0121(.A1(G226), .A2(G3548), .ZN(new_n423_));
  OAI211_X1 g0122(.A(new_n418_), .B(new_n420_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g0123(.A1(new_n380_), .A2(G234), .A3(G435), .ZN(new_n425_));
  INV_X1    g0124(.A(G234), .ZN(new_n426_));
  NAND3_X1  g0125(.A1(new_n426_), .A2(new_n383_), .A3(G435), .ZN(new_n427_));
  INV_X1    g0126(.A(G435), .ZN(new_n428_));
  OAI21_X1  g0127(.A(new_n428_), .B1(new_n426_), .B2(G3546), .ZN(new_n429_));
  NOR2_X1   g0128(.A1(G234), .A2(G3548), .ZN(new_n430_));
  OAI211_X1 g0129(.A(new_n425_), .B(new_n427_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g0130(.A1(new_n380_), .A2(G210), .A3(G457), .ZN(new_n432_));
  INV_X1    g0131(.A(G210), .ZN(new_n433_));
  NAND3_X1  g0132(.A1(new_n433_), .A2(new_n383_), .A3(G457), .ZN(new_n434_));
  INV_X1    g0133(.A(G457), .ZN(new_n435_));
  OAI21_X1  g0134(.A(new_n435_), .B1(new_n433_), .B2(G3546), .ZN(new_n436_));
  NOR2_X1   g0135(.A1(G210), .A2(G3548), .ZN(new_n437_));
  OAI211_X1 g0136(.A(new_n432_), .B(new_n434_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g0137(.A1(new_n417_), .A2(new_n424_), .A3(new_n431_), .A4(new_n438_), .ZN(new_n439_));
  NAND3_X1  g0138(.A1(new_n380_), .A2(G281), .A3(G374), .ZN(new_n440_));
  INV_X1    g0139(.A(G281), .ZN(new_n441_));
  NAND3_X1  g0140(.A1(new_n441_), .A2(new_n383_), .A3(G374), .ZN(new_n442_));
  INV_X1    g0141(.A(G374), .ZN(new_n443_));
  OAI21_X1  g0142(.A(new_n443_), .B1(new_n441_), .B2(G3546), .ZN(new_n444_));
  NOR2_X1   g0143(.A1(G281), .A2(G3548), .ZN(new_n445_));
  OAI211_X1 g0144(.A(new_n440_), .B(new_n442_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g0145(.A1(new_n380_), .A2(G273), .A3(G411), .ZN(new_n447_));
  INV_X1    g0146(.A(G273), .ZN(new_n448_));
  NAND3_X1  g0147(.A1(new_n448_), .A2(new_n383_), .A3(G411), .ZN(new_n449_));
  INV_X1    g0148(.A(G411), .ZN(new_n450_));
  OAI21_X1  g0149(.A(new_n450_), .B1(new_n448_), .B2(G3546), .ZN(new_n451_));
  NOR2_X1   g0150(.A1(G273), .A2(G3548), .ZN(new_n452_));
  OAI211_X1 g0151(.A(new_n447_), .B(new_n449_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g0152(.A1(new_n380_), .A2(G257), .A3(G389), .ZN(new_n454_));
  INV_X1    g0153(.A(G257), .ZN(new_n455_));
  NAND3_X1  g0154(.A1(new_n455_), .A2(new_n383_), .A3(G389), .ZN(new_n456_));
  INV_X1    g0155(.A(G389), .ZN(new_n457_));
  OAI21_X1  g0156(.A(new_n457_), .B1(new_n455_), .B2(G3546), .ZN(new_n458_));
  NOR2_X1   g0157(.A1(G257), .A2(G3548), .ZN(new_n459_));
  OAI211_X1 g0158(.A(new_n454_), .B(new_n456_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g0159(.A1(new_n380_), .A2(G265), .A3(G400), .ZN(new_n461_));
  INV_X1    g0160(.A(G265), .ZN(new_n462_));
  NAND3_X1  g0161(.A1(new_n462_), .A2(new_n383_), .A3(G400), .ZN(new_n463_));
  INV_X1    g0162(.A(G400), .ZN(new_n464_));
  OAI21_X1  g0163(.A(new_n464_), .B1(new_n462_), .B2(G3546), .ZN(new_n465_));
  NOR2_X1   g0164(.A1(G265), .A2(G3548), .ZN(new_n466_));
  OAI211_X1 g0165(.A(new_n461_), .B(new_n463_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g0166(.A1(new_n446_), .A2(new_n453_), .A3(new_n460_), .A4(new_n467_), .ZN(new_n468_));
  AOI21_X1  g0167(.A(G446), .B1(G206), .B2(G242), .ZN(new_n469_));
  OAI21_X1  g0168(.A(new_n469_), .B1(G206), .B2(new_n364_), .ZN(new_n470_));
  NAND3_X1  g0169(.A1(G206), .A2(G248), .A3(G446), .ZN(new_n471_));
  INV_X1    g0170(.A(G206), .ZN(new_n472_));
  NAND3_X1  g0171(.A1(new_n472_), .A2(G251), .A3(G446), .ZN(new_n473_));
  NAND3_X1  g0172(.A1(new_n470_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g0173(.A(new_n474_), .ZN(new_n475_));
  NOR3_X1   g0174(.A1(new_n439_), .A2(new_n468_), .A3(new_n475_), .ZN(G610));
  NAND2_X1  g0175(.A1(G264), .A2(G335), .ZN(new_n477_));
  OAI21_X1  g0176(.A(new_n477_), .B1(new_n455_), .B2(G335), .ZN(new_n478_));
  XNOR2_X1  g0177(.A(new_n478_), .B(new_n457_), .ZN(new_n479_));
  INV_X1    g0178(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g0179(.A1(G272), .A2(G335), .ZN(new_n481_));
  OAI211_X1 g0180(.A(new_n481_), .B(G400), .C1(new_n462_), .C2(G335), .ZN(new_n482_));
  INV_X1    g0181(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g0182(.A(G335), .ZN(new_n484_));
  NAND2_X1  g0183(.A1(new_n484_), .A2(G265), .ZN(new_n485_));
  AOI21_X1  g0184(.A(G400), .B1(new_n485_), .B2(new_n481_), .ZN(new_n486_));
  NOR2_X1   g0185(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g0186(.A1(G241), .A2(G335), .ZN(new_n488_));
  OAI21_X1  g0187(.A(new_n488_), .B1(new_n426_), .B2(G335), .ZN(new_n489_));
  XNOR2_X1  g0188(.A(new_n489_), .B(G435), .ZN(new_n490_));
  NOR3_X1   g0189(.A1(new_n480_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g0190(.A1(G280), .A2(G335), .ZN(new_n492_));
  OAI21_X1  g0191(.A(new_n492_), .B1(new_n448_), .B2(G335), .ZN(new_n493_));
  NAND2_X1  g0192(.A1(new_n493_), .A2(new_n450_), .ZN(new_n494_));
  OAI211_X1 g0193(.A(new_n492_), .B(G411), .C1(new_n448_), .C2(G335), .ZN(new_n495_));
  NAND2_X1  g0194(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g0195(.A1(new_n484_), .A2(G281), .ZN(new_n497_));
  NAND2_X1  g0196(.A1(G288), .A2(G335), .ZN(new_n498_));
  NAND2_X1  g0197(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g0198(.A(new_n499_), .B(new_n443_), .ZN(new_n500_));
  NAND3_X1  g0199(.A1(new_n491_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g0200(.A1(new_n484_), .A2(G226), .ZN(new_n502_));
  NAND2_X1  g0201(.A1(G233), .A2(G335), .ZN(new_n503_));
  NAND2_X1  g0202(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g0203(.A(new_n504_), .B(G422), .ZN(new_n505_));
  INV_X1    g0204(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g0205(.A1(G209), .A2(G335), .ZN(new_n507_));
  OAI21_X1  g0206(.A(new_n507_), .B1(new_n472_), .B2(G335), .ZN(new_n508_));
  XNOR2_X1  g0207(.A(new_n508_), .B(G446), .ZN(new_n509_));
  INV_X1    g0208(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g0209(.A1(new_n484_), .A2(G218), .ZN(new_n511_));
  NAND2_X1  g0210(.A1(G225), .A2(G335), .ZN(new_n512_));
  AND2_X1   g0211(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g0212(.A1(new_n513_), .A2(G468), .ZN(new_n514_));
  NAND2_X1  g0213(.A1(new_n511_), .A2(new_n512_), .ZN(new_n515_));
  NAND2_X1  g0214(.A1(new_n515_), .A2(new_n414_), .ZN(new_n516_));
  NAND2_X1  g0215(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g0216(.A1(G217), .A2(G335), .ZN(new_n518_));
  OAI21_X1  g0217(.A(new_n518_), .B1(new_n433_), .B2(G335), .ZN(new_n519_));
  XNOR2_X1  g0218(.A(new_n519_), .B(new_n435_), .ZN(new_n520_));
  NAND4_X1  g0219(.A1(new_n506_), .A2(new_n510_), .A3(new_n517_), .A4(new_n520_), .ZN(new_n521_));
  NOR2_X1   g0220(.A1(new_n501_), .A2(new_n521_), .ZN(G588));
  INV_X1    g0221(.A(G332), .ZN(new_n523_));
  NAND2_X1  g0222(.A1(new_n523_), .A2(G316), .ZN(new_n524_));
  NAND2_X1  g0223(.A1(G323), .A2(G332), .ZN(new_n525_));
  NAND2_X1  g0224(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g0225(.A(new_n526_), .B(G490), .ZN(new_n527_));
  INV_X1    g0226(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g0227(.A1(G307), .A2(G332), .ZN(new_n529_));
  INV_X1    g0228(.A(G302), .ZN(new_n530_));
  OAI21_X1  g0229(.A(new_n529_), .B1(new_n530_), .B2(G332), .ZN(new_n531_));
  INV_X1    g0230(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g0231(.A1(G299), .A2(G332), .ZN(new_n533_));
  INV_X1    g0232(.A(G293), .ZN(new_n534_));
  OAI21_X1  g0233(.A(new_n533_), .B1(new_n534_), .B2(G332), .ZN(new_n535_));
  INV_X1    g0234(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g0235(.A1(new_n523_), .A2(G308), .ZN(new_n537_));
  NAND2_X1  g0236(.A1(G315), .A2(G332), .ZN(new_n538_));
  NAND2_X1  g0237(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g0238(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g0239(.A1(new_n540_), .A2(G479), .ZN(new_n541_));
  INV_X1    g0240(.A(G479), .ZN(new_n542_));
  NAND2_X1  g0241(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g0242(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g0243(.A1(new_n528_), .A2(new_n532_), .A3(new_n536_), .A4(new_n544_), .ZN(new_n545_));
  NAND2_X1  g0244(.A1(G331), .A2(G332), .ZN(new_n546_));
  OAI21_X1  g0245(.A(new_n546_), .B1(new_n397_), .B2(G332), .ZN(new_n547_));
  XNOR2_X1  g0246(.A(new_n547_), .B(G503), .ZN(new_n548_));
  INV_X1    g0247(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g0248(.A1(G611), .A2(G332), .ZN(new_n550_));
  NAND2_X1  g0249(.A1(new_n550_), .A2(new_n403_), .ZN(new_n551_));
  NAND3_X1  g0250(.A1(G611), .A2(G332), .A3(G514), .ZN(new_n552_));
  NAND2_X1  g0251(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g0252(.A1(new_n523_), .A2(G341), .ZN(new_n554_));
  NAND2_X1  g0253(.A1(G332), .A2(G348), .ZN(new_n555_));
  NAND2_X1  g0254(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g0255(.A1(new_n556_), .A2(new_n385_), .ZN(new_n557_));
  NAND3_X1  g0256(.A1(new_n554_), .A2(G523), .A3(new_n555_), .ZN(new_n558_));
  NAND2_X1  g0257(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g0258(.A1(G332), .A2(G358), .ZN(new_n560_));
  OAI21_X1  g0259(.A(new_n560_), .B1(new_n390_), .B2(G332), .ZN(new_n561_));
  NAND2_X1  g0260(.A1(new_n561_), .A2(new_n392_), .ZN(new_n562_));
  NAND2_X1  g0261(.A1(new_n523_), .A2(G351), .ZN(new_n563_));
  NAND3_X1  g0262(.A1(new_n563_), .A2(G534), .A3(new_n560_), .ZN(new_n564_));
  NAND2_X1  g0263(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g0264(.A1(new_n549_), .A2(new_n553_), .A3(new_n559_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g0265(.A1(G332), .A2(G366), .ZN(new_n567_));
  INV_X1    g0266(.A(G361), .ZN(new_n568_));
  OAI21_X1  g0267(.A(new_n567_), .B1(new_n568_), .B2(G332), .ZN(new_n569_));
  NOR3_X1   g0268(.A1(new_n545_), .A2(new_n566_), .A3(new_n569_), .ZN(G615));
  INV_X1    g0269(.A(new_n558_), .ZN(new_n571_));
  AOI21_X1  g0270(.A(G523), .B1(new_n554_), .B2(new_n555_), .ZN(new_n572_));
  NOR2_X1   g0271(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g0272(.A(new_n553_), .ZN(new_n574_));
  NOR3_X1   g0273(.A1(new_n548_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g0274(.A(new_n569_), .ZN(new_n576_));
  NAND3_X1  g0275(.A1(new_n575_), .A2(new_n576_), .A3(new_n565_), .ZN(new_n577_));
  NAND4_X1  g0276(.A1(new_n528_), .A2(new_n532_), .A3(new_n536_), .A4(new_n544_), .ZN(new_n578_));
  NOR2_X1   g0277(.A1(new_n577_), .A2(new_n578_), .ZN(G626));
  NAND4_X1  g0278(.A1(new_n506_), .A2(new_n510_), .A3(new_n517_), .A4(new_n520_), .ZN(new_n580_));
  INV_X1    g0279(.A(new_n490_), .ZN(new_n581_));
  OAI21_X1  g0280(.A(new_n481_), .B1(new_n462_), .B2(G335), .ZN(new_n582_));
  NAND2_X1  g0281(.A1(new_n582_), .A2(new_n464_), .ZN(new_n583_));
  NAND2_X1  g0282(.A1(new_n583_), .A2(new_n482_), .ZN(new_n584_));
  NAND4_X1  g0283(.A1(new_n581_), .A2(new_n479_), .A3(new_n496_), .A4(new_n584_), .ZN(new_n585_));
  INV_X1    g0284(.A(new_n500_), .ZN(new_n586_));
  NOR3_X1   g0285(.A1(new_n580_), .A2(new_n585_), .A3(new_n586_), .ZN(G632));
  XNOR2_X1  g0286(.A(G341), .B(G351), .ZN(new_n588_));
  INV_X1    g0287(.A(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g0288(.A(G361), .B(G369), .ZN(new_n590_));
  INV_X1    g0289(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g0290(.A1(new_n589_), .A2(new_n591_), .A3(new_n397_), .ZN(new_n592_));
  NAND3_X1  g0291(.A1(new_n591_), .A2(G324), .A3(new_n588_), .ZN(new_n593_));
  NAND3_X1  g0292(.A1(new_n589_), .A2(G324), .A3(new_n590_), .ZN(new_n594_));
  NAND3_X1  g0293(.A1(new_n588_), .A2(new_n590_), .A3(new_n397_), .ZN(new_n595_));
  NAND4_X1  g0294(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g0295(.A(G308), .B(G316), .ZN(new_n597_));
  XNOR2_X1  g0296(.A(G293), .B(G302), .ZN(new_n598_));
  XNOR2_X1  g0297(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g0298(.A(new_n596_), .B(new_n599_), .ZN(G1002));
  XNOR2_X1  g0299(.A(G265), .B(G273), .ZN(new_n601_));
  INV_X1    g0300(.A(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g0301(.A(G234), .B(G257), .ZN(new_n603_));
  INV_X1    g0302(.A(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g0303(.A(G281), .B(G289), .ZN(new_n605_));
  INV_X1    g0304(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g0305(.A1(new_n602_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1  g0306(.A1(new_n606_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n608_));
  NAND3_X1  g0307(.A1(new_n604_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n609_));
  NAND3_X1  g0308(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n610_));
  NAND4_X1  g0309(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .A4(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g0310(.A(G218), .B(G226), .ZN(new_n612_));
  XNOR2_X1  g0311(.A(G206), .B(G210), .ZN(new_n613_));
  XNOR2_X1  g0312(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g0313(.A(new_n611_), .B(new_n614_), .ZN(G1004));
  NAND2_X1  g0314(.A1(new_n519_), .A2(G457), .ZN(new_n616_));
  NOR2_X1   g0315(.A1(new_n509_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g0316(.A(new_n504_), .ZN(new_n618_));
  NOR2_X1   g0317(.A1(new_n618_), .A2(new_n421_), .ZN(new_n619_));
  NAND3_X1  g0318(.A1(new_n517_), .A2(new_n520_), .A3(new_n619_), .ZN(new_n620_));
  NOR2_X1   g0319(.A1(new_n513_), .A2(new_n414_), .ZN(new_n621_));
  NAND2_X1  g0320(.A1(new_n520_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g0321(.A(new_n509_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  AOI211_X1 g0322(.A(new_n617_), .B(new_n623_), .C1(G446), .C2(new_n508_), .ZN(new_n624_));
  AOI21_X1  g0323(.A(new_n443_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n625_));
  INV_X1    g0324(.A(new_n625_), .ZN(new_n626_));
  NOR3_X1   g0325(.A1(new_n480_), .A2(new_n490_), .A3(new_n626_), .ZN(new_n627_));
  NAND3_X1  g0326(.A1(new_n627_), .A2(new_n496_), .A3(new_n584_), .ZN(new_n628_));
  NAND2_X1  g0327(.A1(new_n489_), .A2(G435), .ZN(new_n629_));
  NAND3_X1  g0328(.A1(new_n479_), .A2(G400), .A3(new_n582_), .ZN(new_n630_));
  INV_X1    g0329(.A(new_n630_), .ZN(new_n631_));
  NAND2_X1  g0330(.A1(new_n631_), .A2(new_n581_), .ZN(new_n632_));
  NAND2_X1  g0331(.A1(new_n484_), .A2(G273), .ZN(new_n633_));
  AOI21_X1  g0332(.A(new_n450_), .B1(new_n633_), .B2(new_n492_), .ZN(new_n634_));
  NAND4_X1  g0333(.A1(new_n581_), .A2(new_n479_), .A3(new_n584_), .A4(new_n634_), .ZN(new_n635_));
  NAND4_X1  g0334(.A1(new_n628_), .A2(new_n629_), .A3(new_n632_), .A4(new_n635_), .ZN(new_n636_));
  NAND2_X1  g0335(.A1(new_n478_), .A2(G389), .ZN(new_n637_));
  NOR2_X1   g0336(.A1(new_n490_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g0337(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g0338(.A(new_n624_), .B1(new_n639_), .B2(new_n521_), .ZN(G591));
  INV_X1    g0339(.A(new_n544_), .ZN(new_n641_));
  INV_X1    g0340(.A(new_n526_), .ZN(new_n642_));
  INV_X1    g0341(.A(G490), .ZN(new_n643_));
  NOR2_X1   g0342(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g0343(.A(new_n644_), .ZN(new_n645_));
  NOR3_X1   g0344(.A1(new_n641_), .A2(new_n531_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g0345(.A1(new_n539_), .A2(G479), .ZN(new_n647_));
  NOR2_X1   g0346(.A1(new_n647_), .A2(new_n531_), .ZN(new_n648_));
  NOR4_X1   g0347(.A1(new_n646_), .A2(new_n531_), .A3(new_n535_), .A4(new_n648_), .ZN(new_n649_));
  NOR3_X1   g0348(.A1(new_n548_), .A2(new_n576_), .A3(new_n574_), .ZN(new_n650_));
  NAND3_X1  g0349(.A1(new_n650_), .A2(new_n559_), .A3(new_n565_), .ZN(new_n651_));
  NAND2_X1  g0350(.A1(new_n556_), .A2(G523), .ZN(new_n652_));
  INV_X1    g0351(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g0352(.A1(new_n653_), .A2(new_n553_), .ZN(new_n654_));
  INV_X1    g0353(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g0354(.A1(new_n655_), .A2(new_n549_), .ZN(new_n656_));
  AOI21_X1  g0355(.A(new_n392_), .B1(new_n563_), .B2(new_n560_), .ZN(new_n657_));
  NAND4_X1  g0356(.A1(new_n549_), .A2(new_n553_), .A3(new_n559_), .A4(new_n657_), .ZN(new_n658_));
  NAND2_X1  g0357(.A1(new_n547_), .A2(G503), .ZN(new_n659_));
  NAND4_X1  g0358(.A1(new_n651_), .A2(new_n656_), .A3(new_n658_), .A4(new_n659_), .ZN(new_n660_));
  NAND2_X1  g0359(.A1(new_n550_), .A2(G514), .ZN(new_n661_));
  NOR2_X1   g0360(.A1(new_n548_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g0361(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g0362(.A(new_n649_), .B1(new_n663_), .B2(new_n545_), .ZN(G618));
  OAI21_X1  g0363(.A(new_n624_), .B1(new_n639_), .B2(new_n580_), .ZN(G621));
  OAI21_X1  g0364(.A(new_n649_), .B1(new_n663_), .B2(new_n578_), .ZN(G629));
  XNOR2_X1  g0365(.A(new_n569_), .B(G54), .ZN(new_n667_));
  INV_X1    g0366(.A(G4092), .ZN(new_n668_));
  NAND3_X1  g0367(.A1(new_n667_), .A2(G4091), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g0368(.A(G4091), .ZN(new_n670_));
  NAND3_X1  g0369(.A1(new_n670_), .A2(G131), .A3(G4092), .ZN(new_n671_));
  NAND3_X1  g0370(.A1(new_n409_), .A2(new_n670_), .A3(new_n668_), .ZN(new_n672_));
  AND3_X1   g0371(.A1(new_n669_), .A2(new_n671_), .A3(new_n672_), .ZN(G822));
  OR2_X1    g0372(.A1(new_n569_), .A2(G54), .ZN(new_n674_));
  XOR2_X1   g0373(.A(new_n565_), .B(new_n674_), .Z(new_n675_));
  NAND3_X1  g0374(.A1(new_n675_), .A2(G4091), .A3(new_n668_), .ZN(new_n676_));
  NAND3_X1  g0375(.A1(new_n670_), .A2(G129), .A3(G4092), .ZN(new_n677_));
  OR3_X1    g0376(.A1(new_n395_), .A2(G4091), .A3(G4092), .ZN(new_n678_));
  AND3_X1   g0377(.A1(new_n676_), .A2(new_n677_), .A3(new_n678_), .ZN(G838));
  XNOR2_X1  g0378(.A(new_n500_), .B(G4), .ZN(new_n680_));
  NOR3_X1   g0379(.A1(new_n680_), .A2(new_n670_), .A3(G4092), .ZN(new_n681_));
  OR2_X1    g0380(.A1(new_n446_), .A2(G4092), .ZN(new_n682_));
  NAND2_X1  g0381(.A1(G117), .A2(G4092), .ZN(new_n683_));
  AOI21_X1  g0382(.A(G4091), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g0383(.A1(new_n681_), .A2(new_n684_), .ZN(G861));
  NOR2_X1   g0384(.A1(new_n566_), .A2(new_n569_), .ZN(new_n686_));
  NAND2_X1  g0385(.A1(new_n686_), .A2(G54), .ZN(new_n687_));
  NAND2_X1  g0386(.A1(new_n663_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g0387(.A(new_n688_), .ZN(new_n689_));
  NOR3_X1   g0388(.A1(new_n646_), .A2(new_n531_), .A3(new_n648_), .ZN(new_n690_));
  XNOR2_X1  g0389(.A(new_n690_), .B(new_n536_), .ZN(new_n691_));
  NAND2_X1  g0390(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g0391(.A(new_n544_), .B(new_n532_), .C1(G490), .C2(new_n526_), .ZN(new_n693_));
  NAND3_X1  g0392(.A1(new_n693_), .A2(new_n532_), .A3(new_n647_), .ZN(new_n694_));
  XNOR2_X1  g0393(.A(new_n694_), .B(new_n535_), .ZN(new_n695_));
  NAND2_X1  g0394(.A1(new_n688_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g0395(.A1(new_n692_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g0396(.A(new_n697_), .ZN(G623));
  INV_X1    g0397(.A(G861), .ZN(new_n699_));
  INV_X1    g0398(.A(G4087), .ZN(new_n700_));
  NAND3_X1  g0399(.A1(new_n699_), .A2(new_n700_), .A3(G4088), .ZN(new_n701_));
  OR3_X1    g0400(.A1(G822), .A2(G4087), .A3(G4088), .ZN(new_n702_));
  NAND3_X1  g0401(.A1(G61), .A2(G4087), .A3(G4088), .ZN(new_n703_));
  INV_X1    g0402(.A(G4088), .ZN(new_n704_));
  NAND3_X1  g0403(.A1(new_n704_), .A2(G11), .A3(G4087), .ZN(new_n705_));
  NAND4_X1  g0404(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .A4(new_n705_), .ZN(G722));
  INV_X1    g0405(.A(new_n565_), .ZN(new_n707_));
  NOR3_X1   g0406(.A1(new_n707_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n708_));
  NAND3_X1  g0407(.A1(new_n708_), .A2(G54), .A3(new_n576_), .ZN(new_n709_));
  NAND3_X1  g0408(.A1(new_n559_), .A2(new_n553_), .A3(new_n657_), .ZN(new_n710_));
  NAND4_X1  g0409(.A1(new_n559_), .A2(new_n565_), .A3(new_n553_), .A4(new_n569_), .ZN(new_n711_));
  NAND4_X1  g0410(.A1(new_n709_), .A2(new_n661_), .A3(new_n710_), .A4(new_n711_), .ZN(new_n712_));
  NOR2_X1   g0411(.A1(new_n712_), .A2(new_n655_), .ZN(new_n713_));
  XNOR2_X1  g0412(.A(new_n713_), .B(new_n548_), .ZN(new_n714_));
  NOR3_X1   g0413(.A1(new_n714_), .A2(new_n670_), .A3(G4092), .ZN(new_n715_));
  OR2_X1    g0414(.A1(new_n402_), .A2(G4092), .ZN(new_n716_));
  NAND2_X1  g0415(.A1(G52), .A2(G4092), .ZN(new_n717_));
  AOI21_X1  g0416(.A(G4091), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NOR2_X1   g0417(.A1(new_n715_), .A2(new_n718_), .ZN(G832));
  OAI211_X1 g0418(.A(new_n559_), .B(new_n565_), .C1(G54), .C2(new_n569_), .ZN(new_n720_));
  OAI21_X1  g0419(.A(new_n657_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n721_));
  NAND3_X1  g0420(.A1(new_n720_), .A2(new_n652_), .A3(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g0421(.A(new_n722_), .B(new_n553_), .ZN(new_n723_));
  NOR3_X1   g0422(.A1(new_n723_), .A2(new_n670_), .A3(G4092), .ZN(new_n724_));
  OR2_X1    g0423(.A1(new_n405_), .A2(G4092), .ZN(new_n725_));
  NAND2_X1  g0424(.A1(G130), .A2(G4092), .ZN(new_n726_));
  AOI21_X1  g0425(.A(G4091), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NOR2_X1   g0426(.A1(new_n724_), .A2(new_n727_), .ZN(G834));
  NAND3_X1  g0427(.A1(new_n565_), .A2(G54), .A3(new_n576_), .ZN(new_n729_));
  INV_X1    g0428(.A(new_n657_), .ZN(new_n730_));
  INV_X1    g0429(.A(new_n564_), .ZN(new_n731_));
  AOI21_X1  g0430(.A(G534), .B1(new_n563_), .B2(new_n560_), .ZN(new_n732_));
  OAI21_X1  g0431(.A(new_n569_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g0432(.A1(new_n729_), .A2(new_n730_), .A3(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g0433(.A(new_n734_), .B(new_n559_), .ZN(new_n735_));
  NOR3_X1   g0434(.A1(new_n735_), .A2(new_n670_), .A3(G4092), .ZN(new_n736_));
  OR2_X1    g0435(.A1(new_n388_), .A2(G4092), .ZN(new_n737_));
  NAND2_X1  g0436(.A1(G119), .A2(G4092), .ZN(new_n738_));
  AOI21_X1  g0437(.A(G4091), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g0438(.A1(new_n736_), .A2(new_n739_), .ZN(G836));
  INV_X1    g0439(.A(G4090), .ZN(new_n741_));
  NAND3_X1  g0440(.A1(new_n699_), .A2(G4089), .A3(new_n741_), .ZN(new_n742_));
  OR3_X1    g0441(.A1(G822), .A2(G4089), .A3(G4090), .ZN(new_n743_));
  NAND3_X1  g0442(.A1(G61), .A2(G4089), .A3(G4090), .ZN(new_n744_));
  INV_X1    g0443(.A(G4089), .ZN(new_n745_));
  NAND3_X1  g0444(.A1(new_n745_), .A2(G11), .A3(G4090), .ZN(new_n746_));
  NAND4_X1  g0445(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .A4(new_n746_), .ZN(G859));
  NAND3_X1  g0446(.A1(new_n479_), .A2(new_n584_), .A3(new_n634_), .ZN(new_n748_));
  NAND4_X1  g0447(.A1(new_n479_), .A2(new_n496_), .A3(new_n584_), .A4(new_n625_), .ZN(new_n749_));
  NAND4_X1  g0448(.A1(new_n479_), .A2(G4), .A3(new_n496_), .A4(new_n584_), .ZN(new_n750_));
  OAI211_X1 g0449(.A(new_n748_), .B(new_n749_), .C1(new_n750_), .C2(new_n586_), .ZN(new_n751_));
  INV_X1    g0450(.A(new_n751_), .ZN(new_n752_));
  NAND3_X1  g0451(.A1(new_n752_), .A2(new_n637_), .A3(new_n630_), .ZN(new_n753_));
  XNOR2_X1  g0452(.A(new_n753_), .B(new_n581_), .ZN(new_n754_));
  NOR3_X1   g0453(.A1(new_n754_), .A2(new_n670_), .A3(G4092), .ZN(new_n755_));
  OR2_X1    g0454(.A1(new_n431_), .A2(G4092), .ZN(new_n756_));
  NAND2_X1  g0455(.A1(G122), .A2(G4092), .ZN(new_n757_));
  AOI21_X1  g0456(.A(G4091), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g0457(.A1(new_n755_), .A2(new_n758_), .ZN(G871));
  NAND4_X1  g0458(.A1(new_n500_), .A2(G4), .A3(new_n496_), .A4(new_n584_), .ZN(new_n760_));
  NAND2_X1  g0459(.A1(new_n582_), .A2(G400), .ZN(new_n761_));
  OAI21_X1  g0460(.A(new_n634_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n762_));
  NAND3_X1  g0461(.A1(new_n496_), .A2(new_n584_), .A3(new_n625_), .ZN(new_n763_));
  NAND4_X1  g0462(.A1(new_n760_), .A2(new_n761_), .A3(new_n762_), .A4(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g0463(.A(new_n764_), .B(new_n479_), .ZN(new_n765_));
  NOR3_X1   g0464(.A1(new_n765_), .A2(new_n670_), .A3(G4092), .ZN(new_n766_));
  NOR2_X1   g0465(.A1(new_n460_), .A2(G4092), .ZN(new_n767_));
  INV_X1    g0466(.A(new_n767_), .ZN(new_n768_));
  NAND2_X1  g0467(.A1(G128), .A2(G4092), .ZN(new_n769_));
  AOI21_X1  g0468(.A(G4091), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g0469(.A1(new_n766_), .A2(new_n770_), .ZN(G873));
  NAND3_X1  g0470(.A1(new_n500_), .A2(G4), .A3(new_n496_), .ZN(new_n772_));
  INV_X1    g0471(.A(new_n634_), .ZN(new_n773_));
  INV_X1    g0472(.A(new_n495_), .ZN(new_n774_));
  AOI21_X1  g0473(.A(G411), .B1(new_n633_), .B2(new_n492_), .ZN(new_n775_));
  OAI21_X1  g0474(.A(new_n625_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g0475(.A1(new_n772_), .A2(new_n773_), .A3(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g0476(.A(new_n777_), .B(new_n584_), .ZN(new_n778_));
  NOR3_X1   g0477(.A1(new_n778_), .A2(new_n670_), .A3(G4092), .ZN(new_n779_));
  OR2_X1    g0478(.A1(new_n467_), .A2(G4092), .ZN(new_n780_));
  NAND2_X1  g0479(.A1(G127), .A2(G4092), .ZN(new_n781_));
  AOI21_X1  g0480(.A(G4091), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g0481(.A1(new_n779_), .A2(new_n782_), .ZN(G875));
  AOI21_X1  g0482(.A(new_n625_), .B1(new_n500_), .B2(G4), .ZN(new_n784_));
  INV_X1    g0483(.A(new_n496_), .ZN(new_n785_));
  XNOR2_X1  g0484(.A(new_n784_), .B(new_n785_), .ZN(new_n786_));
  NOR3_X1   g0485(.A1(new_n786_), .A2(new_n670_), .A3(G4092), .ZN(new_n787_));
  OR2_X1    g0486(.A1(new_n453_), .A2(G4092), .ZN(new_n788_));
  NAND2_X1  g0487(.A1(G126), .A2(G4092), .ZN(new_n789_));
  AOI21_X1  g0488(.A(G4091), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g0489(.A1(new_n787_), .A2(new_n790_), .ZN(G877));
  MUX2_X1   g0490(.A(G369), .B(G372), .S(G332), .Z(new_n792_));
  XNOR2_X1  g0491(.A(new_n792_), .B(new_n569_), .ZN(new_n793_));
  XOR2_X1   g0492(.A(new_n556_), .B(new_n561_), .Z(new_n794_));
  XNOR2_X1  g0493(.A(new_n547_), .B(new_n550_), .ZN(new_n795_));
  INV_X1    g0494(.A(new_n795_), .ZN(new_n796_));
  NOR3_X1   g0495(.A1(new_n793_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  NOR2_X1   g0496(.A1(new_n793_), .A2(new_n795_), .ZN(new_n798_));
  AOI21_X1  g0497(.A(new_n797_), .B1(new_n794_), .B2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g0498(.A1(new_n794_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n800_));
  NAND2_X1  g0499(.A1(new_n793_), .A2(new_n796_), .ZN(new_n801_));
  OAI211_X1 g0500(.A(new_n799_), .B(new_n800_), .C1(new_n794_), .C2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g0501(.A(new_n526_), .B(new_n539_), .ZN(new_n803_));
  XNOR2_X1  g0502(.A(new_n531_), .B(new_n535_), .ZN(new_n804_));
  XNOR2_X1  g0503(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g0504(.A(new_n802_), .B(new_n805_), .ZN(G998));
  MUX2_X1   g0505(.A(G289), .B(G292), .S(G335), .Z(new_n807_));
  XNOR2_X1  g0506(.A(new_n807_), .B(new_n508_), .ZN(new_n808_));
  INV_X1    g0507(.A(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g0508(.A(new_n515_), .B(new_n519_), .ZN(new_n810_));
  XNOR2_X1  g0509(.A(new_n504_), .B(new_n489_), .ZN(new_n811_));
  NAND3_X1  g0510(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g0511(.A(new_n810_), .ZN(new_n813_));
  INV_X1    g0512(.A(new_n811_), .ZN(new_n814_));
  NAND3_X1  g0513(.A1(new_n809_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g0514(.A1(new_n814_), .A2(new_n808_), .A3(new_n810_), .ZN(new_n816_));
  NAND3_X1  g0515(.A1(new_n813_), .A2(new_n808_), .A3(new_n811_), .ZN(new_n817_));
  NAND4_X1  g0516(.A1(new_n812_), .A2(new_n815_), .A3(new_n816_), .A4(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g0517(.A(new_n499_), .B(new_n493_), .ZN(new_n819_));
  XNOR2_X1  g0518(.A(new_n582_), .B(new_n478_), .ZN(new_n820_));
  XNOR2_X1  g0519(.A(new_n819_), .B(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g0520(.A(new_n818_), .B(new_n821_), .ZN(G1000));
  NOR2_X1   g0521(.A1(new_n585_), .A2(new_n586_), .ZN(new_n823_));
  NAND2_X1  g0522(.A1(new_n823_), .A2(G4), .ZN(new_n824_));
  NAND2_X1  g0523(.A1(new_n639_), .A2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g0524(.A(new_n825_), .B(new_n506_), .ZN(new_n826_));
  INV_X1    g0525(.A(new_n826_), .ZN(new_n827_));
  INV_X1    g0526(.A(new_n825_), .ZN(new_n828_));
  XOR2_X1   g0527(.A(new_n517_), .B(new_n619_), .Z(new_n829_));
  NAND2_X1  g0528(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g0529(.A1(new_n618_), .A2(new_n421_), .ZN(new_n831_));
  XNOR2_X1  g0530(.A(new_n517_), .B(new_n831_), .ZN(new_n832_));
  OAI21_X1  g0531(.A(new_n830_), .B1(new_n828_), .B2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g0532(.A1(new_n620_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n834_));
  XNOR2_X1  g0533(.A(new_n834_), .B(new_n509_), .ZN(new_n835_));
  NAND2_X1  g0534(.A1(new_n828_), .A2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g0535(.A(new_n517_), .B(new_n520_), .C1(G422), .C2(new_n504_), .ZN(new_n837_));
  NAND3_X1  g0536(.A1(new_n837_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n838_));
  XNOR2_X1  g0537(.A(new_n838_), .B(new_n509_), .ZN(new_n839_));
  NAND2_X1  g0538(.A1(new_n825_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g0539(.A1(new_n836_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g0540(.A1(new_n517_), .A2(new_n619_), .ZN(new_n842_));
  INV_X1    g0541(.A(new_n621_), .ZN(new_n843_));
  NAND2_X1  g0542(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g0543(.A(new_n520_), .ZN(new_n845_));
  XNOR2_X1  g0544(.A(new_n844_), .B(new_n845_), .ZN(new_n846_));
  NAND2_X1  g0545(.A1(new_n828_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g0546(.A(new_n517_), .ZN(new_n848_));
  OAI211_X1 g0547(.A(new_n842_), .B(new_n843_), .C1(new_n848_), .C2(new_n505_), .ZN(new_n849_));
  XNOR2_X1  g0548(.A(new_n849_), .B(new_n845_), .ZN(new_n850_));
  NAND2_X1  g0549(.A1(new_n825_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g0550(.A1(new_n847_), .A2(new_n851_), .ZN(new_n852_));
  NOR4_X1   g0551(.A1(new_n827_), .A2(new_n833_), .A3(new_n841_), .A4(new_n852_), .ZN(new_n853_));
  AND4_X1   g0552(.A1(new_n754_), .A2(new_n853_), .A3(new_n765_), .A4(new_n778_), .ZN(new_n854_));
  AND3_X1   g0553(.A1(new_n854_), .A2(new_n680_), .A3(new_n786_), .ZN(G575));
  XNOR2_X1  g0554(.A(new_n688_), .B(new_n528_), .ZN(new_n856_));
  INV_X1    g0555(.A(new_n856_), .ZN(new_n857_));
  XNOR2_X1  g0556(.A(new_n544_), .B(new_n645_), .ZN(new_n858_));
  NAND2_X1  g0557(.A1(new_n689_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g0558(.A1(new_n642_), .A2(new_n643_), .ZN(new_n860_));
  XNOR2_X1  g0559(.A(new_n544_), .B(new_n860_), .ZN(new_n861_));
  OAI21_X1  g0560(.A(new_n859_), .B1(new_n689_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g0561(.A1(new_n544_), .A2(new_n644_), .ZN(new_n863_));
  NAND2_X1  g0562(.A1(new_n863_), .A2(new_n647_), .ZN(new_n864_));
  XNOR2_X1  g0563(.A(new_n864_), .B(new_n531_), .ZN(new_n865_));
  NAND2_X1  g0564(.A1(new_n689_), .A2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g0565(.A(new_n863_), .B(new_n647_), .C1(new_n641_), .C2(new_n527_), .ZN(new_n867_));
  XNOR2_X1  g0566(.A(new_n867_), .B(new_n531_), .ZN(new_n868_));
  NAND2_X1  g0567(.A1(new_n688_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g0568(.A1(new_n866_), .A2(new_n869_), .ZN(new_n870_));
  NOR4_X1   g0569(.A1(new_n857_), .A2(new_n862_), .A3(new_n697_), .A4(new_n870_), .ZN(new_n871_));
  NAND4_X1  g0570(.A1(new_n871_), .A2(new_n714_), .A3(new_n723_), .A4(new_n735_), .ZN(new_n872_));
  NOR3_X1   g0571(.A1(new_n872_), .A2(new_n667_), .A3(new_n675_), .ZN(G585));
  INV_X1    g0572(.A(G137), .ZN(new_n874_));
  INV_X1    g0573(.A(G1690), .ZN(new_n875_));
  NAND3_X1  g0574(.A1(new_n699_), .A2(G1689), .A3(new_n875_), .ZN(new_n876_));
  NAND3_X1  g0575(.A1(G185), .A2(G1689), .A3(G1690), .ZN(new_n877_));
  NAND2_X1  g0576(.A1(G182), .A2(G1690), .ZN(new_n878_));
  OAI21_X1  g0577(.A(new_n877_), .B1(new_n878_), .B2(G1689), .ZN(new_n879_));
  NOR2_X1   g0578(.A1(G822), .A2(G1690), .ZN(new_n880_));
  INV_X1    g0579(.A(G1689), .ZN(new_n881_));
  AOI21_X1  g0580(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g0581(.A(new_n874_), .B1(new_n876_), .B2(new_n882_), .ZN(G661));
  INV_X1    g0582(.A(G1694), .ZN(new_n884_));
  NAND3_X1  g0583(.A1(new_n699_), .A2(G1691), .A3(new_n884_), .ZN(new_n885_));
  NAND3_X1  g0584(.A1(G185), .A2(G1691), .A3(G1694), .ZN(new_n886_));
  NAND2_X1  g0585(.A1(G182), .A2(G1694), .ZN(new_n887_));
  OAI21_X1  g0586(.A(new_n886_), .B1(new_n887_), .B2(G1691), .ZN(new_n888_));
  NOR2_X1   g0587(.A1(G822), .A2(G1694), .ZN(new_n889_));
  INV_X1    g0588(.A(G1691), .ZN(new_n890_));
  AOI21_X1  g0589(.A(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g0590(.A(new_n874_), .B1(new_n885_), .B2(new_n891_), .ZN(G693));
  INV_X1    g0591(.A(G832), .ZN(new_n893_));
  NAND3_X1  g0592(.A1(new_n893_), .A2(new_n700_), .A3(new_n704_), .ZN(new_n894_));
  INV_X1    g0593(.A(G871), .ZN(new_n895_));
  NAND3_X1  g0594(.A1(new_n895_), .A2(new_n700_), .A3(G4088), .ZN(new_n896_));
  NAND3_X1  g0595(.A1(G37), .A2(G4087), .A3(G4088), .ZN(new_n897_));
  NAND3_X1  g0596(.A1(new_n704_), .A2(G43), .A3(G4087), .ZN(new_n898_));
  NAND4_X1  g0597(.A1(new_n894_), .A2(new_n896_), .A3(new_n897_), .A4(new_n898_), .ZN(G747));
  INV_X1    g0598(.A(G873), .ZN(new_n900_));
  NAND3_X1  g0599(.A1(new_n900_), .A2(new_n700_), .A3(G4088), .ZN(new_n901_));
  INV_X1    g0600(.A(G834), .ZN(new_n902_));
  NAND3_X1  g0601(.A1(new_n902_), .A2(new_n700_), .A3(new_n704_), .ZN(new_n903_));
  NAND3_X1  g0602(.A1(G20), .A2(G4087), .A3(G4088), .ZN(new_n904_));
  NAND3_X1  g0603(.A1(new_n704_), .A2(G76), .A3(G4087), .ZN(new_n905_));
  NAND4_X1  g0604(.A1(new_n901_), .A2(new_n903_), .A3(new_n904_), .A4(new_n905_), .ZN(G752));
  INV_X1    g0605(.A(G875), .ZN(new_n907_));
  NAND3_X1  g0606(.A1(new_n907_), .A2(new_n700_), .A3(G4088), .ZN(new_n908_));
  INV_X1    g0607(.A(G836), .ZN(new_n909_));
  NAND3_X1  g0608(.A1(new_n909_), .A2(new_n700_), .A3(new_n704_), .ZN(new_n910_));
  NAND3_X1  g0609(.A1(G17), .A2(G4087), .A3(G4088), .ZN(new_n911_));
  NAND3_X1  g0610(.A1(new_n704_), .A2(G73), .A3(G4087), .ZN(new_n912_));
  NAND4_X1  g0611(.A1(new_n908_), .A2(new_n910_), .A3(new_n911_), .A4(new_n912_), .ZN(G757));
  INV_X1    g0612(.A(G877), .ZN(new_n914_));
  NAND3_X1  g0613(.A1(new_n914_), .A2(new_n700_), .A3(G4088), .ZN(new_n915_));
  OR3_X1    g0614(.A1(G838), .A2(G4087), .A3(G4088), .ZN(new_n916_));
  NAND3_X1  g0615(.A1(G70), .A2(G4087), .A3(G4088), .ZN(new_n917_));
  NAND3_X1  g0616(.A1(new_n704_), .A2(G67), .A3(G4087), .ZN(new_n918_));
  NAND4_X1  g0617(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .A4(new_n918_), .ZN(G762));
  NAND3_X1  g0618(.A1(new_n893_), .A2(new_n745_), .A3(new_n741_), .ZN(new_n920_));
  NAND3_X1  g0619(.A1(new_n895_), .A2(G4089), .A3(new_n741_), .ZN(new_n921_));
  NAND3_X1  g0620(.A1(G37), .A2(G4089), .A3(G4090), .ZN(new_n922_));
  NAND3_X1  g0621(.A1(new_n745_), .A2(G43), .A3(G4090), .ZN(new_n923_));
  NAND4_X1  g0622(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .A4(new_n923_), .ZN(G787));
  NAND3_X1  g0623(.A1(new_n900_), .A2(G4089), .A3(new_n741_), .ZN(new_n925_));
  NAND3_X1  g0624(.A1(new_n902_), .A2(new_n745_), .A3(new_n741_), .ZN(new_n926_));
  NAND3_X1  g0625(.A1(G20), .A2(G4089), .A3(G4090), .ZN(new_n927_));
  NAND3_X1  g0626(.A1(new_n745_), .A2(G76), .A3(G4090), .ZN(new_n928_));
  NAND4_X1  g0627(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .A4(new_n928_), .ZN(G792));
  NAND3_X1  g0628(.A1(new_n907_), .A2(G4089), .A3(new_n741_), .ZN(new_n930_));
  NAND3_X1  g0629(.A1(new_n909_), .A2(new_n745_), .A3(new_n741_), .ZN(new_n931_));
  NAND3_X1  g0630(.A1(G17), .A2(G4089), .A3(G4090), .ZN(new_n932_));
  NAND3_X1  g0631(.A1(new_n745_), .A2(G73), .A3(G4090), .ZN(new_n933_));
  NAND4_X1  g0632(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .A4(new_n933_), .ZN(G797));
  NAND3_X1  g0633(.A1(new_n914_), .A2(G4089), .A3(new_n741_), .ZN(new_n935_));
  OR3_X1    g0634(.A1(G838), .A2(G4089), .A3(G4090), .ZN(new_n936_));
  NAND3_X1  g0635(.A1(G70), .A2(G4089), .A3(G4090), .ZN(new_n937_));
  NAND3_X1  g0636(.A1(new_n745_), .A2(G67), .A3(G4090), .ZN(new_n938_));
  NAND4_X1  g0637(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .A4(new_n938_), .ZN(G802));
  NAND3_X1  g0638(.A1(G170), .A2(G1689), .A3(G1690), .ZN(new_n940_));
  NAND2_X1  g0639(.A1(G200), .A2(G1690), .ZN(new_n941_));
  OAI21_X1  g0640(.A(new_n940_), .B1(new_n941_), .B2(G1689), .ZN(new_n942_));
  NOR2_X1   g0641(.A1(G832), .A2(G1690), .ZN(new_n943_));
  AOI21_X1  g0642(.A(new_n942_), .B1(new_n943_), .B2(new_n881_), .ZN(new_n944_));
  NAND3_X1  g0643(.A1(new_n895_), .A2(G1689), .A3(new_n875_), .ZN(new_n945_));
  AOI21_X1  g0644(.A(new_n874_), .B1(new_n944_), .B2(new_n945_), .ZN(G642));
  NAND3_X1  g0645(.A1(new_n914_), .A2(G1689), .A3(new_n875_), .ZN(new_n947_));
  NAND3_X1  g0646(.A1(G158), .A2(G1689), .A3(G1690), .ZN(new_n948_));
  NAND2_X1  g0647(.A1(G188), .A2(G1690), .ZN(new_n949_));
  OAI21_X1  g0648(.A(new_n948_), .B1(new_n949_), .B2(G1689), .ZN(new_n950_));
  NOR2_X1   g0649(.A1(G838), .A2(G1690), .ZN(new_n951_));
  AOI21_X1  g0650(.A(new_n950_), .B1(new_n951_), .B2(new_n881_), .ZN(new_n952_));
  AOI21_X1  g0651(.A(new_n874_), .B1(new_n947_), .B2(new_n952_), .ZN(G664));
  NAND3_X1  g0652(.A1(new_n907_), .A2(G1689), .A3(new_n875_), .ZN(new_n954_));
  NAND3_X1  g0653(.A1(G152), .A2(G1689), .A3(G1690), .ZN(new_n955_));
  NAND2_X1  g0654(.A1(G155), .A2(G1690), .ZN(new_n956_));
  OAI21_X1  g0655(.A(new_n955_), .B1(new_n956_), .B2(G1689), .ZN(new_n957_));
  NOR2_X1   g0656(.A1(G836), .A2(G1690), .ZN(new_n958_));
  AOI21_X1  g0657(.A(new_n957_), .B1(new_n958_), .B2(new_n881_), .ZN(new_n959_));
  AOI21_X1  g0658(.A(new_n874_), .B1(new_n954_), .B2(new_n959_), .ZN(G667));
  NAND3_X1  g0659(.A1(G146), .A2(G1689), .A3(G1690), .ZN(new_n961_));
  NAND2_X1  g0660(.A1(G149), .A2(G1690), .ZN(new_n962_));
  OAI21_X1  g0661(.A(new_n961_), .B1(new_n962_), .B2(G1689), .ZN(new_n963_));
  NOR2_X1   g0662(.A1(G834), .A2(G1690), .ZN(new_n964_));
  AOI21_X1  g0663(.A(new_n963_), .B1(new_n964_), .B2(new_n881_), .ZN(new_n965_));
  NAND3_X1  g0664(.A1(new_n900_), .A2(G1689), .A3(new_n875_), .ZN(new_n966_));
  AOI21_X1  g0665(.A(new_n874_), .B1(new_n965_), .B2(new_n966_), .ZN(G670));
  NAND3_X1  g0666(.A1(G170), .A2(G1691), .A3(G1694), .ZN(new_n968_));
  NAND2_X1  g0667(.A1(G200), .A2(G1694), .ZN(new_n969_));
  OAI21_X1  g0668(.A(new_n968_), .B1(new_n969_), .B2(G1691), .ZN(new_n970_));
  NOR2_X1   g0669(.A1(G832), .A2(G1694), .ZN(new_n971_));
  AOI21_X1  g0670(.A(new_n970_), .B1(new_n971_), .B2(new_n890_), .ZN(new_n972_));
  NAND3_X1  g0671(.A1(new_n895_), .A2(G1691), .A3(new_n884_), .ZN(new_n973_));
  AOI21_X1  g0672(.A(new_n874_), .B1(new_n972_), .B2(new_n973_), .ZN(G676));
  NAND3_X1  g0673(.A1(new_n914_), .A2(G1691), .A3(new_n884_), .ZN(new_n975_));
  NAND3_X1  g0674(.A1(G158), .A2(G1691), .A3(G1694), .ZN(new_n976_));
  NAND2_X1  g0675(.A1(G188), .A2(G1694), .ZN(new_n977_));
  OAI21_X1  g0676(.A(new_n976_), .B1(new_n977_), .B2(G1691), .ZN(new_n978_));
  NOR2_X1   g0677(.A1(G838), .A2(G1694), .ZN(new_n979_));
  AOI21_X1  g0678(.A(new_n978_), .B1(new_n979_), .B2(new_n890_), .ZN(new_n980_));
  AOI21_X1  g0679(.A(new_n874_), .B1(new_n975_), .B2(new_n980_), .ZN(G696));
  NAND3_X1  g0680(.A1(new_n907_), .A2(G1691), .A3(new_n884_), .ZN(new_n982_));
  NAND3_X1  g0681(.A1(G152), .A2(G1691), .A3(G1694), .ZN(new_n983_));
  NAND2_X1  g0682(.A1(G155), .A2(G1694), .ZN(new_n984_));
  OAI21_X1  g0683(.A(new_n983_), .B1(new_n984_), .B2(G1691), .ZN(new_n985_));
  NOR2_X1   g0684(.A1(G836), .A2(G1694), .ZN(new_n986_));
  AOI21_X1  g0685(.A(new_n985_), .B1(new_n986_), .B2(new_n890_), .ZN(new_n987_));
  AOI21_X1  g0686(.A(new_n874_), .B1(new_n982_), .B2(new_n987_), .ZN(G699));
  NAND3_X1  g0687(.A1(G146), .A2(G1691), .A3(G1694), .ZN(new_n989_));
  NAND2_X1  g0688(.A1(G149), .A2(G1694), .ZN(new_n990_));
  OAI21_X1  g0689(.A(new_n989_), .B1(new_n990_), .B2(G1691), .ZN(new_n991_));
  NOR2_X1   g0690(.A1(G834), .A2(G1694), .ZN(new_n992_));
  AOI21_X1  g0691(.A(new_n991_), .B1(new_n992_), .B2(new_n890_), .ZN(new_n993_));
  NAND3_X1  g0692(.A1(new_n900_), .A2(G1691), .A3(new_n884_), .ZN(new_n994_));
  AOI21_X1  g0693(.A(new_n874_), .B1(new_n993_), .B2(new_n994_), .ZN(G702));
  NAND3_X1  g0694(.A1(new_n697_), .A2(G3717), .A3(G3724), .ZN(new_n996_));
  INV_X1    g0695(.A(G3717), .ZN(new_n997_));
  INV_X1    g0696(.A(G3724), .ZN(new_n998_));
  NAND3_X1  g0697(.A1(new_n365_), .A2(new_n997_), .A3(new_n998_), .ZN(new_n999_));
  NAND3_X1  g0698(.A1(new_n998_), .A2(G123), .A3(G3717), .ZN(new_n1000_));
  AND3_X1   g0699(.A1(new_n996_), .A2(new_n999_), .A3(new_n1000_), .ZN(new_n1001_));
  XNOR2_X1  g0700(.A(new_n535_), .B(G132), .ZN(new_n1002_));
  NAND3_X1  g0701(.A1(new_n1002_), .A2(new_n997_), .A3(G3724), .ZN(new_n1003_));
  AOI22_X1  g0702(.A1(new_n1001_), .A2(new_n1003_), .B1(G135), .B2(G4115), .ZN(G818));
  XOR2_X1   g0703(.A(new_n697_), .B(new_n1002_), .Z(G813));
  NOR3_X1   g0704(.A1(G623), .A2(new_n670_), .A3(G4092), .ZN(new_n1006_));
  NAND2_X1  g0705(.A1(new_n365_), .A2(new_n668_), .ZN(new_n1007_));
  NAND2_X1  g0706(.A1(G123), .A2(G4092), .ZN(new_n1008_));
  AOI21_X1  g0707(.A(G4091), .B1(new_n1007_), .B2(new_n1008_), .ZN(new_n1009_));
  NOR2_X1   g0708(.A1(new_n1006_), .A2(new_n1009_), .ZN(G824));
  AOI211_X1 g0709(.A(new_n670_), .B(G4092), .C1(new_n866_), .C2(new_n869_), .ZN(new_n1011_));
  NAND2_X1  g0710(.A1(new_n362_), .A2(new_n668_), .ZN(new_n1012_));
  NAND2_X1  g0711(.A1(G121), .A2(G4092), .ZN(new_n1013_));
  AOI21_X1  g0712(.A(G4091), .B1(new_n1012_), .B2(new_n1013_), .ZN(new_n1014_));
  NOR2_X1   g0713(.A1(new_n1011_), .A2(new_n1014_), .ZN(G826));
  AND3_X1   g0714(.A1(new_n862_), .A2(G4091), .A3(new_n668_), .ZN(new_n1016_));
  OR2_X1    g0715(.A1(new_n372_), .A2(G4092), .ZN(new_n1017_));
  NAND2_X1  g0716(.A1(G116), .A2(G4092), .ZN(new_n1018_));
  AOI21_X1  g0717(.A(G4091), .B1(new_n1017_), .B2(new_n1018_), .ZN(new_n1019_));
  NOR2_X1   g0718(.A1(new_n1016_), .A2(new_n1019_), .ZN(G828));
  NOR3_X1   g0719(.A1(new_n856_), .A2(new_n670_), .A3(G4092), .ZN(new_n1021_));
  OR2_X1    g0720(.A1(new_n378_), .A2(G4092), .ZN(new_n1022_));
  NAND2_X1  g0721(.A1(G112), .A2(G4092), .ZN(new_n1023_));
  AOI21_X1  g0722(.A(G4091), .B1(new_n1022_), .B2(new_n1023_), .ZN(new_n1024_));
  NOR2_X1   g0723(.A1(new_n1021_), .A2(new_n1024_), .ZN(G830));
  OR4_X1    g0724(.A1(G850), .A2(G1000), .A3(G1002), .A4(G1004), .ZN(new_n1026_));
  NAND4_X1  g0725(.A1(G386), .A2(G552), .A3(G556), .A4(G559), .ZN(new_n1027_));
  NOR4_X1   g0726(.A1(new_n1026_), .A2(G848), .A3(G998), .A4(new_n1027_), .ZN(G854));
  AOI211_X1 g0727(.A(new_n670_), .B(G4092), .C1(new_n836_), .C2(new_n840_), .ZN(new_n1029_));
  NAND2_X1  g0728(.A1(new_n475_), .A2(new_n668_), .ZN(new_n1030_));
  NAND2_X1  g0729(.A1(G115), .A2(G4092), .ZN(new_n1031_));
  AOI21_X1  g0730(.A(G4091), .B1(new_n1030_), .B2(new_n1031_), .ZN(new_n1032_));
  NOR2_X1   g0731(.A1(new_n1029_), .A2(new_n1032_), .ZN(G863));
  AOI211_X1 g0732(.A(new_n670_), .B(G4092), .C1(new_n847_), .C2(new_n851_), .ZN(new_n1034_));
  NOR2_X1   g0733(.A1(new_n438_), .A2(G4092), .ZN(new_n1035_));
  INV_X1    g0734(.A(new_n1035_), .ZN(new_n1036_));
  NAND2_X1  g0735(.A1(G114), .A2(G4092), .ZN(new_n1037_));
  AOI21_X1  g0736(.A(G4091), .B1(new_n1036_), .B2(new_n1037_), .ZN(new_n1038_));
  NOR2_X1   g0737(.A1(new_n1034_), .A2(new_n1038_), .ZN(G865));
  AND3_X1   g0738(.A1(new_n833_), .A2(G4091), .A3(new_n668_), .ZN(new_n1040_));
  NOR2_X1   g0739(.A1(new_n417_), .A2(G4092), .ZN(new_n1041_));
  INV_X1    g0740(.A(new_n1041_), .ZN(new_n1042_));
  NAND2_X1  g0741(.A1(G53), .A2(G4092), .ZN(new_n1043_));
  AOI21_X1  g0742(.A(G4091), .B1(new_n1042_), .B2(new_n1043_), .ZN(new_n1044_));
  NOR2_X1   g0743(.A1(new_n1040_), .A2(new_n1044_), .ZN(G867));
  NOR3_X1   g0744(.A1(new_n826_), .A2(new_n670_), .A3(G4092), .ZN(new_n1046_));
  NOR2_X1   g0745(.A1(new_n424_), .A2(G4092), .ZN(new_n1047_));
  INV_X1    g0746(.A(new_n1047_), .ZN(new_n1048_));
  NAND2_X1  g0747(.A1(G113), .A2(G4092), .ZN(new_n1049_));
  AOI21_X1  g0748(.A(G4091), .B1(new_n1048_), .B2(new_n1049_), .ZN(new_n1050_));
  NOR2_X1   g0749(.A1(new_n1046_), .A2(new_n1050_), .ZN(G869));
  INV_X1    g0750(.A(G824), .ZN(new_n1052_));
  NAND3_X1  g0751(.A1(new_n1052_), .A2(new_n745_), .A3(new_n741_), .ZN(new_n1053_));
  INV_X1    g0752(.A(G863), .ZN(new_n1054_));
  NAND3_X1  g0753(.A1(new_n1054_), .A2(G4089), .A3(new_n741_), .ZN(new_n1055_));
  NAND3_X1  g0754(.A1(G106), .A2(G4089), .A3(G4090), .ZN(new_n1056_));
  NAND3_X1  g0755(.A1(new_n745_), .A2(G109), .A3(G4090), .ZN(new_n1057_));
  NAND4_X1  g0756(.A1(new_n1053_), .A2(new_n1055_), .A3(new_n1056_), .A4(new_n1057_), .ZN(G712));
  NAND3_X1  g0757(.A1(new_n1052_), .A2(new_n700_), .A3(new_n704_), .ZN(new_n1059_));
  NAND3_X1  g0758(.A1(new_n1054_), .A2(new_n700_), .A3(G4088), .ZN(new_n1060_));
  NAND3_X1  g0759(.A1(G106), .A2(G4087), .A3(G4088), .ZN(new_n1061_));
  NAND3_X1  g0760(.A1(new_n704_), .A2(G109), .A3(G4087), .ZN(new_n1062_));
  NAND4_X1  g0761(.A1(new_n1059_), .A2(new_n1060_), .A3(new_n1061_), .A4(new_n1062_), .ZN(G727));
  INV_X1    g0762(.A(G865), .ZN(new_n1064_));
  NAND3_X1  g0763(.A1(new_n1064_), .A2(new_n700_), .A3(G4088), .ZN(new_n1065_));
  INV_X1    g0764(.A(G826), .ZN(new_n1066_));
  NAND3_X1  g0765(.A1(new_n1066_), .A2(new_n700_), .A3(new_n704_), .ZN(new_n1067_));
  NAND3_X1  g0766(.A1(G49), .A2(G4087), .A3(G4088), .ZN(new_n1068_));
  NAND3_X1  g0767(.A1(new_n704_), .A2(G46), .A3(G4087), .ZN(new_n1069_));
  NAND4_X1  g0768(.A1(new_n1065_), .A2(new_n1067_), .A3(new_n1068_), .A4(new_n1069_), .ZN(G732));
  INV_X1    g0769(.A(G867), .ZN(new_n1071_));
  NAND3_X1  g0770(.A1(new_n1071_), .A2(new_n700_), .A3(G4088), .ZN(new_n1072_));
  INV_X1    g0771(.A(G828), .ZN(new_n1073_));
  NAND3_X1  g0772(.A1(new_n1073_), .A2(new_n700_), .A3(new_n704_), .ZN(new_n1074_));
  NAND3_X1  g0773(.A1(G103), .A2(G4087), .A3(G4088), .ZN(new_n1075_));
  NAND3_X1  g0774(.A1(new_n704_), .A2(G100), .A3(G4087), .ZN(new_n1076_));
  NAND4_X1  g0775(.A1(new_n1072_), .A2(new_n1074_), .A3(new_n1075_), .A4(new_n1076_), .ZN(G737));
  INV_X1    g0776(.A(G869), .ZN(new_n1078_));
  NAND3_X1  g0777(.A1(new_n1078_), .A2(new_n700_), .A3(G4088), .ZN(new_n1079_));
  INV_X1    g0778(.A(G830), .ZN(new_n1080_));
  NAND3_X1  g0779(.A1(new_n1080_), .A2(new_n700_), .A3(new_n704_), .ZN(new_n1081_));
  NAND3_X1  g0780(.A1(G40), .A2(G4087), .A3(G4088), .ZN(new_n1082_));
  NAND3_X1  g0781(.A1(new_n704_), .A2(G91), .A3(G4087), .ZN(new_n1083_));
  NAND4_X1  g0782(.A1(new_n1079_), .A2(new_n1081_), .A3(new_n1082_), .A4(new_n1083_), .ZN(G742));
  NAND3_X1  g0783(.A1(new_n1064_), .A2(G4089), .A3(new_n741_), .ZN(new_n1085_));
  NAND3_X1  g0784(.A1(new_n1066_), .A2(new_n745_), .A3(new_n741_), .ZN(new_n1086_));
  NAND3_X1  g0785(.A1(G49), .A2(G4089), .A3(G4090), .ZN(new_n1087_));
  NAND3_X1  g0786(.A1(new_n745_), .A2(G46), .A3(G4090), .ZN(new_n1088_));
  NAND4_X1  g0787(.A1(new_n1085_), .A2(new_n1086_), .A3(new_n1087_), .A4(new_n1088_), .ZN(G772));
  NAND3_X1  g0788(.A1(new_n1071_), .A2(G4089), .A3(new_n741_), .ZN(new_n1090_));
  NAND3_X1  g0789(.A1(new_n1073_), .A2(new_n745_), .A3(new_n741_), .ZN(new_n1091_));
  NAND3_X1  g0790(.A1(G103), .A2(G4089), .A3(G4090), .ZN(new_n1092_));
  NAND3_X1  g0791(.A1(new_n745_), .A2(G100), .A3(G4090), .ZN(new_n1093_));
  NAND4_X1  g0792(.A1(new_n1090_), .A2(new_n1091_), .A3(new_n1092_), .A4(new_n1093_), .ZN(G777));
  NAND3_X1  g0793(.A1(new_n1078_), .A2(G4089), .A3(new_n741_), .ZN(new_n1095_));
  NAND3_X1  g0794(.A1(new_n1080_), .A2(new_n745_), .A3(new_n741_), .ZN(new_n1096_));
  NAND3_X1  g0795(.A1(G40), .A2(G4089), .A3(G4090), .ZN(new_n1097_));
  NAND3_X1  g0796(.A1(new_n745_), .A2(G91), .A3(G4090), .ZN(new_n1098_));
  NAND4_X1  g0797(.A1(new_n1095_), .A2(new_n1096_), .A3(new_n1097_), .A4(new_n1098_), .ZN(G782));
  NAND3_X1  g0798(.A1(new_n1078_), .A2(G1689), .A3(new_n875_), .ZN(new_n1100_));
  NAND3_X1  g0799(.A1(G173), .A2(G1689), .A3(G1690), .ZN(new_n1101_));
  NAND2_X1  g0800(.A1(G203), .A2(G1690), .ZN(new_n1102_));
  OAI21_X1  g0801(.A(new_n1101_), .B1(new_n1102_), .B2(G1689), .ZN(new_n1103_));
  NOR2_X1   g0802(.A1(G830), .A2(G1690), .ZN(new_n1104_));
  AOI21_X1  g0803(.A(new_n1103_), .B1(new_n1104_), .B2(new_n881_), .ZN(new_n1105_));
  AOI21_X1  g0804(.A(new_n874_), .B1(new_n1100_), .B2(new_n1105_), .ZN(G645));
  NAND3_X1  g0805(.A1(new_n1071_), .A2(G1689), .A3(new_n875_), .ZN(new_n1107_));
  NAND3_X1  g0806(.A1(G167), .A2(G1689), .A3(G1690), .ZN(new_n1108_));
  NAND2_X1  g0807(.A1(G197), .A2(G1690), .ZN(new_n1109_));
  OAI21_X1  g0808(.A(new_n1108_), .B1(new_n1109_), .B2(G1689), .ZN(new_n1110_));
  NOR2_X1   g0809(.A1(G828), .A2(G1690), .ZN(new_n1111_));
  AOI21_X1  g0810(.A(new_n1110_), .B1(new_n1111_), .B2(new_n881_), .ZN(new_n1112_));
  AOI21_X1  g0811(.A(new_n874_), .B1(new_n1107_), .B2(new_n1112_), .ZN(G648));
  NAND3_X1  g0812(.A1(new_n1064_), .A2(G1689), .A3(new_n875_), .ZN(new_n1114_));
  NAND3_X1  g0813(.A1(G164), .A2(G1689), .A3(G1690), .ZN(new_n1115_));
  NAND2_X1  g0814(.A1(G194), .A2(G1690), .ZN(new_n1116_));
  OAI21_X1  g0815(.A(new_n1115_), .B1(new_n1116_), .B2(G1689), .ZN(new_n1117_));
  NOR2_X1   g0816(.A1(G826), .A2(G1690), .ZN(new_n1118_));
  AOI21_X1  g0817(.A(new_n1117_), .B1(new_n1118_), .B2(new_n881_), .ZN(new_n1119_));
  AOI21_X1  g0818(.A(new_n874_), .B1(new_n1114_), .B2(new_n1119_), .ZN(G651));
  NAND3_X1  g0819(.A1(G161), .A2(G1689), .A3(G1690), .ZN(new_n1121_));
  NAND2_X1  g0820(.A1(G191), .A2(G1690), .ZN(new_n1122_));
  OAI21_X1  g0821(.A(new_n1121_), .B1(new_n1122_), .B2(G1689), .ZN(new_n1123_));
  NOR2_X1   g0822(.A1(G824), .A2(G1690), .ZN(new_n1124_));
  AOI21_X1  g0823(.A(new_n1123_), .B1(new_n1124_), .B2(new_n881_), .ZN(new_n1125_));
  NAND3_X1  g0824(.A1(new_n1054_), .A2(G1689), .A3(new_n875_), .ZN(new_n1126_));
  AOI21_X1  g0825(.A(new_n874_), .B1(new_n1125_), .B2(new_n1126_), .ZN(G654));
  NAND3_X1  g0826(.A1(new_n1078_), .A2(G1691), .A3(new_n884_), .ZN(new_n1128_));
  NAND3_X1  g0827(.A1(G173), .A2(G1691), .A3(G1694), .ZN(new_n1129_));
  NAND2_X1  g0828(.A1(G203), .A2(G1694), .ZN(new_n1130_));
  OAI21_X1  g0829(.A(new_n1129_), .B1(new_n1130_), .B2(G1691), .ZN(new_n1131_));
  NOR2_X1   g0830(.A1(G830), .A2(G1694), .ZN(new_n1132_));
  AOI21_X1  g0831(.A(new_n1131_), .B1(new_n1132_), .B2(new_n890_), .ZN(new_n1133_));
  AOI21_X1  g0832(.A(new_n874_), .B1(new_n1128_), .B2(new_n1133_), .ZN(G679));
  NAND3_X1  g0833(.A1(new_n1071_), .A2(G1691), .A3(new_n884_), .ZN(new_n1135_));
  NAND3_X1  g0834(.A1(G167), .A2(G1691), .A3(G1694), .ZN(new_n1136_));
  NAND2_X1  g0835(.A1(G197), .A2(G1694), .ZN(new_n1137_));
  OAI21_X1  g0836(.A(new_n1136_), .B1(new_n1137_), .B2(G1691), .ZN(new_n1138_));
  NOR2_X1   g0837(.A1(G828), .A2(G1694), .ZN(new_n1139_));
  AOI21_X1  g0838(.A(new_n1138_), .B1(new_n1139_), .B2(new_n890_), .ZN(new_n1140_));
  AOI21_X1  g0839(.A(new_n874_), .B1(new_n1135_), .B2(new_n1140_), .ZN(G682));
  NAND3_X1  g0840(.A1(new_n1064_), .A2(G1691), .A3(new_n884_), .ZN(new_n1142_));
  NAND3_X1  g0841(.A1(G164), .A2(G1691), .A3(G1694), .ZN(new_n1143_));
  NAND2_X1  g0842(.A1(G194), .A2(G1694), .ZN(new_n1144_));
  OAI21_X1  g0843(.A(new_n1143_), .B1(new_n1144_), .B2(G1691), .ZN(new_n1145_));
  NOR2_X1   g0844(.A1(G826), .A2(G1694), .ZN(new_n1146_));
  AOI21_X1  g0845(.A(new_n1145_), .B1(new_n1146_), .B2(new_n890_), .ZN(new_n1147_));
  AOI21_X1  g0846(.A(new_n874_), .B1(new_n1142_), .B2(new_n1147_), .ZN(G685));
  NAND3_X1  g0847(.A1(G161), .A2(G1691), .A3(G1694), .ZN(new_n1149_));
  NAND2_X1  g0848(.A1(G191), .A2(G1694), .ZN(new_n1150_));
  OAI21_X1  g0849(.A(new_n1149_), .B1(new_n1150_), .B2(G1691), .ZN(new_n1151_));
  NOR2_X1   g0850(.A1(G824), .A2(G1694), .ZN(new_n1152_));
  AOI21_X1  g0851(.A(new_n1151_), .B1(new_n1152_), .B2(new_n890_), .ZN(new_n1153_));
  NAND3_X1  g0852(.A1(new_n1054_), .A2(G1691), .A3(new_n884_), .ZN(new_n1154_));
  AOI21_X1  g0853(.A(new_n874_), .B1(new_n1153_), .B2(new_n1154_), .ZN(G688));
  NAND4_X1  g0854(.A1(new_n711_), .A2(new_n710_), .A3(new_n661_), .A4(new_n654_), .ZN(new_n1156_));
  OAI211_X1 g0855(.A(new_n652_), .B(new_n721_), .C1(new_n733_), .C2(new_n573_), .ZN(new_n1157_));
  NAND2_X1  g0856(.A1(new_n1157_), .A2(new_n569_), .ZN(new_n1158_));
  AOI21_X1  g0857(.A(new_n657_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n1159_));
  AOI21_X1  g0858(.A(new_n576_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n1160_));
  AOI21_X1  g0859(.A(new_n653_), .B1(new_n1160_), .B2(new_n559_), .ZN(new_n1161_));
  NAND3_X1  g0860(.A1(new_n1161_), .A2(new_n576_), .A3(new_n721_), .ZN(new_n1162_));
  AND3_X1   g0861(.A1(new_n1158_), .A2(new_n1159_), .A3(new_n1162_), .ZN(new_n1163_));
  AOI21_X1  g0862(.A(new_n1159_), .B1(new_n1158_), .B2(new_n1162_), .ZN(new_n1164_));
  OAI21_X1  g0863(.A(new_n1156_), .B1(new_n1163_), .B2(new_n1164_), .ZN(new_n1165_));
  NOR2_X1   g0864(.A1(new_n1157_), .A2(new_n569_), .ZN(new_n1166_));
  AOI21_X1  g0865(.A(new_n576_), .B1(new_n1161_), .B2(new_n721_), .ZN(new_n1167_));
  OAI22_X1  g0866(.A1(new_n1166_), .A2(new_n1167_), .B1(new_n657_), .B2(new_n1160_), .ZN(new_n1168_));
  INV_X1    g0867(.A(new_n1156_), .ZN(new_n1169_));
  NAND3_X1  g0868(.A1(new_n1158_), .A2(new_n1159_), .A3(new_n1162_), .ZN(new_n1170_));
  NAND3_X1  g0869(.A1(new_n1168_), .A2(new_n1169_), .A3(new_n1170_), .ZN(new_n1171_));
  AND3_X1   g0870(.A1(new_n1165_), .A2(new_n576_), .A3(new_n1171_), .ZN(new_n1172_));
  AOI21_X1  g0871(.A(new_n576_), .B1(new_n1165_), .B2(new_n1171_), .ZN(new_n1173_));
  OAI21_X1  g0872(.A(new_n707_), .B1(new_n1172_), .B2(new_n1173_), .ZN(new_n1174_));
  NOR3_X1   g0873(.A1(new_n1163_), .A2(new_n1164_), .A3(new_n1156_), .ZN(new_n1175_));
  AOI21_X1  g0874(.A(new_n1169_), .B1(new_n1168_), .B2(new_n1170_), .ZN(new_n1176_));
  OAI21_X1  g0875(.A(new_n569_), .B1(new_n1175_), .B2(new_n1176_), .ZN(new_n1177_));
  NAND3_X1  g0876(.A1(new_n1165_), .A2(new_n1171_), .A3(new_n576_), .ZN(new_n1178_));
  NAND3_X1  g0877(.A1(new_n1177_), .A2(new_n565_), .A3(new_n1178_), .ZN(new_n1179_));
  AND3_X1   g0878(.A1(new_n1174_), .A2(new_n549_), .A3(new_n1179_), .ZN(new_n1180_));
  AOI21_X1  g0879(.A(new_n549_), .B1(new_n1174_), .B2(new_n1179_), .ZN(new_n1181_));
  NOR3_X1   g0880(.A1(new_n1180_), .A2(new_n1181_), .A3(new_n573_), .ZN(new_n1182_));
  NOR3_X1   g0881(.A1(new_n1172_), .A2(new_n1173_), .A3(new_n707_), .ZN(new_n1183_));
  AOI21_X1  g0882(.A(new_n565_), .B1(new_n1177_), .B2(new_n1178_), .ZN(new_n1184_));
  OAI21_X1  g0883(.A(new_n548_), .B1(new_n1183_), .B2(new_n1184_), .ZN(new_n1185_));
  NAND3_X1  g0884(.A1(new_n1174_), .A2(new_n549_), .A3(new_n1179_), .ZN(new_n1186_));
  AOI21_X1  g0885(.A(new_n559_), .B1(new_n1185_), .B2(new_n1186_), .ZN(new_n1187_));
  OAI21_X1  g0886(.A(new_n574_), .B1(new_n1182_), .B2(new_n1187_), .ZN(new_n1188_));
  INV_X1    g0887(.A(G2174), .ZN(new_n1189_));
  OAI21_X1  g0888(.A(new_n573_), .B1(new_n1180_), .B2(new_n1181_), .ZN(new_n1190_));
  NAND3_X1  g0889(.A1(new_n1185_), .A2(new_n559_), .A3(new_n1186_), .ZN(new_n1191_));
  NAND3_X1  g0890(.A1(new_n1190_), .A2(new_n553_), .A3(new_n1191_), .ZN(new_n1192_));
  NAND3_X1  g0891(.A1(new_n1188_), .A2(new_n1189_), .A3(new_n1192_), .ZN(new_n1193_));
  NAND2_X1  g0892(.A1(new_n1160_), .A2(new_n559_), .ZN(new_n1194_));
  AOI21_X1  g0893(.A(new_n569_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n1195_));
  NAND2_X1  g0894(.A1(new_n1195_), .A2(new_n559_), .ZN(new_n1196_));
  NAND4_X1  g0895(.A1(new_n1194_), .A2(new_n1196_), .A3(new_n652_), .A4(new_n721_), .ZN(new_n1197_));
  NOR3_X1   g0896(.A1(new_n1160_), .A2(new_n1195_), .A3(new_n657_), .ZN(new_n1198_));
  NAND2_X1  g0897(.A1(new_n1197_), .A2(new_n1198_), .ZN(new_n1199_));
  INV_X1    g0898(.A(new_n1195_), .ZN(new_n1200_));
  NAND2_X1  g0899(.A1(new_n1159_), .A2(new_n1200_), .ZN(new_n1201_));
  OAI21_X1  g0900(.A(new_n559_), .B1(new_n1160_), .B2(new_n1195_), .ZN(new_n1202_));
  NAND4_X1  g0901(.A1(new_n1201_), .A2(new_n1202_), .A3(new_n652_), .A4(new_n721_), .ZN(new_n1203_));
  NAND2_X1  g0902(.A1(new_n1199_), .A2(new_n1203_), .ZN(new_n1204_));
  NAND4_X1  g0903(.A1(new_n559_), .A2(new_n565_), .A3(new_n553_), .A4(new_n576_), .ZN(new_n1205_));
  NAND4_X1  g0904(.A1(new_n711_), .A2(new_n1205_), .A3(new_n661_), .A4(new_n710_), .ZN(new_n1206_));
  NOR2_X1   g0905(.A1(new_n1206_), .A2(new_n655_), .ZN(new_n1207_));
  NAND2_X1  g0906(.A1(new_n1204_), .A2(new_n1207_), .ZN(new_n1208_));
  OAI211_X1 g0907(.A(new_n1199_), .B(new_n1203_), .C1(new_n655_), .C2(new_n1206_), .ZN(new_n1209_));
  NAND3_X1  g0908(.A1(new_n1208_), .A2(new_n576_), .A3(new_n1209_), .ZN(new_n1210_));
  INV_X1    g0909(.A(new_n1210_), .ZN(new_n1211_));
  AOI21_X1  g0910(.A(new_n576_), .B1(new_n1208_), .B2(new_n1209_), .ZN(new_n1212_));
  OAI21_X1  g0911(.A(new_n707_), .B1(new_n1211_), .B2(new_n1212_), .ZN(new_n1213_));
  NAND2_X1  g0912(.A1(new_n1208_), .A2(new_n1209_), .ZN(new_n1214_));
  NAND2_X1  g0913(.A1(new_n1214_), .A2(new_n569_), .ZN(new_n1215_));
  NAND3_X1  g0914(.A1(new_n1215_), .A2(new_n565_), .A3(new_n1210_), .ZN(new_n1216_));
  AND3_X1   g0915(.A1(new_n1213_), .A2(new_n1216_), .A3(new_n549_), .ZN(new_n1217_));
  AOI21_X1  g0916(.A(new_n549_), .B1(new_n1213_), .B2(new_n1216_), .ZN(new_n1218_));
  OAI21_X1  g0917(.A(new_n573_), .B1(new_n1217_), .B2(new_n1218_), .ZN(new_n1219_));
  NAND2_X1  g0918(.A1(new_n1213_), .A2(new_n1216_), .ZN(new_n1220_));
  NAND2_X1  g0919(.A1(new_n1220_), .A2(new_n548_), .ZN(new_n1221_));
  NAND3_X1  g0920(.A1(new_n1213_), .A2(new_n1216_), .A3(new_n549_), .ZN(new_n1222_));
  NAND3_X1  g0921(.A1(new_n1221_), .A2(new_n559_), .A3(new_n1222_), .ZN(new_n1223_));
  AND3_X1   g0922(.A1(new_n1219_), .A2(new_n1223_), .A3(new_n553_), .ZN(new_n1224_));
  AOI21_X1  g0923(.A(new_n553_), .B1(new_n1219_), .B2(new_n1223_), .ZN(new_n1225_));
  OAI21_X1  g0924(.A(G2174), .B1(new_n1224_), .B2(new_n1225_), .ZN(new_n1226_));
  NAND2_X1  g0925(.A1(new_n1193_), .A2(new_n1226_), .ZN(new_n1227_));
  INV_X1    g0926(.A(new_n663_), .ZN(new_n1228_));
  OAI211_X1 g0927(.A(new_n643_), .B(new_n642_), .C1(new_n540_), .C2(new_n542_), .ZN(new_n1229_));
  OAI22_X1  g0928(.A1(G479), .A2(new_n539_), .B1(new_n526_), .B2(G490), .ZN(new_n1230_));
  NAND2_X1  g0929(.A1(new_n1229_), .A2(new_n1230_), .ZN(new_n1231_));
  XNOR2_X1  g0930(.A(new_n694_), .B(new_n1231_), .ZN(new_n1232_));
  NAND2_X1  g0931(.A1(new_n1232_), .A2(new_n528_), .ZN(new_n1233_));
  INV_X1    g0932(.A(new_n1233_), .ZN(new_n1234_));
  NOR2_X1   g0933(.A1(new_n1232_), .A2(new_n528_), .ZN(new_n1235_));
  NOR3_X1   g0934(.A1(new_n1234_), .A2(new_n641_), .A3(new_n1235_), .ZN(new_n1236_));
  OR2_X1    g0935(.A1(new_n1232_), .A2(new_n528_), .ZN(new_n1237_));
  AOI21_X1  g0936(.A(new_n544_), .B1(new_n1237_), .B2(new_n1233_), .ZN(new_n1238_));
  OAI21_X1  g0937(.A(new_n535_), .B1(new_n1236_), .B2(new_n1238_), .ZN(new_n1239_));
  OAI21_X1  g0938(.A(new_n641_), .B1(new_n1234_), .B2(new_n1235_), .ZN(new_n1240_));
  NAND3_X1  g0939(.A1(new_n1237_), .A2(new_n544_), .A3(new_n1233_), .ZN(new_n1241_));
  NAND3_X1  g0940(.A1(new_n1240_), .A2(new_n536_), .A3(new_n1241_), .ZN(new_n1242_));
  AND3_X1   g0941(.A1(new_n1239_), .A2(new_n532_), .A3(new_n1242_), .ZN(new_n1243_));
  AOI21_X1  g0942(.A(new_n532_), .B1(new_n1239_), .B2(new_n1242_), .ZN(new_n1244_));
  OAI211_X1 g0943(.A(new_n1189_), .B(new_n1228_), .C1(new_n1243_), .C2(new_n1244_), .ZN(new_n1245_));
  NAND2_X1  g0944(.A1(new_n663_), .A2(new_n577_), .ZN(new_n1246_));
  OAI211_X1 g0945(.A(G2174), .B(new_n1246_), .C1(new_n1243_), .C2(new_n1244_), .ZN(new_n1247_));
  NAND2_X1  g0946(.A1(new_n864_), .A2(new_n644_), .ZN(new_n1248_));
  AOI211_X1 g0947(.A(new_n531_), .B(new_n648_), .C1(new_n544_), .C2(new_n644_), .ZN(new_n1249_));
  OAI21_X1  g0948(.A(new_n645_), .B1(new_n542_), .B2(new_n540_), .ZN(new_n1250_));
  NAND3_X1  g0949(.A1(new_n1248_), .A2(new_n1249_), .A3(new_n1250_), .ZN(new_n1251_));
  INV_X1    g0950(.A(new_n1251_), .ZN(new_n1252_));
  AOI21_X1  g0951(.A(new_n1249_), .B1(new_n1248_), .B2(new_n1250_), .ZN(new_n1253_));
  NOR3_X1   g0952(.A1(new_n1252_), .A2(new_n527_), .A3(new_n1253_), .ZN(new_n1254_));
  NAND2_X1  g0953(.A1(new_n1248_), .A2(new_n1250_), .ZN(new_n1255_));
  INV_X1    g0954(.A(new_n1249_), .ZN(new_n1256_));
  NAND2_X1  g0955(.A1(new_n1255_), .A2(new_n1256_), .ZN(new_n1257_));
  AOI21_X1  g0956(.A(new_n528_), .B1(new_n1257_), .B2(new_n1251_), .ZN(new_n1258_));
  OAI21_X1  g0957(.A(new_n641_), .B1(new_n1254_), .B2(new_n1258_), .ZN(new_n1259_));
  OAI21_X1  g0958(.A(new_n527_), .B1(new_n1252_), .B2(new_n1253_), .ZN(new_n1260_));
  NAND3_X1  g0959(.A1(new_n1257_), .A2(new_n528_), .A3(new_n1251_), .ZN(new_n1261_));
  NAND3_X1  g0960(.A1(new_n1260_), .A2(new_n544_), .A3(new_n1261_), .ZN(new_n1262_));
  NAND2_X1  g0961(.A1(new_n1259_), .A2(new_n1262_), .ZN(new_n1263_));
  NAND2_X1  g0962(.A1(new_n1263_), .A2(new_n535_), .ZN(new_n1264_));
  NAND3_X1  g0963(.A1(new_n1259_), .A2(new_n536_), .A3(new_n1262_), .ZN(new_n1265_));
  AND3_X1   g0964(.A1(new_n1264_), .A2(new_n532_), .A3(new_n1265_), .ZN(new_n1266_));
  AOI21_X1  g0965(.A(new_n532_), .B1(new_n1264_), .B2(new_n1265_), .ZN(new_n1267_));
  OAI211_X1 g0966(.A(new_n1189_), .B(new_n663_), .C1(new_n1266_), .C2(new_n1267_), .ZN(new_n1268_));
  INV_X1    g0967(.A(new_n1246_), .ZN(new_n1269_));
  OAI211_X1 g0968(.A(G2174), .B(new_n1269_), .C1(new_n1266_), .C2(new_n1267_), .ZN(new_n1270_));
  AND4_X1   g0969(.A1(new_n1245_), .A2(new_n1247_), .A3(new_n1268_), .A4(new_n1270_), .ZN(new_n1271_));
  NAND2_X1  g0970(.A1(new_n1227_), .A2(new_n1271_), .ZN(new_n1272_));
  NAND4_X1  g0971(.A1(new_n1245_), .A2(new_n1247_), .A3(new_n1268_), .A4(new_n1270_), .ZN(new_n1273_));
  NAND3_X1  g0972(.A1(new_n1273_), .A2(new_n1193_), .A3(new_n1226_), .ZN(new_n1274_));
  NAND2_X1  g0973(.A1(new_n1272_), .A2(new_n1274_), .ZN(new_n1275_));
  NAND3_X1  g0974(.A1(new_n1275_), .A2(G4091), .A3(new_n668_), .ZN(new_n1276_));
  AOI21_X1  g0975(.A(G534), .B1(G242), .B2(G351), .ZN(new_n1277_));
  OAI21_X1  g0976(.A(new_n1277_), .B1(new_n364_), .B2(G351), .ZN(new_n1278_));
  NAND3_X1  g0977(.A1(G248), .A2(G351), .A3(G534), .ZN(new_n1279_));
  NAND3_X1  g0978(.A1(new_n390_), .A2(G251), .A3(G534), .ZN(new_n1280_));
  NAND3_X1  g0979(.A1(new_n1278_), .A2(new_n1279_), .A3(new_n1280_), .ZN(new_n1281_));
  AOI21_X1  g0980(.A(G523), .B1(G242), .B2(G341), .ZN(new_n1282_));
  OAI21_X1  g0981(.A(new_n1282_), .B1(new_n364_), .B2(G341), .ZN(new_n1283_));
  NAND3_X1  g0982(.A1(G248), .A2(G341), .A3(G523), .ZN(new_n1284_));
  NAND3_X1  g0983(.A1(new_n382_), .A2(G251), .A3(G523), .ZN(new_n1285_));
  NAND3_X1  g0984(.A1(new_n1283_), .A2(new_n1284_), .A3(new_n1285_), .ZN(new_n1286_));
  XNOR2_X1  g0985(.A(new_n1281_), .B(new_n1286_), .ZN(new_n1287_));
  INV_X1    g0986(.A(new_n1287_), .ZN(new_n1288_));
  AOI21_X1  g0987(.A(G503), .B1(G242), .B2(G324), .ZN(new_n1289_));
  OAI21_X1  g0988(.A(new_n1289_), .B1(new_n364_), .B2(G324), .ZN(new_n1290_));
  NAND3_X1  g0989(.A1(G248), .A2(G324), .A3(G503), .ZN(new_n1291_));
  NAND3_X1  g0990(.A1(new_n397_), .A2(G251), .A3(G503), .ZN(new_n1292_));
  NAND3_X1  g0991(.A1(new_n1290_), .A2(new_n1291_), .A3(new_n1292_), .ZN(new_n1293_));
  NOR2_X1   g0992(.A1(G242), .A2(G514), .ZN(new_n1294_));
  AOI21_X1  g0993(.A(new_n1294_), .B1(G248), .B2(G514), .ZN(new_n1295_));
  XNOR2_X1  g0994(.A(new_n1293_), .B(new_n1295_), .ZN(new_n1296_));
  OR3_X1    g0995(.A1(new_n1288_), .A2(new_n409_), .A3(new_n1296_), .ZN(new_n1297_));
  OR3_X1    g0996(.A1(new_n1287_), .A2(new_n1296_), .A3(new_n408_), .ZN(new_n1298_));
  NAND3_X1  g0997(.A1(new_n1287_), .A2(new_n1296_), .A3(new_n409_), .ZN(new_n1299_));
  NAND3_X1  g0998(.A1(new_n1288_), .A2(new_n408_), .A3(new_n1296_), .ZN(new_n1300_));
  NAND4_X1  g0999(.A1(new_n1297_), .A2(new_n1298_), .A3(new_n1299_), .A4(new_n1300_), .ZN(new_n1301_));
  XNOR2_X1  g1000(.A(new_n372_), .B(new_n378_), .ZN(new_n1302_));
  XNOR2_X1  g1001(.A(new_n362_), .B(new_n365_), .ZN(new_n1303_));
  XNOR2_X1  g1002(.A(new_n1302_), .B(new_n1303_), .ZN(new_n1304_));
  XNOR2_X1  g1003(.A(new_n1301_), .B(new_n1304_), .ZN(new_n1305_));
  OR3_X1    g1004(.A1(new_n1305_), .A2(G4091), .A3(G4092), .ZN(new_n1306_));
  OAI21_X1  g1005(.A(G4092), .B1(G120), .B2(G4091), .ZN(new_n1307_));
  NAND3_X1  g1006(.A1(new_n1276_), .A2(new_n1306_), .A3(new_n1307_), .ZN(G843));
  INV_X1    g1007(.A(G1497), .ZN(new_n1309_));
  INV_X1    g1008(.A(new_n639_), .ZN(new_n1310_));
  OAI211_X1 g1009(.A(new_n618_), .B(new_n421_), .C1(new_n513_), .C2(new_n414_), .ZN(new_n1311_));
  OAI22_X1  g1010(.A1(G422), .A2(new_n504_), .B1(new_n515_), .B2(G468), .ZN(new_n1312_));
  NAND2_X1  g1011(.A1(new_n1311_), .A2(new_n1312_), .ZN(new_n1313_));
  XNOR2_X1  g1012(.A(new_n838_), .B(new_n1313_), .ZN(new_n1314_));
  NAND2_X1  g1013(.A1(new_n1314_), .A2(new_n506_), .ZN(new_n1315_));
  INV_X1    g1014(.A(new_n1315_), .ZN(new_n1316_));
  NOR2_X1   g1015(.A1(new_n1314_), .A2(new_n506_), .ZN(new_n1317_));
  NOR3_X1   g1016(.A1(new_n1316_), .A2(new_n848_), .A3(new_n1317_), .ZN(new_n1318_));
  OR2_X1    g1017(.A1(new_n1314_), .A2(new_n506_), .ZN(new_n1319_));
  AOI21_X1  g1018(.A(new_n517_), .B1(new_n1319_), .B2(new_n1315_), .ZN(new_n1320_));
  OAI21_X1  g1019(.A(new_n509_), .B1(new_n1318_), .B2(new_n1320_), .ZN(new_n1321_));
  OAI21_X1  g1020(.A(new_n848_), .B1(new_n1316_), .B2(new_n1317_), .ZN(new_n1322_));
  NAND3_X1  g1021(.A1(new_n1319_), .A2(new_n517_), .A3(new_n1315_), .ZN(new_n1323_));
  NAND3_X1  g1022(.A1(new_n1322_), .A2(new_n510_), .A3(new_n1323_), .ZN(new_n1324_));
  AND3_X1   g1023(.A1(new_n1321_), .A2(new_n520_), .A3(new_n1324_), .ZN(new_n1325_));
  AOI21_X1  g1024(.A(new_n520_), .B1(new_n1321_), .B2(new_n1324_), .ZN(new_n1326_));
  OAI211_X1 g1025(.A(new_n1309_), .B(new_n1310_), .C1(new_n1325_), .C2(new_n1326_), .ZN(new_n1327_));
  OAI21_X1  g1026(.A(new_n619_), .B1(G468), .B2(new_n515_), .ZN(new_n1328_));
  INV_X1    g1027(.A(new_n1328_), .ZN(new_n1329_));
  AOI21_X1  g1028(.A(new_n619_), .B1(G468), .B2(new_n515_), .ZN(new_n1330_));
  NOR2_X1   g1029(.A1(new_n1329_), .A2(new_n1330_), .ZN(new_n1331_));
  NAND3_X1  g1030(.A1(new_n517_), .A2(new_n520_), .A3(new_n619_), .ZN(new_n1332_));
  NAND3_X1  g1031(.A1(new_n1332_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n1333_));
  XNOR2_X1  g1032(.A(new_n1331_), .B(new_n1333_), .ZN(new_n1334_));
  OR2_X1    g1033(.A1(new_n1334_), .A2(new_n506_), .ZN(new_n1335_));
  NAND2_X1  g1034(.A1(new_n1334_), .A2(new_n506_), .ZN(new_n1336_));
  NAND3_X1  g1035(.A1(new_n1335_), .A2(new_n517_), .A3(new_n1336_), .ZN(new_n1337_));
  INV_X1    g1036(.A(new_n1337_), .ZN(new_n1338_));
  AOI21_X1  g1037(.A(new_n517_), .B1(new_n1335_), .B2(new_n1336_), .ZN(new_n1339_));
  OAI21_X1  g1038(.A(new_n509_), .B1(new_n1338_), .B2(new_n1339_), .ZN(new_n1340_));
  XNOR2_X1  g1039(.A(new_n1334_), .B(new_n506_), .ZN(new_n1341_));
  NAND2_X1  g1040(.A1(new_n1341_), .A2(new_n848_), .ZN(new_n1342_));
  NAND3_X1  g1041(.A1(new_n1342_), .A2(new_n510_), .A3(new_n1337_), .ZN(new_n1343_));
  AND3_X1   g1042(.A1(new_n1340_), .A2(new_n520_), .A3(new_n1343_), .ZN(new_n1344_));
  AOI21_X1  g1043(.A(new_n520_), .B1(new_n1340_), .B2(new_n1343_), .ZN(new_n1345_));
  OAI211_X1 g1044(.A(new_n1309_), .B(new_n639_), .C1(new_n1344_), .C2(new_n1345_), .ZN(new_n1346_));
  NAND2_X1  g1045(.A1(new_n639_), .A2(new_n501_), .ZN(new_n1347_));
  INV_X1    g1046(.A(new_n1347_), .ZN(new_n1348_));
  OAI211_X1 g1047(.A(G1497), .B(new_n1348_), .C1(new_n1344_), .C2(new_n1345_), .ZN(new_n1349_));
  OAI211_X1 g1048(.A(G1497), .B(new_n1347_), .C1(new_n1325_), .C2(new_n1326_), .ZN(new_n1350_));
  AND4_X1   g1049(.A1(new_n1327_), .A2(new_n1346_), .A3(new_n1349_), .A4(new_n1350_), .ZN(new_n1351_));
  NAND4_X1  g1050(.A1(new_n500_), .A2(new_n479_), .A3(new_n496_), .A4(new_n584_), .ZN(new_n1352_));
  NAND4_X1  g1051(.A1(new_n1352_), .A2(new_n749_), .A3(new_n637_), .A4(new_n748_), .ZN(new_n1353_));
  NOR2_X1   g1052(.A1(new_n1353_), .A2(new_n631_), .ZN(new_n1354_));
  OAI211_X1 g1053(.A(new_n496_), .B(new_n584_), .C1(G374), .C2(new_n499_), .ZN(new_n1355_));
  NAND3_X1  g1054(.A1(new_n1355_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n1356_));
  INV_X1    g1055(.A(new_n499_), .ZN(new_n1357_));
  NAND2_X1  g1056(.A1(new_n1357_), .A2(new_n443_), .ZN(new_n1358_));
  NAND2_X1  g1057(.A1(new_n1356_), .A2(new_n1358_), .ZN(new_n1359_));
  NAND2_X1  g1058(.A1(new_n776_), .A2(new_n773_), .ZN(new_n1360_));
  INV_X1    g1059(.A(new_n1360_), .ZN(new_n1361_));
  OAI21_X1  g1060(.A(new_n1361_), .B1(new_n785_), .B2(new_n586_), .ZN(new_n1362_));
  INV_X1    g1061(.A(new_n1358_), .ZN(new_n1363_));
  NAND4_X1  g1062(.A1(new_n1355_), .A2(new_n761_), .A3(new_n762_), .A4(new_n1363_), .ZN(new_n1364_));
  AND3_X1   g1063(.A1(new_n1359_), .A2(new_n1362_), .A3(new_n1364_), .ZN(new_n1365_));
  AOI21_X1  g1064(.A(new_n1362_), .B1(new_n1359_), .B2(new_n1364_), .ZN(new_n1366_));
  OAI21_X1  g1065(.A(new_n1354_), .B1(new_n1365_), .B2(new_n1366_), .ZN(new_n1367_));
  NAND2_X1  g1066(.A1(new_n1359_), .A2(new_n1364_), .ZN(new_n1368_));
  INV_X1    g1067(.A(new_n1362_), .ZN(new_n1369_));
  NAND2_X1  g1068(.A1(new_n1368_), .A2(new_n1369_), .ZN(new_n1370_));
  OR2_X1    g1069(.A1(new_n1353_), .A2(new_n631_), .ZN(new_n1371_));
  NAND3_X1  g1070(.A1(new_n1359_), .A2(new_n1362_), .A3(new_n1364_), .ZN(new_n1372_));
  NAND3_X1  g1071(.A1(new_n1370_), .A2(new_n1371_), .A3(new_n1372_), .ZN(new_n1373_));
  AND3_X1   g1072(.A1(new_n1367_), .A2(new_n1373_), .A3(new_n500_), .ZN(new_n1374_));
  AOI21_X1  g1073(.A(new_n500_), .B1(new_n1367_), .B2(new_n1373_), .ZN(new_n1375_));
  OAI21_X1  g1074(.A(new_n785_), .B1(new_n1374_), .B2(new_n1375_), .ZN(new_n1376_));
  NOR3_X1   g1075(.A1(new_n1365_), .A2(new_n1366_), .A3(new_n1354_), .ZN(new_n1377_));
  AOI21_X1  g1076(.A(new_n1371_), .B1(new_n1370_), .B2(new_n1372_), .ZN(new_n1378_));
  OAI21_X1  g1077(.A(new_n586_), .B1(new_n1377_), .B2(new_n1378_), .ZN(new_n1379_));
  NAND3_X1  g1078(.A1(new_n1367_), .A2(new_n1373_), .A3(new_n500_), .ZN(new_n1380_));
  NAND3_X1  g1079(.A1(new_n1379_), .A2(new_n496_), .A3(new_n1380_), .ZN(new_n1381_));
  AND3_X1   g1080(.A1(new_n1376_), .A2(new_n581_), .A3(new_n1381_), .ZN(new_n1382_));
  AOI21_X1  g1081(.A(new_n581_), .B1(new_n1376_), .B2(new_n1381_), .ZN(new_n1383_));
  NOR3_X1   g1082(.A1(new_n1382_), .A2(new_n1383_), .A3(new_n487_), .ZN(new_n1384_));
  NOR3_X1   g1083(.A1(new_n1374_), .A2(new_n1375_), .A3(new_n785_), .ZN(new_n1385_));
  AOI21_X1  g1084(.A(new_n496_), .B1(new_n1379_), .B2(new_n1380_), .ZN(new_n1386_));
  OAI21_X1  g1085(.A(new_n490_), .B1(new_n1385_), .B2(new_n1386_), .ZN(new_n1387_));
  NAND3_X1  g1086(.A1(new_n1376_), .A2(new_n1381_), .A3(new_n581_), .ZN(new_n1388_));
  AOI21_X1  g1087(.A(new_n584_), .B1(new_n1387_), .B2(new_n1388_), .ZN(new_n1389_));
  OAI21_X1  g1088(.A(new_n480_), .B1(new_n1384_), .B2(new_n1389_), .ZN(new_n1390_));
  OAI21_X1  g1089(.A(new_n487_), .B1(new_n1382_), .B2(new_n1383_), .ZN(new_n1391_));
  NAND3_X1  g1090(.A1(new_n1387_), .A2(new_n584_), .A3(new_n1388_), .ZN(new_n1392_));
  NAND3_X1  g1091(.A1(new_n1391_), .A2(new_n479_), .A3(new_n1392_), .ZN(new_n1393_));
  AOI21_X1  g1092(.A(new_n1309_), .B1(new_n1390_), .B2(new_n1393_), .ZN(new_n1394_));
  NAND4_X1  g1093(.A1(new_n749_), .A2(new_n630_), .A3(new_n748_), .A4(new_n637_), .ZN(new_n1395_));
  OAI211_X1 g1094(.A(new_n761_), .B(new_n762_), .C1(new_n776_), .C2(new_n487_), .ZN(new_n1396_));
  NAND2_X1  g1095(.A1(new_n1396_), .A2(new_n625_), .ZN(new_n1397_));
  NAND4_X1  g1096(.A1(new_n763_), .A2(new_n761_), .A3(new_n626_), .A4(new_n762_), .ZN(new_n1398_));
  AND3_X1   g1097(.A1(new_n1397_), .A2(new_n1361_), .A3(new_n1398_), .ZN(new_n1399_));
  AOI21_X1  g1098(.A(new_n1361_), .B1(new_n1397_), .B2(new_n1398_), .ZN(new_n1400_));
  OAI21_X1  g1099(.A(new_n1395_), .B1(new_n1399_), .B2(new_n1400_), .ZN(new_n1401_));
  NAND2_X1  g1100(.A1(new_n1397_), .A2(new_n1398_), .ZN(new_n1402_));
  NAND2_X1  g1101(.A1(new_n1402_), .A2(new_n1360_), .ZN(new_n1403_));
  INV_X1    g1102(.A(new_n1395_), .ZN(new_n1404_));
  NAND3_X1  g1103(.A1(new_n1397_), .A2(new_n1361_), .A3(new_n1398_), .ZN(new_n1405_));
  NAND3_X1  g1104(.A1(new_n1403_), .A2(new_n1404_), .A3(new_n1405_), .ZN(new_n1406_));
  AND3_X1   g1105(.A1(new_n1401_), .A2(new_n1406_), .A3(new_n500_), .ZN(new_n1407_));
  AOI21_X1  g1106(.A(new_n500_), .B1(new_n1401_), .B2(new_n1406_), .ZN(new_n1408_));
  OAI21_X1  g1107(.A(new_n785_), .B1(new_n1407_), .B2(new_n1408_), .ZN(new_n1409_));
  NOR3_X1   g1108(.A1(new_n1399_), .A2(new_n1400_), .A3(new_n1395_), .ZN(new_n1410_));
  AOI21_X1  g1109(.A(new_n1404_), .B1(new_n1403_), .B2(new_n1405_), .ZN(new_n1411_));
  OAI21_X1  g1110(.A(new_n586_), .B1(new_n1410_), .B2(new_n1411_), .ZN(new_n1412_));
  NAND3_X1  g1111(.A1(new_n1401_), .A2(new_n1406_), .A3(new_n500_), .ZN(new_n1413_));
  NAND3_X1  g1112(.A1(new_n1412_), .A2(new_n496_), .A3(new_n1413_), .ZN(new_n1414_));
  AND3_X1   g1113(.A1(new_n1409_), .A2(new_n581_), .A3(new_n1414_), .ZN(new_n1415_));
  AOI21_X1  g1114(.A(new_n581_), .B1(new_n1409_), .B2(new_n1414_), .ZN(new_n1416_));
  OAI21_X1  g1115(.A(new_n487_), .B1(new_n1415_), .B2(new_n1416_), .ZN(new_n1417_));
  NOR3_X1   g1116(.A1(new_n1407_), .A2(new_n1408_), .A3(new_n785_), .ZN(new_n1418_));
  AOI21_X1  g1117(.A(new_n496_), .B1(new_n1412_), .B2(new_n1413_), .ZN(new_n1419_));
  OAI21_X1  g1118(.A(new_n490_), .B1(new_n1418_), .B2(new_n1419_), .ZN(new_n1420_));
  NAND3_X1  g1119(.A1(new_n1409_), .A2(new_n1414_), .A3(new_n581_), .ZN(new_n1421_));
  NAND3_X1  g1120(.A1(new_n1420_), .A2(new_n584_), .A3(new_n1421_), .ZN(new_n1422_));
  AND3_X1   g1121(.A1(new_n1417_), .A2(new_n479_), .A3(new_n1422_), .ZN(new_n1423_));
  AOI21_X1  g1122(.A(new_n479_), .B1(new_n1417_), .B2(new_n1422_), .ZN(new_n1424_));
  NOR3_X1   g1123(.A1(new_n1423_), .A2(new_n1424_), .A3(G1497), .ZN(new_n1425_));
  OAI21_X1  g1124(.A(new_n1351_), .B1(new_n1394_), .B2(new_n1425_), .ZN(new_n1426_));
  AND3_X1   g1125(.A1(new_n1391_), .A2(new_n479_), .A3(new_n1392_), .ZN(new_n1427_));
  AOI21_X1  g1126(.A(new_n479_), .B1(new_n1391_), .B2(new_n1392_), .ZN(new_n1428_));
  OAI21_X1  g1127(.A(G1497), .B1(new_n1427_), .B2(new_n1428_), .ZN(new_n1429_));
  INV_X1    g1128(.A(new_n1424_), .ZN(new_n1430_));
  NAND3_X1  g1129(.A1(new_n1417_), .A2(new_n479_), .A3(new_n1422_), .ZN(new_n1431_));
  NAND3_X1  g1130(.A1(new_n1430_), .A2(new_n1309_), .A3(new_n1431_), .ZN(new_n1432_));
  NAND4_X1  g1131(.A1(new_n1346_), .A2(new_n1349_), .A3(new_n1327_), .A4(new_n1350_), .ZN(new_n1433_));
  NAND3_X1  g1132(.A1(new_n1429_), .A2(new_n1432_), .A3(new_n1433_), .ZN(new_n1434_));
  NAND2_X1  g1133(.A1(new_n1426_), .A2(new_n1434_), .ZN(new_n1435_));
  NAND3_X1  g1134(.A1(new_n1435_), .A2(G4091), .A3(new_n668_), .ZN(new_n1436_));
  AOI21_X1  g1135(.A(G389), .B1(G242), .B2(G257), .ZN(new_n1437_));
  OAI21_X1  g1136(.A(new_n1437_), .B1(new_n364_), .B2(G257), .ZN(new_n1438_));
  NAND3_X1  g1137(.A1(G248), .A2(G257), .A3(G389), .ZN(new_n1439_));
  NAND3_X1  g1138(.A1(new_n455_), .A2(G251), .A3(G389), .ZN(new_n1440_));
  NAND3_X1  g1139(.A1(new_n1438_), .A2(new_n1439_), .A3(new_n1440_), .ZN(new_n1441_));
  AOI21_X1  g1140(.A(G435), .B1(G234), .B2(G242), .ZN(new_n1442_));
  OAI21_X1  g1141(.A(new_n1442_), .B1(G234), .B2(new_n364_), .ZN(new_n1443_));
  NAND3_X1  g1142(.A1(G234), .A2(G248), .A3(G435), .ZN(new_n1444_));
  NAND3_X1  g1143(.A1(new_n426_), .A2(G251), .A3(G435), .ZN(new_n1445_));
  NAND3_X1  g1144(.A1(new_n1443_), .A2(new_n1444_), .A3(new_n1445_), .ZN(new_n1446_));
  XOR2_X1   g1145(.A(new_n1441_), .B(new_n1446_), .Z(new_n1447_));
  AOI21_X1  g1146(.A(G411), .B1(G242), .B2(G273), .ZN(new_n1448_));
  OAI21_X1  g1147(.A(new_n1448_), .B1(new_n364_), .B2(G273), .ZN(new_n1449_));
  NAND3_X1  g1148(.A1(G248), .A2(G273), .A3(G411), .ZN(new_n1450_));
  NAND3_X1  g1149(.A1(new_n448_), .A2(G251), .A3(G411), .ZN(new_n1451_));
  NAND3_X1  g1150(.A1(new_n1449_), .A2(new_n1450_), .A3(new_n1451_), .ZN(new_n1452_));
  AOI21_X1  g1151(.A(G400), .B1(G242), .B2(G265), .ZN(new_n1453_));
  OAI21_X1  g1152(.A(new_n1453_), .B1(new_n364_), .B2(G265), .ZN(new_n1454_));
  NAND3_X1  g1153(.A1(G248), .A2(G265), .A3(G400), .ZN(new_n1455_));
  NAND3_X1  g1154(.A1(new_n462_), .A2(G251), .A3(G400), .ZN(new_n1456_));
  NAND3_X1  g1155(.A1(new_n1454_), .A2(new_n1455_), .A3(new_n1456_), .ZN(new_n1457_));
  XNOR2_X1  g1156(.A(new_n1452_), .B(new_n1457_), .ZN(new_n1458_));
  AOI21_X1  g1157(.A(G374), .B1(G242), .B2(G281), .ZN(new_n1459_));
  OAI21_X1  g1158(.A(new_n1459_), .B1(new_n364_), .B2(G281), .ZN(new_n1460_));
  NAND3_X1  g1159(.A1(G248), .A2(G281), .A3(G374), .ZN(new_n1461_));
  NAND3_X1  g1160(.A1(new_n441_), .A2(G251), .A3(G374), .ZN(new_n1462_));
  NAND3_X1  g1161(.A1(new_n1460_), .A2(new_n1461_), .A3(new_n1462_), .ZN(new_n1463_));
  NOR3_X1   g1162(.A1(new_n1447_), .A2(new_n1458_), .A3(new_n1463_), .ZN(new_n1464_));
  INV_X1    g1163(.A(new_n1458_), .ZN(new_n1465_));
  AND2_X1   g1164(.A1(new_n1465_), .A2(new_n1447_), .ZN(new_n1466_));
  AOI21_X1  g1165(.A(new_n1464_), .B1(new_n1466_), .B2(new_n1463_), .ZN(new_n1467_));
  INV_X1    g1166(.A(new_n1463_), .ZN(new_n1468_));
  OR3_X1    g1167(.A1(new_n1465_), .A2(new_n1447_), .A3(new_n1468_), .ZN(new_n1469_));
  NAND3_X1  g1168(.A1(new_n1447_), .A2(new_n1458_), .A3(new_n1468_), .ZN(new_n1470_));
  NAND3_X1  g1169(.A1(new_n1467_), .A2(new_n1469_), .A3(new_n1470_), .ZN(new_n1471_));
  AOI21_X1  g1170(.A(G468), .B1(G218), .B2(G242), .ZN(new_n1472_));
  OAI21_X1  g1171(.A(new_n1472_), .B1(G218), .B2(new_n364_), .ZN(new_n1473_));
  NAND3_X1  g1172(.A1(G218), .A2(G248), .A3(G468), .ZN(new_n1474_));
  OAI211_X1 g1173(.A(new_n1473_), .B(new_n1474_), .C1(new_n360_), .C2(new_n413_), .ZN(new_n1475_));
  AOI21_X1  g1174(.A(G422), .B1(G226), .B2(G242), .ZN(new_n1476_));
  OAI21_X1  g1175(.A(new_n1476_), .B1(G226), .B2(new_n364_), .ZN(new_n1477_));
  NAND3_X1  g1176(.A1(G226), .A2(G248), .A3(G422), .ZN(new_n1478_));
  NAND3_X1  g1177(.A1(new_n419_), .A2(G251), .A3(G422), .ZN(new_n1479_));
  NAND3_X1  g1178(.A1(new_n1477_), .A2(new_n1478_), .A3(new_n1479_), .ZN(new_n1480_));
  XNOR2_X1  g1179(.A(new_n1475_), .B(new_n1480_), .ZN(new_n1481_));
  AOI21_X1  g1180(.A(G457), .B1(G210), .B2(G242), .ZN(new_n1482_));
  OAI21_X1  g1181(.A(new_n1482_), .B1(G210), .B2(new_n364_), .ZN(new_n1483_));
  NAND3_X1  g1182(.A1(G210), .A2(G248), .A3(G457), .ZN(new_n1484_));
  NAND3_X1  g1183(.A1(new_n433_), .A2(G251), .A3(G457), .ZN(new_n1485_));
  NAND3_X1  g1184(.A1(new_n1483_), .A2(new_n1484_), .A3(new_n1485_), .ZN(new_n1486_));
  XNOR2_X1  g1185(.A(new_n474_), .B(new_n1486_), .ZN(new_n1487_));
  XNOR2_X1  g1186(.A(new_n1481_), .B(new_n1487_), .ZN(new_n1488_));
  XOR2_X1   g1187(.A(new_n1471_), .B(new_n1488_), .Z(new_n1489_));
  NAND3_X1  g1188(.A1(new_n1489_), .A2(new_n670_), .A3(new_n668_), .ZN(new_n1490_));
  OAI21_X1  g1189(.A(G4092), .B1(G118), .B2(G4091), .ZN(new_n1491_));
  NAND3_X1  g1190(.A1(new_n1436_), .A2(new_n1490_), .A3(new_n1491_), .ZN(G882));
  NAND3_X1  g1191(.A1(new_n1426_), .A2(new_n1434_), .A3(G4091), .ZN(new_n1493_));
  OR2_X1    g1192(.A1(new_n1489_), .A2(G4091), .ZN(new_n1494_));
  AOI21_X1  g1193(.A(G4092), .B1(new_n1493_), .B2(new_n1494_), .ZN(new_n1495_));
  AND2_X1   g1194(.A1(G97), .A2(G4092), .ZN(new_n1496_));
  OAI211_X1 g1195(.A(new_n700_), .B(G4088), .C1(new_n1495_), .C2(new_n1496_), .ZN(new_n1497_));
  NAND3_X1  g1196(.A1(new_n1272_), .A2(G4091), .A3(new_n1274_), .ZN(new_n1498_));
  NAND2_X1  g1197(.A1(new_n1305_), .A2(new_n670_), .ZN(new_n1499_));
  AOI21_X1  g1198(.A(G4092), .B1(new_n1498_), .B2(new_n1499_), .ZN(new_n1500_));
  AND2_X1   g1199(.A1(G94), .A2(G4092), .ZN(new_n1501_));
  OAI211_X1 g1200(.A(new_n700_), .B(new_n704_), .C1(new_n1500_), .C2(new_n1501_), .ZN(new_n1502_));
  NAND3_X1  g1201(.A1(G64), .A2(G4087), .A3(G4088), .ZN(new_n1503_));
  NAND3_X1  g1202(.A1(new_n704_), .A2(G14), .A3(G4087), .ZN(new_n1504_));
  NAND4_X1  g1203(.A1(new_n1497_), .A2(new_n1502_), .A3(new_n1503_), .A4(new_n1504_), .ZN(G767));
  OAI211_X1 g1204(.A(G4089), .B(new_n741_), .C1(new_n1495_), .C2(new_n1496_), .ZN(new_n1506_));
  OAI211_X1 g1205(.A(new_n745_), .B(new_n741_), .C1(new_n1500_), .C2(new_n1501_), .ZN(new_n1507_));
  NAND3_X1  g1206(.A1(G64), .A2(G4089), .A3(G4090), .ZN(new_n1508_));
  NAND3_X1  g1207(.A1(new_n745_), .A2(G14), .A3(G4090), .ZN(new_n1509_));
  NAND4_X1  g1208(.A1(new_n1506_), .A2(new_n1507_), .A3(new_n1508_), .A4(new_n1509_), .ZN(G807));
  OAI211_X1 g1209(.A(G1689), .B(new_n875_), .C1(new_n1495_), .C2(new_n1496_), .ZN(new_n1511_));
  OAI211_X1 g1210(.A(new_n881_), .B(new_n875_), .C1(new_n1500_), .C2(new_n1501_), .ZN(new_n1512_));
  NAND3_X1  g1211(.A1(new_n881_), .A2(G176), .A3(G1690), .ZN(new_n1513_));
  NAND3_X1  g1212(.A1(G179), .A2(G1689), .A3(G1690), .ZN(new_n1514_));
  AND2_X1   g1213(.A1(new_n1513_), .A2(new_n1514_), .ZN(new_n1515_));
  NAND3_X1  g1214(.A1(new_n1511_), .A2(new_n1512_), .A3(new_n1515_), .ZN(new_n1516_));
  NAND2_X1  g1215(.A1(new_n1516_), .A2(G137), .ZN(G658));
  OAI211_X1 g1216(.A(G1691), .B(new_n884_), .C1(new_n1495_), .C2(new_n1496_), .ZN(new_n1518_));
  OAI211_X1 g1217(.A(new_n890_), .B(new_n884_), .C1(new_n1500_), .C2(new_n1501_), .ZN(new_n1519_));
  NAND3_X1  g1218(.A1(new_n890_), .A2(G176), .A3(G1694), .ZN(new_n1520_));
  NAND3_X1  g1219(.A1(G179), .A2(G1691), .A3(G1694), .ZN(new_n1521_));
  AND2_X1   g1220(.A1(new_n1520_), .A2(new_n1521_), .ZN(new_n1522_));
  NAND3_X1  g1221(.A1(new_n1518_), .A2(new_n1519_), .A3(new_n1522_), .ZN(new_n1523_));
  NAND2_X1  g1222(.A1(new_n1523_), .A2(G137), .ZN(G690));
endmodule


