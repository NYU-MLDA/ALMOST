//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_;
  INV_X1    g000(.A(KEYINPUT104), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT23), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G183gat), .A3(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n204_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT22), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(KEYINPUT22), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n214_), .B(new_n217_), .C1(new_n218_), .C2(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n203_), .A2(KEYINPUT24), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n223_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n209_), .A2(KEYINPUT82), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n232_), .A2(new_n208_), .A3(G183gat), .A4(G190gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n230_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n220_), .B1(new_n229_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT30), .ZN(new_n236_));
  INV_X1    g035(.A(G99gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT31), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n236_), .B(G99gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT31), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(KEYINPUT84), .B(KEYINPUT85), .Z(new_n243_));
  XNOR2_X1  g042(.A(G15gat), .B(G43gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G71gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n245_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT86), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n249_), .B(new_n250_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n254_), .B2(new_n252_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n248_), .B(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n239_), .A2(new_n242_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G8gat), .B(G36gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n262_), .B(new_n263_), .Z(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT22), .B(G169gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n204_), .B1(new_n265_), .B2(new_n214_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n234_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT98), .A3(new_n212_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT98), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n234_), .B2(new_n211_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n267_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n225_), .B1(new_n224_), .B2(KEYINPUT96), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(KEYINPUT96), .B2(new_n224_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n223_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n210_), .A2(new_n228_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(KEYINPUT97), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(KEYINPUT97), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n275_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n272_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G197gat), .B(G204gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT21), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n282_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n286_), .A3(new_n284_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n280_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT20), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n285_), .A2(new_n287_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n293_), .B1(new_n235_), .B2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(new_n292_), .A3(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n294_), .B1(new_n272_), .B2(new_n279_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n229_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n298_), .A2(new_n268_), .B1(new_n219_), .B2(new_n213_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n293_), .B1(new_n288_), .B2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n292_), .B1(new_n297_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT99), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n296_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n301_), .A2(new_n302_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n264_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n297_), .A2(new_n300_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT99), .B1(new_n306_), .B2(new_n292_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n302_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n264_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .A4(new_n296_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT4), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT87), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT87), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(G141gat), .A3(G148gat), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n314_), .B(new_n316_), .C1(G141gat), .C2(G148gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT1), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n318_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT1), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n317_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n314_), .A2(new_n316_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G141gat), .ZN(new_n329_));
  INV_X1    g128(.A(G148gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(KEYINPUT3), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n332_), .B1(G141gat), .B2(G148gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n328_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT89), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(KEYINPUT89), .A3(new_n328_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n323_), .A2(new_n322_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n326_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n254_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n340_), .A2(KEYINPUT89), .A3(new_n328_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT89), .B1(new_n340_), .B2(new_n328_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n343_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n326_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n255_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n312_), .B1(new_n345_), .B2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT4), .B1(new_n350_), .B2(new_n255_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n345_), .B2(new_n351_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G1gat), .B(G29gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n360_), .A2(KEYINPUT33), .A3(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n355_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT102), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n345_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n370_), .A2(new_n365_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n368_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT33), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n358_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n365_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n311_), .A2(new_n367_), .A3(new_n374_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n360_), .A2(new_n366_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n365_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n309_), .A2(KEYINPUT32), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n307_), .A2(new_n308_), .A3(new_n296_), .A4(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n289_), .A2(new_n295_), .ZN(new_n384_));
  MUX2_X1   g183(.A(new_n384_), .B(new_n306_), .S(new_n292_), .Z(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(KEYINPUT32), .A3(new_n309_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n381_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n259_), .B1(new_n378_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT91), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G228gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n393_), .A2(new_n395_), .A3(new_n288_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n343_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT29), .B1(new_n398_), .B2(new_n326_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n394_), .B1(new_n399_), .B2(new_n294_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n391_), .B1(new_n396_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n395_), .B1(new_n393_), .B2(new_n288_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n394_), .A3(new_n294_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n390_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT28), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n344_), .B2(new_n392_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n348_), .A2(new_n349_), .A3(new_n406_), .A4(new_n392_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT90), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G22gat), .B(G50gat), .Z(new_n411_));
  NAND3_X1  g210(.A1(new_n348_), .A2(new_n349_), .A3(new_n392_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT28), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n408_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n410_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n411_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n413_), .A2(new_n414_), .A3(new_n408_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n414_), .B1(new_n413_), .B2(new_n408_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n405_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n404_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n401_), .A2(KEYINPUT92), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n402_), .A2(new_n403_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT92), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n391_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n420_), .A2(new_n416_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n428_), .A2(KEYINPUT93), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT93), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n426_), .B1(new_n425_), .B2(new_n391_), .ZN(new_n432_));
  AOI211_X1 g231(.A(KEYINPUT92), .B(new_n390_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n404_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n418_), .A2(new_n419_), .A3(new_n417_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n411_), .B1(new_n410_), .B2(new_n415_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n431_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n422_), .B1(new_n430_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT94), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT93), .B1(new_n428_), .B2(new_n429_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n434_), .A2(new_n437_), .A3(new_n431_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(KEYINPUT94), .A3(new_n422_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n388_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n259_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT94), .B1(new_n444_), .B2(new_n422_), .ZN(new_n448_));
  AOI211_X1 g247(.A(new_n440_), .B(new_n421_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n441_), .A2(new_n445_), .A3(new_n259_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n311_), .A2(KEYINPUT27), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n385_), .A2(KEYINPUT103), .A3(new_n264_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT103), .B1(new_n385_), .B2(new_n264_), .ZN(new_n455_));
  OAI211_X1 g254(.A(KEYINPUT27), .B(new_n310_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n381_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n446_), .B1(new_n452_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G229gat), .A2(G233gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT78), .B(G15gat), .ZN(new_n463_));
  INV_X1    g262(.A(G22gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT79), .B(G1gat), .ZN(new_n466_));
  INV_X1    g265(.A(G8gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT14), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G1gat), .B(G8gat), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n465_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n469_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G29gat), .B(G36gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT81), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n465_), .A2(new_n468_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n469_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n465_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n478_), .B1(new_n483_), .B2(new_n475_), .ZN(new_n484_));
  AOI211_X1 g283(.A(KEYINPUT81), .B(new_n476_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n462_), .B(new_n477_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT81), .B1(new_n472_), .B2(new_n476_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n478_), .A3(new_n475_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n475_), .B(new_n490_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n487_), .A2(new_n488_), .B1(new_n472_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n486_), .B1(new_n492_), .B2(new_n462_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G113gat), .B(G141gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G169gat), .B(G197gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n486_), .B(new_n498_), .C1(new_n492_), .C2(new_n462_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n202_), .B1(new_n460_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n458_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT104), .B(new_n500_), .C1(new_n503_), .C2(new_n446_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT37), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT76), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT77), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G232gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT34), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT35), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT70), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT75), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT70), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n511_), .A2(new_n515_), .A3(KEYINPUT35), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n513_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n514_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n520_), .B(new_n521_), .C1(G99gat), .C2(G106gat), .ZN(new_n522_));
  INV_X1    g321(.A(G106gat), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n237_), .B(new_n523_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT67), .B1(new_n536_), .B2(new_n531_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n530_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT65), .B1(new_n527_), .B2(new_n528_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G99gat), .A2(G106gat), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT65), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n526_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n540_), .A2(new_n525_), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT8), .B1(new_n535_), .B2(new_n537_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n539_), .A2(KEYINPUT8), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT10), .B(G99gat), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n540_), .B(new_n545_), .C1(G106gat), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT9), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n534_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT64), .B(G92gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(G85gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n532_), .A2(KEYINPUT9), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n552_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n548_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n475_), .B(new_n489_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n519_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n539_), .A2(KEYINPUT8), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n547_), .A2(new_n546_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n550_), .A2(new_n556_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n475_), .A3(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n511_), .A2(KEYINPUT35), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n560_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n513_), .A2(new_n516_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT72), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n571_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n566_), .B1(new_n558_), .B2(new_n475_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n563_), .A2(new_n564_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(KEYINPUT72), .A3(new_n491_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n569_), .B1(new_n570_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT73), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT36), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n576_), .A2(new_n570_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n569_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(KEYINPUT74), .A3(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n581_), .A2(KEYINPUT36), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n577_), .A2(KEYINPUT74), .A3(new_n587_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n583_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n506_), .A2(KEYINPUT76), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n509_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n577_), .A2(new_n582_), .ZN(new_n594_));
  AND4_X1   g393(.A1(KEYINPUT74), .A2(new_n584_), .A3(new_n585_), .A4(new_n587_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n587_), .B1(new_n577_), .B2(KEYINPUT74), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n592_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n508_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n593_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G57gat), .B(G64gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT69), .ZN(new_n602_));
  INV_X1    g401(.A(G71gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT68), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT68), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G71gat), .ZN(new_n606_));
  INV_X1    g405(.A(G78gat), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n602_), .A2(KEYINPUT11), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT69), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n601_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT11), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n614_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n604_), .A2(new_n606_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(G78gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(KEYINPUT11), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n613_), .A2(new_n615_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n611_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(new_n483_), .ZN(new_n624_));
  XOR2_X1   g423(.A(G127gat), .B(G155gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n624_), .A2(KEYINPUT17), .A3(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(KEYINPUT17), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n624_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n600_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G230gat), .A2(G233gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n621_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n611_), .B(new_n620_), .C1(new_n548_), .C2(new_n557_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(KEYINPUT12), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT12), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n574_), .A2(new_n640_), .A3(new_n611_), .A4(new_n620_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n635_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G120gat), .B(G148gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT5), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n647_), .B(new_n648_), .Z(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n643_), .A2(new_n645_), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT13), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n634_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n457_), .A2(KEYINPUT105), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n381_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(new_n466_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n505_), .A2(new_n656_), .A3(new_n662_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n663_), .A2(KEYINPUT106), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(KEYINPUT106), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(KEYINPUT38), .A3(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n460_), .A2(new_n597_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n633_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n655_), .A2(new_n501_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n670_), .B2(new_n457_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n666_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT38), .B1(new_n664_), .B2(new_n665_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT107), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n673_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n675_), .A2(new_n676_), .A3(new_n671_), .A4(new_n666_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(G1324gat));
  NAND2_X1  g477(.A1(new_n453_), .A2(new_n456_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G8gat), .B1(new_n670_), .B2(new_n680_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT39), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n681_), .A2(KEYINPUT39), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n505_), .A2(new_n656_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(new_n467_), .ZN(new_n686_));
  OAI22_X1  g485(.A1(new_n683_), .A2(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n670_), .B2(new_n447_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT41), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n685_), .A2(G15gat), .A3(new_n447_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1326gat));
  NOR2_X1   g492(.A1(new_n448_), .A2(new_n449_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G22gat), .B1(new_n670_), .B2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n464_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n685_), .B2(new_n699_), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n668_), .A2(new_n597_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n655_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT110), .B1(new_n505_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704_));
  INV_X1    g503(.A(new_n702_), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n704_), .B(new_n705_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n703_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G29gat), .B1(new_n707_), .B2(new_n381_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n600_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n503_), .B2(new_n446_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT43), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT109), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(new_n713_), .A3(KEYINPUT43), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n715_), .B(new_n709_), .C1(new_n503_), .C2(new_n446_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n712_), .A2(new_n714_), .A3(new_n716_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n655_), .A2(new_n501_), .A3(new_n633_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(KEYINPUT44), .A3(new_n718_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n719_), .A2(G29gat), .A3(new_n661_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n718_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n708_), .B1(new_n720_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n680_), .A2(G36gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n707_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n727_), .ZN(new_n729_));
  NOR4_X1   g528(.A1(new_n703_), .A2(new_n706_), .A3(KEYINPUT45), .A4(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n718_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n716_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(KEYINPUT109), .B2(new_n711_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n735_), .B2(new_n714_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n680_), .B1(new_n736_), .B2(KEYINPUT44), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n732_), .B1(new_n737_), .B2(new_n723_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n725_), .B1(new_n731_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n703_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n706_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n727_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT45), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n707_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n719_), .A2(new_n679_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n736_), .A2(KEYINPUT44), .ZN(new_n747_));
  OAI21_X1  g546(.A(G36gat), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(new_n748_), .A3(KEYINPUT46), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n739_), .A2(new_n749_), .ZN(G1329gat));
  NAND2_X1  g549(.A1(new_n707_), .A2(new_n259_), .ZN(new_n751_));
  INV_X1    g550(.A(G43gat), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n723_), .A2(G43gat), .A3(new_n259_), .A4(new_n719_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT47), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n753_), .A2(new_n754_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1330gat));
  AOI21_X1  g558(.A(G50gat), .B1(new_n707_), .B2(new_n698_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n719_), .A2(G50gat), .A3(new_n698_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n723_), .ZN(G1331gat));
  NOR2_X1   g561(.A1(new_n460_), .A2(new_n500_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n634_), .A2(new_n654_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT111), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G57gat), .B1(new_n767_), .B2(new_n661_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n667_), .A2(new_n501_), .A3(new_n655_), .A4(new_n633_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT112), .B(G57gat), .Z(new_n770_));
  NOR3_X1   g569(.A1(new_n769_), .A2(new_n457_), .A3(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n768_), .A2(new_n771_), .ZN(G1332gat));
  OAI21_X1  g571(.A(G64gat), .B1(new_n769_), .B2(new_n680_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT48), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n680_), .A2(G64gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n766_), .B2(new_n775_), .ZN(G1333gat));
  OAI21_X1  g575(.A(G71gat), .B1(new_n769_), .B2(new_n447_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT49), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n767_), .A2(new_n603_), .A3(new_n259_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1334gat));
  OAI21_X1  g579(.A(G78gat), .B1(new_n769_), .B2(new_n694_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT50), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n767_), .A2(new_n607_), .A3(new_n698_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1335gat));
  NOR2_X1   g583(.A1(new_n701_), .A2(new_n654_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n763_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(G85gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n661_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n717_), .A2(KEYINPUT113), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n735_), .A2(new_n791_), .A3(new_n714_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n655_), .A2(new_n501_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(new_n633_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n790_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n795_), .A2(new_n381_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n789_), .B1(new_n796_), .B2(new_n788_), .ZN(G1336gat));
  AOI21_X1  g596(.A(G92gat), .B1(new_n787_), .B2(new_n679_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n679_), .A2(new_n553_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n795_), .B2(new_n799_), .ZN(G1337gat));
  NAND4_X1  g599(.A1(new_n790_), .A2(new_n792_), .A3(new_n259_), .A4(new_n794_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G99gat), .ZN(new_n802_));
  OR3_X1    g601(.A1(new_n786_), .A2(new_n447_), .A3(new_n549_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT51), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n802_), .A2(new_n806_), .A3(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1338gat));
  XNOR2_X1  g607(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811_));
  OAI21_X1  g610(.A(G106gat), .B1(new_n811_), .B2(KEYINPUT114), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n694_), .A2(new_n793_), .A3(new_n633_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n717_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(KEYINPUT114), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n787_), .A2(new_n523_), .A3(new_n698_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n810_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n814_), .A2(new_n815_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n821_), .A2(new_n816_), .A3(new_n818_), .A4(new_n809_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1339gat));
  NAND4_X1  g622(.A1(new_n600_), .A2(new_n501_), .A3(new_n654_), .A4(new_n633_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n639_), .A2(new_n641_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n635_), .ZN(new_n831_));
  AOI211_X1 g630(.A(KEYINPUT55), .B(new_n636_), .C1(new_n639_), .C2(new_n641_), .ZN(new_n832_));
  OAI22_X1  g631(.A1(new_n831_), .A2(new_n832_), .B1(new_n635_), .B2(new_n830_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n649_), .A3(new_n834_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n642_), .A2(new_n644_), .A3(new_n649_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n499_), .B2(new_n497_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n834_), .B1(new_n833_), .B2(new_n649_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n828_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n833_), .A2(new_n649_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n834_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n843_), .A2(KEYINPUT117), .A3(new_n835_), .A4(new_n837_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n496_), .B1(new_n492_), .B2(new_n462_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n477_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n461_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n493_), .A2(new_n496_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n848_), .A2(new_n653_), .A3(KEYINPUT118), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT118), .B1(new_n848_), .B2(new_n653_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n840_), .A2(new_n844_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n591_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT57), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n855_), .A3(new_n591_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n841_), .A2(KEYINPUT56), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT56), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n833_), .A2(new_n858_), .A3(new_n649_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n857_), .A2(new_n651_), .A3(new_n848_), .A4(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(KEYINPUT119), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(KEYINPUT119), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n600_), .B1(new_n863_), .B2(KEYINPUT58), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n854_), .A2(new_n856_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n827_), .B1(new_n865_), .B2(new_n633_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n451_), .A2(new_n679_), .A3(new_n660_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n865_), .A2(KEYINPUT120), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n668_), .B1(new_n865_), .B2(KEYINPUT120), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n827_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n873_), .A2(new_n868_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n869_), .B1(new_n874_), .B2(new_n867_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875_), .B2(new_n501_), .ZN(new_n876_));
  INV_X1    g675(.A(G113gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n877_), .A3(new_n500_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1340gat));
  OAI21_X1  g678(.A(G120gat), .B1(new_n875_), .B2(new_n654_), .ZN(new_n880_));
  INV_X1    g679(.A(G120gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n654_), .B2(KEYINPUT60), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n874_), .B(new_n882_), .C1(KEYINPUT60), .C2(new_n881_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(G1341gat));
  OAI21_X1  g683(.A(G127gat), .B1(new_n875_), .B2(new_n668_), .ZN(new_n885_));
  INV_X1    g684(.A(G127gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n874_), .A2(new_n886_), .A3(new_n633_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1342gat));
  OAI21_X1  g687(.A(G134gat), .B1(new_n875_), .B2(new_n600_), .ZN(new_n889_));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n874_), .A2(new_n890_), .A3(new_n597_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1343gat));
  INV_X1    g691(.A(new_n450_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n873_), .A2(new_n893_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n894_), .A2(new_n679_), .A3(new_n660_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n500_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n655_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n633_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT61), .B(G155gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  INV_X1    g701(.A(G162gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n895_), .A2(new_n903_), .A3(new_n597_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n895_), .A2(new_n709_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n903_), .ZN(G1347gat));
  NAND2_X1  g705(.A1(new_n864_), .A2(new_n862_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n852_), .A2(new_n855_), .A3(new_n591_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n855_), .B1(new_n852_), .B2(new_n591_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n907_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n826_), .B1(new_n910_), .B2(new_n668_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n447_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n912_), .A2(new_n913_), .A3(new_n679_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n912_), .B2(new_n679_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n694_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n911_), .A2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n216_), .B1(new_n917_), .B2(new_n500_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT62), .Z(new_n919_));
  INV_X1    g718(.A(new_n916_), .ZN(new_n920_));
  AOI21_X1  g719(.A(KEYINPUT122), .B1(new_n866_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n911_), .A2(new_n922_), .A3(new_n916_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n921_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n925_), .A2(new_n265_), .A3(new_n500_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n919_), .A2(new_n926_), .ZN(G1348gat));
  AND2_X1   g726(.A1(new_n873_), .A2(new_n694_), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n914_), .A2(new_n915_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n928_), .A2(G176gat), .A3(new_n655_), .A4(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n655_), .B1(new_n921_), .B2(new_n923_), .ZN(new_n931_));
  AOI21_X1  g730(.A(KEYINPUT123), .B1(new_n931_), .B2(new_n214_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n922_), .B1(new_n911_), .B2(new_n916_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n854_), .A2(new_n856_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n633_), .B1(new_n934_), .B2(new_n907_), .ZN(new_n935_));
  OAI211_X1 g734(.A(KEYINPUT122), .B(new_n920_), .C1(new_n935_), .C2(new_n826_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n654_), .B1(new_n933_), .B2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n937_), .A2(new_n938_), .A3(G176gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n930_), .B1(new_n932_), .B2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n930_), .B(KEYINPUT124), .C1(new_n932_), .C2(new_n939_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1349gat));
  NOR3_X1   g743(.A1(new_n924_), .A2(new_n221_), .A3(new_n668_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n928_), .A2(new_n633_), .A3(new_n929_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n205_), .B2(new_n946_), .ZN(G1350gat));
  OAI21_X1  g746(.A(G190gat), .B1(new_n924_), .B2(new_n600_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n597_), .A2(new_n222_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n924_), .B2(new_n949_), .ZN(G1351gat));
  NOR2_X1   g749(.A1(new_n680_), .A2(new_n381_), .ZN(new_n951_));
  NAND4_X1  g750(.A1(new_n873_), .A2(new_n893_), .A3(new_n500_), .A4(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(G197gat), .ZN(new_n953_));
  AND3_X1   g752(.A1(new_n952_), .A2(KEYINPUT125), .A3(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(KEYINPUT125), .B1(new_n952_), .B2(new_n953_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n952_), .A2(new_n953_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n954_), .A2(new_n955_), .A3(new_n956_), .ZN(G1352gat));
  INV_X1    g756(.A(new_n951_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n894_), .A2(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n654_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n962_));
  XOR2_X1   g761(.A(new_n961_), .B(new_n962_), .Z(G1353gat));
  NAND2_X1  g762(.A1(new_n959_), .A2(new_n633_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(KEYINPUT63), .B(G211gat), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(new_n964_), .B2(new_n967_), .ZN(G1354gat));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n969_));
  NOR3_X1   g768(.A1(new_n894_), .A2(new_n600_), .A3(new_n958_), .ZN(new_n970_));
  INV_X1    g769(.A(G218gat), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  NOR4_X1   g771(.A1(new_n894_), .A2(G218gat), .A3(new_n591_), .A4(new_n958_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n969_), .B1(new_n972_), .B2(new_n973_), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n959_), .A2(new_n971_), .A3(new_n597_), .ZN(new_n975_));
  OAI211_X1 g774(.A(new_n975_), .B(KEYINPUT127), .C1(new_n970_), .C2(new_n971_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n974_), .A2(new_n976_), .ZN(G1355gat));
endmodule


