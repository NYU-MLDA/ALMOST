//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n967_, new_n969_, new_n970_, new_n971_, new_n972_, new_n974_,
    new_n975_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n988_,
    new_n990_, new_n991_, new_n993_, new_n994_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1018_,
    new_n1019_, new_n1020_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XOR2_X1   g001(.A(G8gat), .B(G36gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G64gat), .B(G92gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT92), .ZN(new_n208_));
  INV_X1    g007(.A(G197gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(G204gat), .ZN(new_n210_));
  INV_X1    g009(.A(G204gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G197gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT92), .B1(new_n211_), .B2(G197gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G211gat), .B(G218gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n209_), .A2(G204gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n212_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT21), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n214_), .A2(new_n210_), .A3(new_n217_), .A4(new_n212_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT93), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n222_), .B(new_n216_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n223_), .A2(new_n224_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n219_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT94), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G183gat), .ZN(new_n230_));
  INV_X1    g029(.A(G190gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT23), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT83), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(G183gat), .A3(G190gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n234_), .A2(KEYINPUT83), .A3(G183gat), .A4(G190gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT79), .B(G190gat), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n236_), .B(new_n237_), .C1(G183gat), .C2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT80), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(G169gat), .A3(G176gat), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G176gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT22), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G169gat), .ZN(new_n247_));
  INV_X1    g046(.A(G169gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT81), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G169gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n246_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n245_), .B(new_n247_), .C1(new_n252_), .C2(KEYINPUT82), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n251_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT22), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT82), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n239_), .B(new_n244_), .C1(new_n253_), .C2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n244_), .A2(new_n260_), .ZN(new_n261_));
  NOR3_X1   g060(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(new_n238_), .B2(KEYINPUT26), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n230_), .A2(KEYINPUT25), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G183gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n261_), .B(new_n263_), .C1(new_n265_), .C2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n258_), .A2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n219_), .B(KEYINPUT94), .C1(new_n225_), .C2(new_n226_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n229_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G226gat), .A2(G233gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT19), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT20), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n248_), .A2(KEYINPUT22), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n247_), .A2(new_n277_), .A3(new_n245_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n244_), .A2(new_n278_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n232_), .A2(new_n235_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT97), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n232_), .A2(new_n235_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n230_), .A2(new_n231_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT97), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(new_n244_), .A4(new_n278_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n236_), .A2(new_n237_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n262_), .B1(new_n260_), .B2(new_n240_), .ZN(new_n288_));
  AND2_X1   g087(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n266_), .B(new_n268_), .C1(new_n289_), .C2(new_n264_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n281_), .A2(new_n286_), .B1(new_n287_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n216_), .B1(new_n293_), .B2(new_n217_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n223_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(KEYINPUT93), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n223_), .A2(new_n224_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n296_), .A2(new_n297_), .B1(new_n215_), .B2(new_n218_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n276_), .B1(new_n292_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT98), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n273_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n241_), .A2(new_n243_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n247_), .A2(new_n245_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n252_), .A2(KEYINPUT82), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n302_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n265_), .A2(new_n269_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n261_), .A2(new_n263_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n306_), .A2(new_n239_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n272_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n213_), .A2(KEYINPUT93), .A3(new_n217_), .A4(new_n214_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n294_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(new_n297_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT94), .B1(new_n313_), .B2(new_n219_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n309_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n281_), .A2(new_n286_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n288_), .A2(new_n236_), .A3(new_n237_), .A4(new_n290_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n316_), .B1(new_n319_), .B2(new_n227_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n275_), .B1(new_n315_), .B2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n301_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n273_), .A2(new_n299_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT98), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n207_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n275_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n271_), .B1(new_n229_), .B2(new_n272_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT20), .B1(new_n292_), .B2(new_n298_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n273_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n324_), .A2(new_n329_), .A3(new_n207_), .A4(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n202_), .B1(new_n325_), .B2(new_n332_), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n327_), .A2(new_n328_), .A3(new_n326_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n284_), .A2(new_n244_), .A3(new_n278_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(KEYINPUT104), .A3(new_n318_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT104), .B1(new_n335_), .B2(new_n318_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n227_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT105), .B1(new_n339_), .B2(new_n316_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n338_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n298_), .A3(new_n336_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT105), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(KEYINPUT20), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n273_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n334_), .B1(new_n345_), .B2(new_n326_), .ZN(new_n346_));
  OAI211_X1 g145(.A(KEYINPUT27), .B(new_n331_), .C1(new_n346_), .C2(new_n207_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n333_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G134gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G127gat), .ZN(new_n353_));
  INV_X1    g152(.A(G127gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G134gat), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n353_), .A2(new_n355_), .A3(new_n350_), .ZN(new_n356_));
  INV_X1    g155(.A(G120gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G113gat), .ZN(new_n358_));
  INV_X1    g157(.A(G113gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G120gat), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n358_), .A2(new_n360_), .A3(KEYINPUT86), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT86), .B1(new_n358_), .B2(new_n360_), .ZN(new_n362_));
  OAI22_X1  g161(.A1(new_n351_), .A2(new_n356_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT87), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n362_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n353_), .A2(new_n355_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT85), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n349_), .A2(new_n350_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n358_), .A2(new_n360_), .A3(KEYINPUT86), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n366_), .A2(new_n368_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n365_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT31), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT84), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G227gat), .A2(G233gat), .ZN(new_n377_));
  INV_X1    g176(.A(G15gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT30), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n309_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n376_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G71gat), .B(G99gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G43gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n382_), .B(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G141gat), .A2(G148gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G141gat), .A2(G148gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(KEYINPUT1), .B2(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n390_), .A2(KEYINPUT1), .ZN(new_n392_));
  AOI211_X1 g191(.A(new_n387_), .B(new_n388_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(new_n371_), .B2(new_n363_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT90), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT2), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n386_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n386_), .A2(KEYINPUT89), .A3(new_n396_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT88), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n387_), .A2(KEYINPUT2), .B1(new_n388_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT88), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n388_), .B2(new_n403_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n401_), .A2(new_n402_), .A3(new_n404_), .A4(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G155gat), .B(G162gat), .Z(new_n408_));
  AOI21_X1  g207(.A(new_n395_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n388_), .A2(new_n403_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n406_), .A2(new_n402_), .A3(new_n410_), .A4(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n386_), .A2(KEYINPUT89), .A3(new_n396_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT89), .B1(new_n386_), .B2(new_n396_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n395_), .B(new_n408_), .C1(new_n412_), .C2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n394_), .B1(new_n409_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT100), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n393_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(new_n409_), .B2(new_n417_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n373_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n408_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT90), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n416_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(KEYINPUT100), .A3(new_n394_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n420_), .A2(new_n423_), .A3(KEYINPUT4), .A4(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT101), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n426_), .A2(new_n421_), .B1(new_n365_), .B2(new_n372_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n428_), .A2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n420_), .A2(new_n423_), .A3(new_n429_), .A4(new_n427_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(G85gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT0), .B(G57gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT106), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n435_), .A2(new_n436_), .A3(new_n441_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n437_), .A2(KEYINPUT106), .A3(new_n442_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OR3_X1    g247(.A1(new_n422_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT28), .B1(new_n422_), .B2(KEYINPUT29), .ZN(new_n450_));
  XOR2_X1   g249(.A(G22gat), .B(G50gat), .Z(new_n451_));
  AND3_X1   g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G228gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT91), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n422_), .B2(KEYINPUT29), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT95), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n229_), .A2(new_n272_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n458_), .A2(new_n459_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n393_), .B1(new_n425_), .B2(new_n416_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT29), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n456_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT95), .B1(new_n465_), .B2(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n462_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G78gat), .B(G106gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n468_), .B(KEYINPUT96), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n227_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n457_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n467_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n470_), .B1(new_n467_), .B2(new_n472_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n454_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n459_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n465_), .A2(KEYINPUT95), .A3(new_n460_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n472_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n469_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n452_), .A2(new_n453_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n467_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n475_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n348_), .A2(new_n385_), .A3(new_n448_), .A4(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n420_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n441_), .B1(new_n486_), .B2(new_n430_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT102), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n432_), .A2(new_n433_), .B1(G225gat), .B2(G233gat), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n428_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n488_), .B1(new_n428_), .B2(new_n489_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n487_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT103), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n445_), .A2(KEYINPUT33), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT33), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n435_), .A2(new_n495_), .A3(new_n436_), .A4(new_n441_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n325_), .A2(new_n332_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT103), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n499_), .B(new_n487_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n493_), .A2(new_n497_), .A3(new_n498_), .A4(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n207_), .A2(KEYINPUT32), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n322_), .A2(new_n502_), .A3(new_n324_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n345_), .A2(new_n326_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n334_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n502_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n446_), .A2(new_n447_), .A3(new_n503_), .A4(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n501_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n483_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n483_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(new_n448_), .A3(new_n348_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n385_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n485_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT13), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT9), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G85gat), .B(G92gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT65), .B(G85gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(G92gat), .ZN(new_n521_));
  OAI22_X1  g320(.A1(new_n518_), .A2(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT66), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT66), .ZN(new_n524_));
  OAI221_X1 g323(.A(new_n524_), .B1(new_n519_), .B2(new_n518_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n525_));
  OR2_X1    g324(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT64), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT6), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n530_), .B2(new_n529_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n523_), .A2(new_n525_), .A3(new_n531_), .A4(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n519_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT7), .ZN(new_n538_));
  INV_X1    g337(.A(G99gat), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(new_n527_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n537_), .B1(new_n534_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n544_), .B(new_n537_), .C1(new_n534_), .C2(new_n542_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n536_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT69), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n536_), .A2(new_n548_), .A3(KEYINPUT69), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT68), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n553_), .A2(new_n556_), .A3(KEYINPUT11), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n559_));
  XOR2_X1   g358(.A(G71gat), .B(G78gat), .Z(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n555_), .A2(new_n559_), .A3(new_n560_), .A4(new_n557_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n551_), .A2(KEYINPUT12), .A3(new_n552_), .A4(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT12), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n536_), .A2(new_n548_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n567_), .B1(new_n568_), .B2(new_n564_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n564_), .A2(new_n548_), .A3(new_n536_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n566_), .A2(new_n569_), .A3(new_n570_), .A4(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n570_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n571_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n564_), .B1(new_n548_), .B2(new_n536_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT5), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n578_), .B(new_n579_), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n572_), .A2(new_n576_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n517_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n572_), .A2(new_n576_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n580_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n572_), .A2(new_n576_), .A3(new_n581_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(KEYINPUT13), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT70), .ZN(new_n591_));
  XOR2_X1   g390(.A(G1gat), .B(G8gat), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G15gat), .B(G22gat), .ZN(new_n594_));
  INV_X1    g393(.A(G1gat), .ZN(new_n595_));
  INV_X1    g394(.A(G8gat), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT14), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n592_), .A2(new_n597_), .A3(new_n594_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G29gat), .B(G36gat), .Z(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(KEYINPUT71), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G29gat), .B(G36gat), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT71), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G43gat), .B(G50gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n603_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n602_), .A2(KEYINPUT71), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n605_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n607_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT15), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n609_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n608_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n610_), .A2(new_n611_), .A3(new_n607_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT15), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n601_), .B1(new_n614_), .B2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n615_), .A2(new_n616_), .A3(new_n599_), .A4(new_n600_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n601_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n619_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n620_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT76), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT76), .ZN(new_n627_));
  AOI211_X1 g426(.A(new_n627_), .B(new_n620_), .C1(new_n623_), .C2(new_n619_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n622_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT77), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT77), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n622_), .B(new_n631_), .C1(new_n626_), .C2(new_n628_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G169gat), .B(G197gat), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n633_), .B(new_n634_), .Z(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n630_), .A2(new_n632_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT78), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n630_), .A2(KEYINPUT78), .A3(new_n632_), .A4(new_n636_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n629_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n635_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n640_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n591_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n516_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT74), .ZN(new_n649_));
  INV_X1    g448(.A(new_n617_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n615_), .A2(KEYINPUT15), .A3(new_n616_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n551_), .A2(new_n652_), .A3(new_n552_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n615_), .A2(new_n616_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT35), .ZN(new_n656_));
  NAND2_X1  g455(.A1(G232gat), .A2(G233gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT34), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n568_), .A2(new_n655_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n656_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n653_), .A2(new_n660_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n653_), .B2(new_n660_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n649_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n653_), .A2(new_n660_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n661_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(KEYINPUT74), .A3(new_n663_), .ZN(new_n669_));
  XOR2_X1   g468(.A(G190gat), .B(G218gat), .Z(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT72), .ZN(new_n671_));
  XNOR2_X1  g470(.A(G134gat), .B(G162gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT36), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n666_), .A2(new_n669_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT37), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT36), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n673_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT73), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n668_), .A2(new_n663_), .A3(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n675_), .A2(new_n676_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT75), .ZN(new_n682_));
  INV_X1    g481(.A(new_n680_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n674_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n668_), .B2(new_n663_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT37), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n681_), .A2(new_n682_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n682_), .B1(new_n681_), .B2(new_n686_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(G231gat), .A2(G233gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n601_), .B(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(new_n564_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT17), .ZN(new_n693_));
  XOR2_X1   g492(.A(G127gat), .B(G155gat), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT16), .ZN(new_n695_));
  XNOR2_X1  g494(.A(G183gat), .B(G211gat), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n692_), .A2(new_n693_), .A3(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n693_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n692_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n689_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n648_), .A2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n446_), .A2(new_n447_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n595_), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n675_), .A2(new_n680_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NOR4_X1   g507(.A1(new_n516_), .A2(new_n647_), .A3(new_n708_), .A4(new_n702_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(new_n705_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n710_), .B2(new_n595_), .ZN(new_n711_));
  MUX2_X1   g510(.A(new_n706_), .B(new_n711_), .S(KEYINPUT38), .Z(G1324gat));
  INV_X1    g511(.A(new_n348_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n704_), .A2(new_n596_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT39), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n709_), .A2(new_n713_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(G8gat), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT39), .B(new_n596_), .C1(new_n709_), .C2(new_n713_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT40), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(G1325gat));
  AOI21_X1  g520(.A(new_n378_), .B1(new_n709_), .B2(new_n385_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT41), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n704_), .A2(new_n378_), .A3(new_n385_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1326gat));
  INV_X1    g524(.A(G22gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n709_), .B2(new_n512_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n704_), .A2(new_n726_), .A3(new_n512_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1327gat));
  NOR2_X1   g530(.A1(new_n707_), .A2(new_n701_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n648_), .A2(new_n732_), .ZN(new_n733_));
  OR3_X1    g532(.A1(new_n733_), .A2(G29gat), .A3(new_n448_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n647_), .A2(new_n701_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n687_), .A2(new_n688_), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT43), .B1(new_n516_), .B2(new_n737_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n501_), .A2(new_n509_), .B1(new_n482_), .B2(new_n475_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n475_), .A2(new_n333_), .A3(new_n482_), .A4(new_n347_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n705_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n515_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n484_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n689_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n736_), .B1(new_n738_), .B2(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(KEYINPUT44), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(new_n448_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n743_), .B2(new_n689_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT43), .B(new_n737_), .C1(new_n742_), .C2(new_n484_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT44), .B(new_n735_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT108), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n738_), .A2(new_n745_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(KEYINPUT44), .A4(new_n735_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n748_), .A2(KEYINPUT109), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(G29gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT109), .B1(new_n748_), .B2(new_n756_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n734_), .B1(new_n758_), .B2(new_n759_), .ZN(G1328gat));
  INV_X1    g559(.A(KEYINPUT46), .ZN(new_n761_));
  INV_X1    g560(.A(G36gat), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n753_), .A2(new_n735_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n348_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n762_), .B1(new_n756_), .B2(new_n765_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n648_), .A2(new_n762_), .A3(new_n713_), .A4(new_n732_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT45), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n761_), .B1(new_n766_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n713_), .B1(new_n746_), .B2(KEYINPUT44), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n752_), .B2(new_n755_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT46), .B(new_n768_), .C1(new_n772_), .C2(new_n762_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(G1329gat));
  NAND2_X1  g573(.A1(new_n763_), .A2(new_n764_), .ZN(new_n775_));
  INV_X1    g574(.A(G43gat), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n515_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n754_), .B1(new_n746_), .B2(KEYINPUT44), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n751_), .A2(KEYINPUT108), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n775_), .B(new_n777_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n733_), .B2(new_n515_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT110), .B(new_n776_), .C1(new_n733_), .C2(new_n515_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n780_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT47), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n780_), .A2(new_n788_), .A3(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1330gat));
  INV_X1    g589(.A(new_n733_), .ZN(new_n791_));
  AOI21_X1  g590(.A(G50gat), .B1(new_n791_), .B2(new_n512_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n747_), .B1(new_n752_), .B2(new_n755_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n512_), .A2(G50gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(G1331gat));
  NOR2_X1   g594(.A1(new_n516_), .A2(new_n708_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n591_), .A2(new_n702_), .A3(new_n646_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(G57gat), .B1(new_n799_), .B2(new_n448_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n516_), .A2(new_n646_), .A3(new_n591_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n801_), .A2(new_n703_), .ZN(new_n802_));
  INV_X1    g601(.A(G57gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n705_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(new_n804_), .ZN(G1332gat));
  NOR2_X1   g604(.A1(new_n348_), .A2(G64gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT111), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n802_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(G64gat), .B1(new_n799_), .B2(new_n348_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(KEYINPUT48), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(KEYINPUT48), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n808_), .B1(new_n810_), .B2(new_n811_), .ZN(G1333gat));
  INV_X1    g611(.A(G71gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n385_), .A2(new_n813_), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n814_), .B(KEYINPUT112), .Z(new_n815_));
  NAND2_X1  g614(.A1(new_n802_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n798_), .A2(new_n385_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(G71gat), .ZN(new_n819_));
  AOI211_X1 g618(.A(KEYINPUT49), .B(new_n813_), .C1(new_n798_), .C2(new_n385_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT113), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n823_), .B(new_n816_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1334gat));
  INV_X1    g624(.A(G78gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n798_), .B2(new_n512_), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT50), .Z(new_n828_));
  NAND3_X1  g627(.A1(new_n802_), .A2(new_n826_), .A3(new_n512_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1335gat));
  AND2_X1   g629(.A1(new_n801_), .A2(new_n732_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G85gat), .B1(new_n831_), .B2(new_n705_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n591_), .A2(new_n701_), .A3(new_n646_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n753_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n448_), .A2(new_n520_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n834_), .B2(new_n835_), .ZN(G1336gat));
  INV_X1    g635(.A(G92gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n831_), .A2(new_n837_), .A3(new_n713_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n713_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n840_), .B2(new_n837_), .ZN(G1337gat));
  AOI21_X1  g640(.A(new_n539_), .B1(new_n834_), .B2(new_n385_), .ZN(new_n842_));
  AND4_X1   g641(.A1(new_n526_), .A2(new_n831_), .A3(new_n528_), .A4(new_n385_), .ZN(new_n843_));
  OR3_X1    g642(.A1(new_n842_), .A2(new_n843_), .A3(KEYINPUT51), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT51), .B1(new_n842_), .B2(new_n843_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1338gat));
  NAND3_X1  g645(.A1(new_n831_), .A2(new_n527_), .A3(new_n512_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n753_), .A2(new_n512_), .A3(new_n833_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n848_), .A2(new_n849_), .A3(G106gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n848_), .B2(G106gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n847_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT53), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n854_), .B(new_n847_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1339gat));
  NOR3_X1   g655(.A1(new_n713_), .A2(new_n515_), .A3(new_n448_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n641_), .A2(new_n643_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n582_), .B1(new_n858_), .B2(new_n639_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n564_), .A2(new_n567_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n551_), .A2(new_n552_), .A3(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n571_), .B1(new_n575_), .B2(KEYINPUT12), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n573_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT55), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n572_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n861_), .A2(new_n862_), .A3(new_n866_), .A4(new_n573_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n865_), .A2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT56), .B1(new_n869_), .B2(new_n580_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT56), .ZN(new_n871_));
  AOI211_X1 g670(.A(new_n871_), .B(new_n581_), .C1(new_n865_), .C2(new_n868_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n859_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n618_), .A2(new_n619_), .A3(new_n625_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n635_), .B1(new_n624_), .B2(new_n620_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n642_), .A2(new_n635_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n878_), .B2(new_n707_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880_));
  AOI211_X1 g679(.A(new_n880_), .B(new_n708_), .C1(new_n873_), .C2(new_n877_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n876_), .A2(new_n587_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT116), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n876_), .A2(new_n885_), .A3(new_n587_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n572_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(KEYINPUT55), .B2(new_n863_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n580_), .B1(new_n889_), .B2(new_n867_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n871_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n869_), .A2(KEYINPUT56), .A3(new_n580_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n887_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT58), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n870_), .A2(new_n872_), .ZN(new_n897_));
  OAI211_X1 g696(.A(KEYINPUT117), .B(new_n896_), .C1(new_n897_), .C2(new_n887_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(new_n898_), .A3(new_n689_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n701_), .B1(new_n882_), .B2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT115), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n639_), .A2(new_n701_), .A3(new_n643_), .A4(new_n641_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n589_), .B1(KEYINPUT114), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n858_), .A2(new_n904_), .A3(new_n701_), .A4(new_n639_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n901_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n902_), .A2(KEYINPUT114), .ZN(new_n907_));
  AND4_X1   g706(.A1(new_n901_), .A2(new_n907_), .A3(new_n590_), .A4(new_n905_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n737_), .B1(new_n906_), .B2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(KEYINPUT54), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n907_), .A2(new_n590_), .A3(new_n905_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT115), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n903_), .A2(new_n901_), .A3(new_n905_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n911_), .B1(new_n915_), .B2(new_n737_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n910_), .A2(new_n916_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n483_), .B(new_n857_), .C1(new_n900_), .C2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n919_), .A2(new_n359_), .A3(new_n646_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n587_), .B1(new_n640_), .B2(new_n644_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n877_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n707_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n880_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n878_), .A2(KEYINPUT57), .A3(new_n707_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n899_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n702_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n909_), .A2(KEYINPUT54), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n915_), .A2(new_n911_), .A3(new_n737_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n512_), .B1(new_n930_), .B2(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n934_), .A2(KEYINPUT59), .A3(new_n857_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n645_), .B1(new_n922_), .B2(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n920_), .B1(new_n936_), .B2(new_n359_), .ZN(G1340gat));
  OAI21_X1  g736(.A(new_n357_), .B1(new_n591_), .B2(KEYINPUT60), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n919_), .B(new_n938_), .C1(KEYINPUT60), .C2(new_n357_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n591_), .B1(new_n922_), .B2(new_n935_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n357_), .ZN(G1341gat));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n942_));
  AND2_X1   g741(.A1(new_n354_), .A2(KEYINPUT118), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n354_), .A2(KEYINPUT118), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n701_), .B2(new_n944_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n945_), .B1(new_n922_), .B2(new_n935_), .ZN(new_n946_));
  AOI21_X1  g745(.A(G127gat), .B1(new_n919_), .B2(new_n701_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n942_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n945_), .ZN(new_n949_));
  AOI21_X1  g748(.A(KEYINPUT59), .B1(new_n934_), .B2(new_n857_), .ZN(new_n950_));
  AOI22_X1  g749(.A1(new_n929_), .A2(new_n702_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n857_), .ZN(new_n952_));
  NOR4_X1   g751(.A1(new_n951_), .A2(new_n921_), .A3(new_n512_), .A4(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n949_), .B1(new_n950_), .B2(new_n953_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n354_), .B1(new_n918_), .B2(new_n702_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n954_), .A2(KEYINPUT119), .A3(new_n955_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n948_), .A2(new_n956_), .ZN(G1342gat));
  NAND3_X1  g756(.A1(new_n919_), .A2(new_n352_), .A3(new_n708_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n737_), .B1(new_n922_), .B2(new_n935_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n959_), .B2(new_n352_), .ZN(G1343gat));
  INV_X1    g759(.A(new_n951_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n740_), .A2(new_n385_), .A3(new_n448_), .ZN(new_n962_));
  XOR2_X1   g761(.A(new_n962_), .B(KEYINPUT120), .Z(new_n963_));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n963_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(new_n645_), .ZN(new_n965_));
  XOR2_X1   g764(.A(new_n965_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g765(.A1(new_n964_), .A2(new_n591_), .ZN(new_n967_));
  XOR2_X1   g766(.A(new_n967_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g767(.A1(new_n964_), .A2(new_n702_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(KEYINPUT61), .B(G155gat), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(KEYINPUT121), .ZN(new_n971_));
  XOR2_X1   g770(.A(new_n971_), .B(KEYINPUT122), .Z(new_n972_));
  XNOR2_X1  g771(.A(new_n969_), .B(new_n972_), .ZN(G1346gat));
  OAI21_X1  g772(.A(G162gat), .B1(new_n964_), .B2(new_n737_), .ZN(new_n974_));
  OR2_X1    g773(.A1(new_n707_), .A2(G162gat), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n974_), .B1(new_n964_), .B2(new_n975_), .ZN(G1347gat));
  NOR3_X1   g775(.A1(new_n515_), .A2(new_n348_), .A3(new_n705_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n934_), .A2(new_n977_), .ZN(new_n978_));
  INV_X1    g777(.A(new_n978_), .ZN(new_n979_));
  NAND4_X1  g778(.A1(new_n979_), .A2(new_n247_), .A3(new_n277_), .A4(new_n646_), .ZN(new_n980_));
  INV_X1    g779(.A(new_n934_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n977_), .A2(new_n646_), .ZN(new_n982_));
  XNOR2_X1  g781(.A(new_n982_), .B(KEYINPUT123), .ZN(new_n983_));
  OAI21_X1  g782(.A(G169gat), .B1(new_n981_), .B2(new_n983_), .ZN(new_n984_));
  AND2_X1   g783(.A1(new_n984_), .A2(KEYINPUT62), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n984_), .A2(KEYINPUT62), .ZN(new_n986_));
  OAI21_X1  g785(.A(new_n980_), .B1(new_n985_), .B2(new_n986_), .ZN(G1348gat));
  NOR2_X1   g786(.A1(new_n978_), .A2(new_n591_), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(new_n245_), .ZN(G1349gat));
  NOR2_X1   g788(.A1(new_n978_), .A2(new_n702_), .ZN(new_n990_));
  NOR2_X1   g789(.A1(new_n990_), .A2(G183gat), .ZN(new_n991_));
  AOI21_X1  g790(.A(new_n991_), .B1(new_n269_), .B2(new_n990_), .ZN(G1350gat));
  OAI21_X1  g791(.A(G190gat), .B1(new_n978_), .B2(new_n737_), .ZN(new_n993_));
  OAI21_X1  g792(.A(new_n708_), .B1(new_n264_), .B2(new_n289_), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n993_), .B1(new_n978_), .B2(new_n994_), .ZN(G1351gat));
  INV_X1    g794(.A(KEYINPUT125), .ZN(new_n996_));
  NOR4_X1   g795(.A1(new_n705_), .A2(new_n348_), .A3(new_n385_), .A4(new_n483_), .ZN(new_n997_));
  NAND3_X1  g796(.A1(new_n961_), .A2(new_n646_), .A3(new_n997_), .ZN(new_n998_));
  INV_X1    g797(.A(new_n998_), .ZN(new_n999_));
  OAI21_X1  g798(.A(new_n996_), .B1(new_n999_), .B2(G197gat), .ZN(new_n1000_));
  NAND3_X1  g799(.A1(new_n998_), .A2(KEYINPUT125), .A3(new_n209_), .ZN(new_n1001_));
  NAND3_X1  g800(.A1(new_n999_), .A2(KEYINPUT124), .A3(G197gat), .ZN(new_n1002_));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n1003_));
  OAI21_X1  g802(.A(new_n1003_), .B1(new_n998_), .B2(new_n209_), .ZN(new_n1004_));
  AOI22_X1  g803(.A1(new_n1000_), .A2(new_n1001_), .B1(new_n1002_), .B2(new_n1004_), .ZN(G1352gat));
  NAND2_X1  g804(.A1(new_n961_), .A2(new_n997_), .ZN(new_n1006_));
  NOR2_X1   g805(.A1(new_n1006_), .A2(new_n591_), .ZN(new_n1007_));
  NAND2_X1  g806(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n1008_));
  NAND2_X1  g807(.A1(new_n1007_), .A2(new_n1008_), .ZN(new_n1009_));
  XOR2_X1   g808(.A(KEYINPUT126), .B(G204gat), .Z(new_n1010_));
  OAI21_X1  g809(.A(new_n1009_), .B1(new_n1007_), .B2(new_n1010_), .ZN(G1353gat));
  NOR2_X1   g810(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1012_));
  AND2_X1   g811(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1013_));
  NOR4_X1   g812(.A1(new_n1006_), .A2(new_n702_), .A3(new_n1012_), .A4(new_n1013_), .ZN(new_n1014_));
  AND2_X1   g813(.A1(new_n961_), .A2(new_n997_), .ZN(new_n1015_));
  NAND2_X1  g814(.A1(new_n1015_), .A2(new_n701_), .ZN(new_n1016_));
  AOI21_X1  g815(.A(new_n1014_), .B1(new_n1016_), .B2(new_n1012_), .ZN(G1354gat));
  AOI21_X1  g816(.A(G218gat), .B1(new_n1015_), .B2(new_n708_), .ZN(new_n1018_));
  NAND2_X1  g817(.A1(new_n689_), .A2(G218gat), .ZN(new_n1019_));
  XOR2_X1   g818(.A(new_n1019_), .B(KEYINPUT127), .Z(new_n1020_));
  AOI21_X1  g819(.A(new_n1018_), .B1(new_n1015_), .B2(new_n1020_), .ZN(G1355gat));
endmodule


