//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n962_, new_n963_, new_n965_, new_n966_,
    new_n967_, new_n969_, new_n970_, new_n971_, new_n973_, new_n974_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT73), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(new_n204_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n203_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT36), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT74), .B1(new_n206_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT75), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n206_), .A2(new_n210_), .A3(KEYINPUT74), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n214_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT75), .B1(new_n216_), .B2(new_n211_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G85gat), .B(G92gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT7), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT6), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n219_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT65), .B(G92gat), .Z(new_n229_));
  INV_X1    g028(.A(G85gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232_));
  OAI22_X1  g031(.A1(new_n232_), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n232_), .B2(KEYINPUT9), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n228_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT6), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n222_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G106gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(KEYINPUT10), .B(G99gat), .Z(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n226_), .A2(new_n227_), .B1(new_n235_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT7), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n220_), .B(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(new_n237_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT66), .B1(new_n244_), .B2(new_n219_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n224_), .A2(new_n225_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(KEYINPUT8), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G29gat), .B(G36gat), .Z(new_n249_));
  XOR2_X1   g048(.A(G43gat), .B(G50gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT15), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT15), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n248_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT34), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n248_), .B2(new_n252_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n264_), .B(new_n261_), .C1(new_n248_), .C2(new_n252_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n259_), .A2(new_n260_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n265_), .B(new_n266_), .C1(new_n256_), .C2(new_n262_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n218_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n210_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n268_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT37), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT76), .ZN(new_n274_));
  INV_X1    g073(.A(new_n272_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT37), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n268_), .A2(new_n269_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n216_), .B2(new_n211_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n280_), .B(KEYINPUT37), .C1(new_n270_), .C2(new_n272_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n274_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G1gat), .ZN(new_n284_));
  INV_X1    g083(.A(G8gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT14), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT77), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(KEYINPUT77), .B(KEYINPUT14), .C1(new_n284_), .C2(new_n285_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G15gat), .B(G22gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G1gat), .B(G8gat), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n288_), .A2(new_n292_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G231gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G57gat), .B(G64gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n300_));
  XOR2_X1   g099(.A(G71gat), .B(G78gat), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n300_), .A2(new_n301_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n298_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G127gat), .B(G155gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G183gat), .B(G211gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT17), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n308_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT79), .Z(new_n317_));
  AND2_X1   g116(.A1(new_n313_), .A2(new_n314_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n308_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n283_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G230gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n241_), .A2(new_n306_), .A3(new_n247_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n241_), .A2(KEYINPUT67), .A3(new_n306_), .A4(new_n247_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n306_), .B1(new_n241_), .B2(new_n247_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n323_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n324_), .A2(new_n322_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT12), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n248_), .B2(new_n307_), .ZN(new_n333_));
  AOI211_X1 g132(.A(KEYINPUT12), .B(new_n306_), .C1(new_n241_), .C2(new_n247_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n331_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT69), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G120gat), .B(G148gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G176gat), .B(G204gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n336_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n330_), .A2(new_n335_), .A3(new_n342_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(KEYINPUT13), .ZN(new_n348_));
  XOR2_X1   g147(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n321_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n253_), .A2(new_n296_), .A3(new_n255_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n252_), .A2(new_n296_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G229gat), .A2(G233gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n356_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n251_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT80), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n357_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G113gat), .B(G141gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G169gat), .B(G197gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n362_), .A2(KEYINPUT81), .A3(new_n364_), .A4(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n357_), .A2(new_n360_), .A3(new_n367_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n367_), .B1(new_n361_), .B2(KEYINPUT80), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT81), .B1(new_n372_), .B2(new_n364_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT82), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n362_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n370_), .A4(new_n369_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n384_));
  INV_X1    g183(.A(G190gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT84), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G190gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n383_), .B(new_n384_), .C1(new_n389_), .C2(G183gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G169gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n383_), .A2(new_n384_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n389_), .B2(KEYINPUT26), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT25), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT83), .B1(new_n398_), .B2(G183gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n400_));
  INV_X1    g199(.A(G183gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT25), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(G183gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n395_), .B1(new_n397_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT24), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n407_), .A2(G169gat), .A3(G176gat), .ZN(new_n408_));
  INV_X1    g207(.A(G169gat), .ZN(new_n409_));
  INV_X1    g208(.A(G176gat), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT85), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n406_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n406_), .B1(G169gat), .B2(G176gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n409_), .A2(new_n410_), .A3(KEYINPUT85), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n407_), .B1(G169gat), .B2(G176gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n393_), .B1(new_n405_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(G71gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G99gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n418_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G127gat), .B(G134gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G120gat), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n424_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n424_), .A3(KEYINPUT87), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n422_), .B(new_n430_), .Z(new_n431_));
  XNOR2_X1  g230(.A(G15gat), .B(G43gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT86), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT30), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT31), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n431_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(G218gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G211gat), .ZN(new_n442_));
  INV_X1    g241(.A(G211gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G218gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT21), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G197gat), .B(G204gat), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G197gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G204gat), .ZN(new_n451_));
  INV_X1    g250(.A(G204gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G197gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n453_), .A3(KEYINPUT90), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT90), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(new_n450_), .A3(G204gat), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n454_), .A2(KEYINPUT91), .A3(KEYINPUT21), .A4(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n445_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n456_), .A2(KEYINPUT21), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT91), .B1(new_n460_), .B2(new_n454_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n449_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G183gat), .A2(G190gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n392_), .B1(new_n394_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n401_), .A2(KEYINPUT25), .ZN(new_n466_));
  AND2_X1   g265(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n466_), .B(new_n403_), .C1(new_n467_), .C2(new_n396_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n412_), .A2(new_n395_), .A3(new_n416_), .A4(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT95), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n467_), .A2(new_n396_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT25), .B(G183gat), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n394_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n474_), .A2(KEYINPUT95), .A3(new_n412_), .A4(new_n416_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n463_), .B1(new_n465_), .B2(new_n476_), .ZN(new_n477_));
  OR3_X1    g276(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n457_), .A2(new_n458_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n461_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT20), .B1(new_n418_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n440_), .B1(new_n477_), .B2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G8gat), .B(G36gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT18), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G64gat), .B(G92gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n463_), .A2(new_n476_), .A3(new_n465_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(new_n418_), .B2(new_n480_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n489_), .A3(new_n439_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n482_), .A2(new_n486_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT27), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n477_), .A2(new_n481_), .A3(new_n440_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n463_), .A2(new_n465_), .A3(new_n469_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n439_), .B1(new_n494_), .B2(new_n489_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT100), .B1(new_n493_), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(KEYINPUT100), .B2(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n486_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n492_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT24), .B1(new_n414_), .B2(new_n415_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n408_), .A2(new_n411_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(new_n413_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT95), .B1(new_n502_), .B2(new_n474_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n469_), .A2(new_n470_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n465_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n480_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n404_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n396_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT84), .B(G190gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT26), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n394_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n512_), .A2(new_n502_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n488_), .B1(new_n463_), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n439_), .B1(new_n506_), .B2(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n487_), .A2(new_n489_), .A3(new_n439_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n498_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT96), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n491_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT27), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n482_), .A2(new_n490_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(KEYINPUT96), .A3(new_n498_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT103), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT103), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n519_), .A2(new_n525_), .A3(new_n522_), .A4(new_n520_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n499_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G155gat), .A2(G162gat), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(G155gat), .A2(G162gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G141gat), .ZN(new_n534_));
  INV_X1    g333(.A(G148gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT3), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT3), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(G141gat), .B2(G148gat), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G141gat), .A2(G148gat), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT2), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT88), .B1(new_n539_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n536_), .A2(new_n538_), .ZN(new_n546_));
  AND3_X1   g345(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n546_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n533_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n531_), .B1(KEYINPUT1), .B2(new_n529_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n529_), .A2(KEYINPUT1), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(G141gat), .A2(G148gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n555_), .A2(new_n557_), .A3(new_n540_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n528_), .B1(new_n552_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT4), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n546_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n550_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n532_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n557_), .A3(new_n540_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(KEYINPUT89), .A3(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n559_), .A2(new_n560_), .A3(new_n565_), .A4(new_n430_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G225gat), .A2(G233gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n559_), .A2(new_n430_), .A3(new_n565_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT97), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n545_), .A2(new_n551_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n558_), .B1(new_n572_), .B2(new_n532_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n425_), .A2(new_n427_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n571_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n563_), .A2(new_n564_), .A3(new_n574_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT97), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n570_), .B(KEYINPUT4), .C1(new_n575_), .C2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n569_), .A2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n570_), .B(new_n567_), .C1(new_n575_), .C2(new_n577_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G1gat), .B(G29gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(G85gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT0), .B(G57gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(new_n584_));
  NAND4_X1  g383(.A1(new_n579_), .A2(KEYINPUT101), .A3(new_n580_), .A4(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n552_), .A2(new_n528_), .A3(new_n558_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT89), .B1(new_n563_), .B2(new_n564_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n576_), .A2(KEYINPUT97), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n573_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n588_), .A2(new_n430_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n578_), .A2(new_n569_), .B1(new_n591_), .B2(new_n567_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n585_), .B1(new_n592_), .B2(new_n584_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT101), .B1(new_n592_), .B2(new_n584_), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT102), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n579_), .A2(new_n580_), .A3(new_n584_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT101), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n579_), .A2(new_n580_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n584_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n598_), .A2(new_n601_), .A3(new_n602_), .A4(new_n585_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G228gat), .A2(G233gat), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT29), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT92), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n480_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT29), .B1(new_n552_), .B2(new_n558_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(KEYINPUT92), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n605_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G78gat), .B(G106gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n559_), .A2(KEYINPUT29), .A3(new_n565_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n463_), .A2(new_n605_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n559_), .A2(new_n565_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G22gat), .B(G50gat), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT28), .Z(new_n623_));
  AND3_X1   g422(.A1(new_n621_), .A2(new_n606_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n621_), .B2(new_n606_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n463_), .B1(new_n610_), .B2(KEYINPUT92), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n607_), .A2(new_n608_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n604_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n615_), .A2(new_n616_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n613_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n620_), .A2(new_n626_), .B1(new_n618_), .B2(new_n631_), .ZN(new_n632_));
  AND4_X1   g431(.A1(KEYINPUT93), .A2(new_n631_), .A3(new_n618_), .A4(new_n626_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n527_), .A2(new_n595_), .A3(new_n603_), .A4(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n634_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n486_), .A2(KEYINPUT32), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n521_), .B2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT32), .B(new_n486_), .C1(new_n521_), .C2(KEYINPUT99), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n639_), .B1(new_n497_), .B2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n641_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n578_), .A2(new_n567_), .A3(new_n566_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n591_), .A2(new_n568_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(new_n600_), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT98), .B(new_n584_), .C1(new_n591_), .C2(new_n568_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n519_), .A2(new_n522_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n592_), .A2(KEYINPUT33), .A3(new_n584_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT33), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n596_), .A2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .A4(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n642_), .A2(new_n653_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n635_), .A2(KEYINPUT104), .B1(new_n636_), .B2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n595_), .A2(new_n603_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n656_), .A2(new_n657_), .A3(new_n634_), .A4(new_n527_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n436_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n527_), .A2(new_n636_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n595_), .A2(new_n436_), .A3(new_n603_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n660_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n527_), .A2(new_n636_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n665_), .A2(KEYINPUT105), .A3(new_n662_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n380_), .B1(new_n659_), .B2(new_n667_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT106), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(KEYINPUT106), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n352_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n656_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n284_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT38), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n524_), .A2(new_n526_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n499_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n595_), .A2(new_n634_), .A3(new_n603_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT104), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n654_), .A2(new_n636_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n658_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n436_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT105), .B1(new_n665_), .B2(new_n662_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n661_), .A2(new_n660_), .A3(new_n663_), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n682_), .A2(new_n683_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n275_), .A2(new_n278_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n351_), .A2(new_n380_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n320_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G1gat), .B1(new_n692_), .B2(new_n656_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n673_), .A2(new_n674_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n675_), .A2(new_n693_), .A3(new_n694_), .ZN(G1324gat));
  NAND3_X1  g494(.A1(new_n671_), .A2(new_n285_), .A3(new_n678_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G8gat), .B1(new_n692_), .B2(new_n527_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT39), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT39), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g500(.A(G15gat), .B1(new_n692_), .B2(new_n683_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT41), .Z(new_n703_));
  INV_X1    g502(.A(new_n671_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n683_), .A2(G15gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(G1326gat));
  OAI21_X1  g505(.A(G22gat), .B1(new_n692_), .B2(new_n636_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT42), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n636_), .A2(G22gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n704_), .B2(new_n709_), .ZN(G1327gat));
  NOR2_X1   g509(.A1(new_n317_), .A2(new_n319_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n711_), .A2(new_n687_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n351_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G29gat), .B1(new_n714_), .B2(new_n672_), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n686_), .B2(new_n282_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n717_), .B(new_n283_), .C1(new_n659_), .C2(new_n667_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n690_), .A2(new_n711_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(KEYINPUT44), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT44), .B1(new_n719_), .B2(new_n720_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n672_), .A2(G29gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n715_), .B1(new_n723_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n527_), .A2(G36gat), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n714_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n714_), .B2(new_n728_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n721_), .A2(new_n722_), .A3(new_n527_), .ZN(new_n732_));
  INV_X1    g531(.A(G36gat), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n726_), .B1(new_n731_), .B2(new_n734_), .ZN(new_n735_));
  OAI221_X1 g534(.A(KEYINPUT46), .B1(new_n732_), .B2(new_n733_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1329gat));
  XNOR2_X1  g536(.A(KEYINPUT108), .B(G43gat), .ZN(new_n738_));
  INV_X1    g537(.A(new_n714_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n683_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n436_), .A2(G43gat), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n721_), .A2(new_n722_), .A3(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n743_), .A2(new_n741_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT47), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n743_), .A2(new_n741_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n743_), .A2(new_n741_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .A4(new_n740_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n750_), .ZN(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n714_), .B2(new_n634_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n634_), .A2(G50gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n723_), .B2(new_n753_), .ZN(G1331gat));
  INV_X1    g553(.A(new_n351_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n321_), .A2(new_n755_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT109), .Z(new_n757_));
  NOR2_X1   g556(.A1(new_n686_), .A2(new_n380_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G57gat), .B1(new_n759_), .B2(new_n672_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT110), .ZN(new_n761_));
  INV_X1    g560(.A(new_n380_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n689_), .A2(new_n762_), .A3(new_n755_), .A4(new_n711_), .ZN(new_n763_));
  XOR2_X1   g562(.A(KEYINPUT111), .B(G57gat), .Z(new_n764_));
  NOR3_X1   g563(.A1(new_n763_), .A2(new_n656_), .A3(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n761_), .A2(new_n765_), .ZN(G1332gat));
  OAI21_X1  g565(.A(G64gat), .B1(new_n763_), .B2(new_n527_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT48), .ZN(new_n768_));
  INV_X1    g567(.A(new_n759_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n527_), .A2(G64gat), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT112), .Z(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n769_), .B2(new_n771_), .ZN(G1333gat));
  OAI21_X1  g571(.A(G71gat), .B1(new_n763_), .B2(new_n683_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT49), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n683_), .A2(G71gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n769_), .B2(new_n775_), .ZN(G1334gat));
  OAI21_X1  g575(.A(G78gat), .B1(new_n763_), .B2(new_n636_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT50), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n636_), .A2(G78gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n769_), .B2(new_n779_), .ZN(G1335gat));
  NOR3_X1   g579(.A1(new_n351_), .A2(new_n711_), .A3(new_n687_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n758_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n230_), .A3(new_n672_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n351_), .A2(new_n380_), .A3(new_n711_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n787_), .A2(KEYINPUT113), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(KEYINPUT113), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n656_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n784_), .B1(new_n791_), .B2(new_n230_), .ZN(G1336gat));
  AOI21_X1  g591(.A(G92gat), .B1(new_n783_), .B2(new_n678_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n790_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n527_), .A2(new_n229_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(G1337gat));
  NAND2_X1  g595(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n436_), .A2(new_n239_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n782_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n790_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n436_), .B1(new_n800_), .B2(new_n788_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n801_), .B2(G99gat), .ZN(new_n802_));
  NOR2_X1   g601(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(G1338gat));
  NAND3_X1  g603(.A1(new_n783_), .A2(new_n238_), .A3(new_n634_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n636_), .B(new_n786_), .C1(new_n716_), .C2(new_n718_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n238_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n787_), .B2(new_n634_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n806_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n719_), .A2(new_n808_), .A3(new_n634_), .A4(new_n785_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(G106gat), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n814_), .A2(KEYINPUT52), .A3(new_n810_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n805_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT53), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n805_), .C1(new_n812_), .C2(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1339gat));
  NOR3_X1   g619(.A1(new_n665_), .A2(new_n656_), .A3(new_n683_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n353_), .A2(new_n355_), .A3(new_n358_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n356_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n368_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n370_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n345_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT118), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n345_), .A2(new_n826_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n326_), .B(new_n327_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n323_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n335_), .A2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n331_), .B(KEYINPUT55), .C1(new_n333_), .C2(new_n334_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n832_), .B1(new_n838_), .B2(new_n343_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n323_), .A2(new_n833_), .B1(new_n335_), .B2(new_n835_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n342_), .B1(new_n841_), .B2(new_n837_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n832_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n831_), .A2(new_n840_), .A3(new_n843_), .A4(KEYINPUT58), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT119), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n838_), .A2(new_n832_), .A3(new_n343_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n839_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(KEYINPUT58), .A4(new_n831_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n845_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT58), .B1(new_n847_), .B2(new_n831_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n282_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n838_), .A2(new_n343_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT117), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n856_), .A2(new_n832_), .B1(new_n839_), .B2(KEYINPUT117), .ZN(new_n857_));
  INV_X1    g656(.A(new_n345_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n859_));
  AOI22_X1  g658(.A1(new_n857_), .A2(new_n859_), .B1(new_n346_), .B2(new_n826_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n854_), .B1(new_n860_), .B2(new_n688_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n832_), .B1(new_n842_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n839_), .A2(KEYINPUT117), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n346_), .A2(new_n826_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT57), .A3(new_n687_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n853_), .A2(new_n861_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n853_), .A2(new_n861_), .A3(KEYINPUT120), .A4(new_n868_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n320_), .A3(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n762_), .A2(KEYINPUT116), .A3(new_n711_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n320_), .B2(new_n380_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n282_), .A2(new_n351_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n877_), .A2(new_n878_), .A3(KEYINPUT54), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n822_), .B1(new_n873_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(G113gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n380_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n867_), .A2(new_n687_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n854_), .A2(new_n889_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n711_), .B1(new_n890_), .B2(new_n868_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n888_), .B(new_n821_), .C1(new_n891_), .C2(new_n883_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n885_), .B2(new_n888_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n380_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n887_), .B1(new_n896_), .B2(new_n886_), .ZN(G1340gat));
  OAI211_X1 g696(.A(new_n755_), .B(new_n892_), .C1(new_n885_), .C2(new_n888_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT121), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n351_), .A2(G120gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n885_), .B1(KEYINPUT60), .B2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n711_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n883_), .B1(new_n902_), .B2(new_n872_), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT59), .B1(new_n903_), .B2(new_n822_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n904_), .A2(new_n905_), .A3(new_n755_), .A4(new_n892_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n899_), .A2(new_n901_), .A3(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G120gat), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n901_), .A2(KEYINPUT60), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1341gat));
  INV_X1    g709(.A(G127gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n885_), .A2(new_n911_), .A3(new_n711_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n894_), .A2(new_n711_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n914_), .B2(new_n911_), .ZN(G1342gat));
  OAI21_X1  g714(.A(G134gat), .B1(new_n893_), .B2(new_n282_), .ZN(new_n916_));
  INV_X1    g715(.A(G134gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n885_), .A2(new_n917_), .A3(new_n688_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n916_), .A2(KEYINPUT122), .A3(new_n918_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1343gat));
  NOR2_X1   g722(.A1(new_n903_), .A2(new_n436_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n924_), .A2(new_n672_), .A3(new_n634_), .A4(new_n527_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n762_), .ZN(new_n926_));
  XOR2_X1   g725(.A(KEYINPUT123), .B(G141gat), .Z(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1344gat));
  NOR2_X1   g727(.A1(new_n925_), .A2(new_n351_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(new_n535_), .ZN(G1345gat));
  NOR2_X1   g729(.A1(new_n925_), .A2(new_n320_), .ZN(new_n931_));
  XOR2_X1   g730(.A(KEYINPUT61), .B(G155gat), .Z(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1346gat));
  OAI21_X1  g732(.A(G162gat), .B1(new_n925_), .B2(new_n282_), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n687_), .A2(G162gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n925_), .B2(new_n935_), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n662_), .A2(new_n527_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n634_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n380_), .B(new_n939_), .C1(new_n891_), .C2(new_n883_), .ZN(new_n940_));
  XOR2_X1   g739(.A(KEYINPUT22), .B(G169gat), .Z(new_n941_));
  OR2_X1    g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n409_), .B1(new_n940_), .B2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n869_), .A2(new_n320_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n884_), .A2(new_n946_), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n947_), .A2(KEYINPUT124), .A3(new_n380_), .A4(new_n939_), .ZN(new_n948_));
  AND3_X1   g747(.A1(new_n944_), .A2(new_n945_), .A3(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n945_), .B1(new_n944_), .B2(new_n948_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n942_), .B1(new_n949_), .B2(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  OAI211_X1 g752(.A(KEYINPUT125), .B(new_n942_), .C1(new_n949_), .C2(new_n950_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1348gat));
  NAND2_X1  g754(.A1(new_n947_), .A2(new_n939_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(G176gat), .B1(new_n957_), .B2(new_n755_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n903_), .A2(new_n634_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n938_), .A2(new_n351_), .A3(new_n410_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n958_), .B1(new_n959_), .B2(new_n960_), .ZN(G1349gat));
  NOR3_X1   g760(.A1(new_n956_), .A2(new_n473_), .A3(new_n320_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n959_), .A2(new_n711_), .A3(new_n937_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n962_), .B1(new_n963_), .B2(new_n401_), .ZN(G1350gat));
  OAI21_X1  g763(.A(G190gat), .B1(new_n956_), .B2(new_n282_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n688_), .A2(new_n472_), .ZN(new_n966_));
  XOR2_X1   g765(.A(new_n966_), .B(KEYINPUT126), .Z(new_n967_));
  OAI21_X1  g766(.A(new_n965_), .B1(new_n956_), .B2(new_n967_), .ZN(G1351gat));
  NOR2_X1   g767(.A1(new_n679_), .A2(new_n527_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n924_), .A2(new_n969_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n970_), .A2(new_n762_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(new_n450_), .ZN(G1352gat));
  NOR2_X1   g771(.A1(new_n970_), .A2(new_n351_), .ZN(new_n973_));
  XOR2_X1   g772(.A(KEYINPUT127), .B(G204gat), .Z(new_n974_));
  XNOR2_X1  g773(.A(new_n973_), .B(new_n974_), .ZN(G1353gat));
  NAND3_X1  g774(.A1(new_n924_), .A2(new_n711_), .A3(new_n969_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  AND2_X1   g776(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n978_));
  NOR3_X1   g777(.A1(new_n976_), .A2(new_n977_), .A3(new_n978_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n979_), .B1(new_n976_), .B2(new_n977_), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n970_), .B2(new_n282_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n688_), .A2(new_n441_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n970_), .B2(new_n982_), .ZN(G1355gat));
endmodule


