//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT82), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G155gat), .A3(G162gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n211_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(KEYINPUT1), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT83), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n213_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n212_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT83), .B1(new_n219_), .B2(new_n214_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n207_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n214_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n215_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n203_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT84), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227_));
  OAI22_X1  g026(.A1(new_n205_), .A2(new_n227_), .B1(new_n203_), .B2(new_n224_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n223_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT85), .B1(new_n221_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n217_), .A3(new_n222_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n213_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n220_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n206_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT85), .ZN(new_n238_));
  INV_X1    g037(.A(new_n231_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT28), .B1(new_n241_), .B2(KEYINPUT29), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n232_), .A2(new_n240_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT28), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G22gat), .B(G50gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n242_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n248_), .B1(new_n242_), .B2(new_n246_), .ZN(new_n250_));
  INV_X1    g049(.A(G218gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G211gat), .ZN(new_n252_));
  INV_X1    g051(.A(G211gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G218gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n254_), .A3(KEYINPUT87), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT87), .B1(new_n252_), .B2(new_n254_), .ZN(new_n257_));
  INV_X1    g056(.A(G197gat), .ZN(new_n258_));
  INV_X1    g057(.A(G204gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G197gat), .A2(G204gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT21), .A3(new_n261_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n256_), .A2(new_n257_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  INV_X1    g063(.A(new_n261_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G197gat), .A2(G204gat), .ZN(new_n266_));
  OAI211_X1 g065(.A(KEYINPUT86), .B(new_n264_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n260_), .A2(new_n261_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT86), .B1(new_n269_), .B2(new_n264_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n262_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n257_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(new_n255_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n263_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G228gat), .A2(G233gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G78gat), .B(G106gat), .Z(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n245_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n277_), .B1(new_n282_), .B2(new_n275_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n279_), .A2(new_n281_), .A3(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n281_), .B1(new_n279_), .B2(new_n283_), .ZN(new_n285_));
  OR4_X1    g084(.A1(new_n249_), .A2(new_n250_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  OAI22_X1  g085(.A1(new_n249_), .A2(new_n250_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G127gat), .B(G134gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(G113gat), .B(G120gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n232_), .A2(new_n240_), .A3(new_n292_), .ZN(new_n293_));
  OR3_X1    g092(.A1(new_n221_), .A2(new_n231_), .A3(new_n292_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT91), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G57gat), .B(G85gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT94), .ZN(new_n300_));
  XOR2_X1   g099(.A(G1gat), .B(G29gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT92), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n293_), .A2(KEYINPUT4), .A3(new_n294_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n232_), .A2(new_n240_), .A3(new_n308_), .A4(new_n292_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n296_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n306_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n309_), .A2(new_n296_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n293_), .A2(KEYINPUT4), .A3(new_n294_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(KEYINPUT92), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n305_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n307_), .A2(new_n306_), .A3(new_n310_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT92), .B1(new_n312_), .B2(new_n313_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n298_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n304_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n315_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT19), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT25), .B(G183gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(KEYINPUT24), .A3(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n327_), .A2(KEYINPUT24), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n326_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT23), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(G183gat), .A3(G190gat), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT88), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n335_), .A2(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n334_), .A2(KEYINPUT78), .A3(G183gat), .A4(G190gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n333_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n342_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n344_), .A2(new_n345_), .B1(KEYINPUT23), .B2(new_n332_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n351_), .A2(KEYINPUT88), .A3(new_n348_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n341_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n337_), .B1(new_n353_), .B2(KEYINPUT89), .ZN(new_n354_));
  INV_X1    g153(.A(new_n341_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n347_), .A2(new_n342_), .A3(new_n349_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT88), .B1(new_n351_), .B2(new_n348_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT89), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n275_), .B1(new_n354_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n341_), .B1(new_n336_), .B2(new_n348_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n331_), .B2(new_n351_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(KEYINPUT79), .B(new_n362_), .C1(new_n331_), .C2(new_n351_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n275_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT20), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n323_), .B1(new_n361_), .B2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n275_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT20), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n323_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT90), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n353_), .A2(KEYINPUT89), .ZN(new_n375_));
  INV_X1    g174(.A(new_n337_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n375_), .A2(new_n360_), .A3(new_n275_), .A4(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n373_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n374_), .B1(new_n373_), .B2(new_n377_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n370_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT18), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n370_), .B(new_n384_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT27), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n376_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n353_), .A2(KEYINPUT89), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n368_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n369_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n323_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n367_), .A2(new_n368_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n353_), .A2(new_n275_), .A3(new_n376_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(KEYINPUT20), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n323_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n394_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n385_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n387_), .A2(new_n400_), .A3(KEYINPUT27), .ZN(new_n401_));
  NOR4_X1   g200(.A1(new_n289_), .A2(new_n321_), .A3(new_n388_), .A4(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT95), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n315_), .B2(KEYINPUT33), .ZN(new_n404_));
  INV_X1    g203(.A(new_n305_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT33), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(KEYINPUT95), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n313_), .A2(new_n297_), .A3(new_n309_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n293_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n319_), .A3(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n386_), .A2(new_n387_), .A3(new_n412_), .ZN(new_n413_));
  AOI211_X1 g212(.A(new_n407_), .B(new_n305_), .C1(new_n311_), .C2(new_n314_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT96), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT96), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n409_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n380_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n384_), .A2(KEYINPUT32), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n421_), .B(KEYINPUT97), .Z(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n420_), .A2(new_n422_), .B1(new_n399_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n321_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n417_), .A2(new_n419_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n402_), .B1(new_n426_), .B2(new_n289_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n367_), .B(KEYINPUT30), .ZN(new_n428_));
  INV_X1    g227(.A(G99gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT31), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G15gat), .B(G43gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(G71gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n434_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(new_n292_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n431_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n202_), .B1(new_n427_), .B2(new_n441_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n416_), .A2(KEYINPUT96), .B1(new_n321_), .B2(new_n424_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n288_), .B1(new_n443_), .B2(new_n419_), .ZN(new_n444_));
  OAI211_X1 g243(.A(KEYINPUT98), .B(new_n440_), .C1(new_n444_), .C2(new_n402_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT27), .ZN(new_n446_));
  INV_X1    g245(.A(new_n379_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n373_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n384_), .B1(new_n449_), .B2(new_n370_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n387_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n446_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n387_), .A2(new_n400_), .A3(KEYINPUT27), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT99), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT99), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n388_), .A2(new_n401_), .A3(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n289_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT100), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n289_), .B(KEYINPUT100), .C1(new_n454_), .C2(new_n456_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n459_), .A2(new_n320_), .A3(new_n441_), .A4(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT101), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n440_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n464_), .A2(KEYINPUT101), .A3(new_n320_), .A4(new_n460_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n442_), .A2(new_n445_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT75), .B(G8gat), .Z(new_n467_));
  INV_X1    g266(.A(G1gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT14), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G15gat), .B(G22gat), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G1gat), .B(G8gat), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n472_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G231gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G57gat), .B(G64gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT11), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT69), .ZN(new_n480_));
  XOR2_X1   g279(.A(G71gat), .B(G78gat), .Z(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(KEYINPUT11), .B2(new_n478_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n480_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n477_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G127gat), .B(G155gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT16), .ZN(new_n487_));
  XOR2_X1   g286(.A(G183gat), .B(G211gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT17), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n489_), .A2(new_n490_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n485_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n494_), .A2(KEYINPUT76), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(KEYINPUT76), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G190gat), .B(G218gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT72), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G134gat), .B(G162gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT36), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G232gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT34), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT35), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(KEYINPUT35), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n509_));
  INV_X1    g308(.A(G106gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n429_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n509_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT66), .ZN(new_n513_));
  NOR2_X1   g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT7), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(G85gat), .A2(G92gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n522_));
  OR2_X1    g321(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n516_), .A2(new_n521_), .A3(new_n522_), .A4(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n520_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n525_), .B1(new_n526_), .B2(KEYINPUT68), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(KEYINPUT68), .B2(new_n526_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT9), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n519_), .A2(KEYINPUT64), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT64), .B1(new_n519_), .B2(new_n530_), .ZN(new_n532_));
  OAI221_X1 g331(.A(new_n518_), .B1(new_n530_), .B2(new_n519_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT10), .B(G99gat), .Z(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n510_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n513_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n529_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G29gat), .B(G36gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n508_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n529_), .A2(new_n536_), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n540_), .B(KEYINPUT15), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n507_), .B1(new_n542_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n507_), .A3(new_n545_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n504_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n502_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(KEYINPUT36), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n547_), .A2(new_n552_), .A3(new_n548_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n498_), .B1(new_n554_), .B2(KEYINPUT37), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n547_), .A2(new_n552_), .A3(new_n548_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(new_n549_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT37), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(KEYINPUT74), .A3(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n503_), .B(KEYINPUT73), .ZN(new_n560_));
  INV_X1    g359(.A(new_n548_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n560_), .B1(new_n561_), .B2(new_n546_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n553_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n555_), .A2(new_n559_), .B1(KEYINPUT37), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n543_), .A2(new_n484_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n483_), .B1(new_n529_), .B2(new_n536_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT70), .B(new_n570_), .C1(new_n537_), .C2(new_n483_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n567_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT70), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT12), .B1(new_n568_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n569_), .B1(new_n575_), .B2(new_n566_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G120gat), .B(G148gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n576_), .B(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n583_), .A2(KEYINPUT13), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(KEYINPUT13), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n544_), .A2(new_n474_), .A3(new_n473_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n475_), .A2(new_n541_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n475_), .B(new_n541_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(new_n592_), .B2(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT77), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G169gat), .B(G197gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n594_), .B(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n586_), .A2(new_n598_), .ZN(new_n599_));
  NOR4_X1   g398(.A1(new_n466_), .A2(new_n497_), .A3(new_n564_), .A4(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n468_), .A3(new_n321_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT38), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n554_), .B(KEYINPUT102), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR4_X1   g404(.A1(new_n466_), .A2(new_n497_), .A3(new_n599_), .A4(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n468_), .B1(new_n606_), .B2(new_n321_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n602_), .B2(new_n601_), .ZN(G1324gat));
  NOR2_X1   g408(.A1(new_n454_), .A2(new_n456_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n600_), .A2(new_n467_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n606_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n610_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G8gat), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n614_), .A2(KEYINPUT39), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(KEYINPUT39), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n611_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT40), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(G1325gat));
  INV_X1    g418(.A(G15gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n600_), .A2(new_n620_), .A3(new_n441_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n606_), .A2(new_n441_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n622_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT41), .B1(new_n622_), .B2(G15gat), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n621_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT103), .Z(G1326gat));
  INV_X1    g425(.A(G22gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n627_), .B1(new_n606_), .B2(new_n288_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT42), .Z(new_n629_));
  NAND3_X1  g428(.A1(new_n600_), .A2(new_n627_), .A3(new_n288_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1327gat));
  INV_X1    g430(.A(new_n497_), .ZN(new_n632_));
  NOR4_X1   g431(.A1(new_n466_), .A2(new_n632_), .A3(new_n599_), .A4(new_n604_), .ZN(new_n633_));
  AOI21_X1  g432(.A(G29gat), .B1(new_n633_), .B2(new_n321_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n586_), .A2(new_n497_), .A3(new_n598_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n442_), .A2(new_n445_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n463_), .A2(new_n465_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n637_), .B1(new_n640_), .B2(new_n564_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n563_), .A2(KEYINPUT37), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n554_), .A2(new_n498_), .A3(KEYINPUT37), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT74), .B1(new_n557_), .B2(new_n558_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n466_), .A2(KEYINPUT43), .A3(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n636_), .B1(new_n641_), .B2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT44), .B1(new_n647_), .B2(KEYINPUT104), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n640_), .A2(new_n637_), .A3(new_n564_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT43), .B1(new_n466_), .B2(new_n645_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n635_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI22_X1  g452(.A1(new_n648_), .A2(new_n653_), .B1(KEYINPUT44), .B2(new_n651_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n321_), .A2(G29gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n634_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT107), .B1(new_n657_), .B2(KEYINPUT106), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n651_), .A2(KEYINPUT44), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n647_), .A2(KEYINPUT104), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n610_), .B(new_n660_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G36gat), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n613_), .A2(G36gat), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n633_), .A2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n668_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n633_), .A2(new_n666_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n657_), .A2(KEYINPUT107), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n659_), .B1(new_n665_), .B2(new_n675_), .ZN(new_n676_));
  AOI211_X1 g475(.A(new_n658_), .B(new_n674_), .C1(new_n664_), .C2(G36gat), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1329gat));
  INV_X1    g477(.A(KEYINPUT47), .ZN(new_n679_));
  INV_X1    g478(.A(G43gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n654_), .B2(new_n441_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n633_), .A2(new_n680_), .A3(new_n441_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n660_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G43gat), .B1(new_n685_), .B2(new_n440_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(KEYINPUT47), .A3(new_n682_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(G1330gat));
  AOI21_X1  g487(.A(G50gat), .B1(new_n633_), .B2(new_n288_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n288_), .A2(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n654_), .B2(new_n690_), .ZN(G1331gat));
  INV_X1    g490(.A(new_n586_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n497_), .A2(new_n598_), .ZN(new_n693_));
  AND4_X1   g492(.A1(new_n640_), .A2(new_n692_), .A3(new_n604_), .A4(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(G57gat), .A3(new_n321_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n696_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n466_), .A2(new_n586_), .A3(new_n598_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n564_), .A2(new_n497_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n320_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n697_), .B(new_n698_), .C1(G57gat), .C2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT109), .ZN(G1332gat));
  INV_X1    g503(.A(G64gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n694_), .B2(new_n610_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT48), .Z(new_n707_));
  INV_X1    g506(.A(new_n701_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n705_), .A3(new_n610_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1333gat));
  AOI21_X1  g509(.A(new_n436_), .B1(new_n694_), .B2(new_n441_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT49), .Z(new_n712_));
  NAND3_X1  g511(.A1(new_n708_), .A2(new_n436_), .A3(new_n441_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1334gat));
  INV_X1    g513(.A(G78gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n694_), .B2(new_n288_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n708_), .A2(new_n715_), .A3(new_n288_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1335gat));
  NAND2_X1  g519(.A1(new_n649_), .A2(new_n650_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n598_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n692_), .A2(new_n497_), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725_), .B2(new_n320_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n604_), .A2(new_n632_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n699_), .A2(new_n727_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n728_), .A2(G85gat), .A3(new_n320_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(G1336gat));
  OAI21_X1  g529(.A(G92gat), .B1(new_n725_), .B2(new_n613_), .ZN(new_n731_));
  OR3_X1    g530(.A1(new_n728_), .A2(G92gat), .A3(new_n613_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1337gat));
  OAI21_X1  g532(.A(G99gat), .B1(new_n725_), .B2(new_n440_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n441_), .A2(new_n534_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n728_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g536(.A1(new_n699_), .A2(new_n510_), .A3(new_n288_), .A4(new_n727_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n289_), .B(new_n723_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n510_), .B1(new_n740_), .B2(KEYINPUT111), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n723_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT111), .B1(new_n742_), .B2(new_n288_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n739_), .B1(new_n741_), .B2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n721_), .A2(KEYINPUT111), .A3(new_n288_), .A4(new_n724_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G106gat), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n743_), .A3(KEYINPUT52), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n738_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n738_), .C1(new_n745_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1339gat));
  XNOR2_X1  g552(.A(new_n693_), .B(KEYINPUT112), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n645_), .A3(new_n586_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT54), .Z(new_n756_));
  OR2_X1    g555(.A1(new_n576_), .A2(new_n582_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(new_n598_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT56), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(KEYINPUT113), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n575_), .B2(new_n566_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n575_), .A2(new_n566_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n575_), .A2(new_n762_), .A3(new_n566_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n582_), .B(new_n761_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n763_), .A2(new_n764_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n766_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n581_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n760_), .A2(KEYINPUT113), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT56), .B(new_n582_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(new_n759_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n758_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n593_), .A2(new_n597_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n589_), .B1(new_n475_), .B2(new_n541_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n591_), .A2(new_n589_), .B1(new_n587_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n778_), .B2(new_n597_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n583_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n605_), .B1(new_n775_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT57), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n773_), .A2(new_n759_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(new_n767_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n785_), .A2(new_n758_), .B1(new_n583_), .B2(new_n779_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n786_), .B2(new_n605_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n757_), .A2(new_n779_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n582_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n760_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n791_), .B2(new_n773_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n564_), .B(new_n788_), .C1(new_n792_), .C2(KEYINPUT58), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(KEYINPUT58), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n792_), .A2(KEYINPUT58), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n788_), .B1(new_n796_), .B2(new_n564_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n782_), .B(new_n787_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n756_), .B1(new_n798_), .B2(new_n497_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n464_), .A2(new_n321_), .A3(new_n460_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(G113gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n598_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT59), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n800_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n781_), .A2(KEYINPUT57), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n783_), .B(new_n605_), .C1(new_n775_), .C2(new_n780_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n796_), .A2(new_n564_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT115), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n793_), .A2(new_n794_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n632_), .B1(new_n809_), .B2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT59), .B(new_n806_), .C1(new_n814_), .C2(new_n756_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n805_), .A2(new_n815_), .A3(KEYINPUT116), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT116), .B1(new_n805_), .B2(new_n815_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n722_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n803_), .B1(new_n818_), .B2(new_n802_), .ZN(G1340gat));
  INV_X1    g618(.A(G120gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n586_), .B2(KEYINPUT60), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT117), .B1(new_n820_), .B2(KEYINPUT60), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n801_), .B(new_n823_), .C1(new_n824_), .C2(new_n821_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n586_), .B1(new_n805_), .B2(new_n815_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n820_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n801_), .B2(new_n632_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n816_), .A2(new_n817_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(G127gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n632_), .A2(KEYINPUT118), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(G127gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n828_), .B1(new_n829_), .B2(new_n833_), .ZN(G1342gat));
  INV_X1    g633(.A(G134gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n801_), .A2(new_n835_), .A3(new_n605_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n816_), .A2(new_n817_), .A3(new_n645_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n835_), .ZN(G1343gat));
  NAND3_X1  g637(.A1(new_n613_), .A2(new_n321_), .A3(new_n288_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n799_), .A2(new_n441_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n598_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n692_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT119), .B(G148gat), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1345gat));
  NAND2_X1  g644(.A1(new_n840_), .A2(new_n632_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT61), .B(G155gat), .Z(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n847_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n840_), .A2(new_n632_), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT120), .B(KEYINPUT121), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n848_), .A2(new_n852_), .A3(new_n850_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1346gat));
  AND3_X1   g655(.A1(new_n840_), .A2(G162gat), .A3(new_n564_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G162gat), .B1(new_n840_), .B2(new_n605_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n859_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n857_), .B1(new_n860_), .B2(new_n861_), .ZN(G1347gat));
  INV_X1    g661(.A(new_n799_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n613_), .A2(new_n321_), .A3(new_n440_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n598_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT123), .Z(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n289_), .A3(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n867_), .A2(new_n868_), .A3(G169gat), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n867_), .B2(G169gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n863_), .A2(new_n289_), .A3(new_n864_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT22), .B(G169gat), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n598_), .A2(new_n872_), .ZN(new_n873_));
  OAI22_X1  g672(.A1(new_n869_), .A2(new_n870_), .B1(new_n871_), .B2(new_n873_), .ZN(G1348gat));
  NOR2_X1   g673(.A1(new_n871_), .A2(new_n586_), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(G176gat), .Z(G1349gat));
  NOR2_X1   g675(.A1(new_n871_), .A2(new_n497_), .ZN(new_n877_));
  MUX2_X1   g676(.A(G183gat), .B(new_n324_), .S(new_n877_), .Z(G1350gat));
  OAI21_X1  g677(.A(G190gat), .B1(new_n871_), .B2(new_n645_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n605_), .A2(new_n325_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n871_), .B2(new_n880_), .ZN(G1351gat));
  NOR2_X1   g680(.A1(new_n799_), .A2(new_n441_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n613_), .A2(new_n321_), .A3(new_n289_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n722_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n258_), .ZN(G1352gat));
  AND3_X1   g685(.A1(new_n882_), .A2(new_n692_), .A3(new_n883_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT124), .B1(new_n887_), .B2(new_n259_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n889_), .B(G204gat), .C1(new_n884_), .C2(new_n586_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n882_), .A2(new_n259_), .A3(new_n692_), .A4(new_n883_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT125), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1353gat));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n253_), .A3(KEYINPUT126), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n895_), .B2(new_n253_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n884_), .A2(new_n497_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n898_), .B(new_n900_), .ZN(G1354gat));
  INV_X1    g700(.A(new_n884_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G218gat), .B1(new_n902_), .B2(new_n605_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n564_), .A2(G218gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT127), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n902_), .B2(new_n905_), .ZN(G1355gat));
endmodule


