//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT89), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n203_), .B(KEYINPUT89), .C1(G183gat), .C2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(KEYINPUT88), .A2(G169gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT87), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n209_), .B(KEYINPUT22), .C1(new_n210_), .C2(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n210_), .A2(KEYINPUT22), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n211_), .B(new_n212_), .C1(new_n209_), .C2(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .A4(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT85), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(new_n212_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n208_), .A3(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n218_), .B1(new_n219_), .B2(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n225_), .A2(KEYINPUT86), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n223_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n219_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n203_), .B(new_n228_), .C1(new_n225_), .C2(KEYINPUT86), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n215_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G15gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n230_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G71gat), .B(G99gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(G43gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT31), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(KEYINPUT91), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n237_), .B(new_n238_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(KEYINPUT91), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n236_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n233_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT90), .B(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT92), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n246_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G1gat), .B(G29gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G85gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT0), .B(G57gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(G155gat), .A3(G162gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT94), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G155gat), .ZN(new_n262_));
  INV_X1    g061(.A(G162gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT1), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT93), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT93), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(G155gat), .B2(G162gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n255_), .B(new_n257_), .C1(new_n261_), .C2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n267_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(G155gat), .B2(G162gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n256_), .B(KEYINPUT3), .Z(new_n272_));
  XOR2_X1   g071(.A(new_n255_), .B(KEYINPUT2), .Z(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n242_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n275_), .A2(new_n242_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n269_), .A2(new_n274_), .A3(new_n241_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(KEYINPUT4), .A3(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n280_), .A2(KEYINPUT103), .A3(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n282_), .A3(new_n278_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT103), .B1(new_n280_), .B2(new_n283_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n254_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT103), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n281_), .A2(KEYINPUT4), .A3(new_n282_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n277_), .A2(new_n279_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n292_), .A2(new_n284_), .A3(new_n253_), .A4(new_n285_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n249_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G197gat), .B(G204gat), .Z(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(KEYINPUT21), .ZN(new_n298_));
  XOR2_X1   g097(.A(G211gat), .B(G218gat), .Z(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G197gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT95), .A3(G204gat), .ZN(new_n302_));
  OAI211_X1 g101(.A(KEYINPUT21), .B(new_n302_), .C1(new_n297_), .C2(KEYINPUT95), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n297_), .A2(KEYINPUT21), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n300_), .A2(new_n303_), .B1(new_n299_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n230_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n308_));
  NOR2_X1   g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n203_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT100), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(KEYINPUT100), .A3(new_n203_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n224_), .A2(new_n308_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT98), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n216_), .B(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n318_), .B2(new_n217_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT22), .B(G169gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n212_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n208_), .B(KEYINPUT101), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n204_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(new_n305_), .A3(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n307_), .A2(KEYINPUT20), .A3(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n320_), .A2(new_n324_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n306_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n215_), .B(new_n305_), .C1(new_n226_), .C2(new_n229_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n329_), .B(KEYINPUT97), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n333_), .A2(KEYINPUT20), .A3(new_n334_), .A4(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G8gat), .B(G36gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(G64gat), .B(G92gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n335_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n324_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT20), .B1(new_n347_), .B2(new_n305_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n334_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n345_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n307_), .A2(KEYINPUT20), .A3(new_n325_), .A4(new_n329_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n342_), .A3(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n344_), .A2(KEYINPUT106), .A3(KEYINPUT27), .A4(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT27), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n350_), .A2(new_n342_), .A3(new_n351_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n342_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT107), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT28), .B1(new_n275_), .B2(KEYINPUT29), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n269_), .A2(new_n274_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n305_), .B1(new_n275_), .B2(KEYINPUT29), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n360_), .B(new_n363_), .C1(new_n367_), .C2(new_n305_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(G78gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G106gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G22gat), .B(G50gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n369_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n366_), .A2(new_n368_), .A3(new_n376_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT106), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n352_), .A2(KEYINPUT27), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n342_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n358_), .A2(new_n359_), .A3(new_n381_), .A4(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n353_), .A2(new_n385_), .A3(new_n381_), .A4(new_n357_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT107), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n296_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT105), .ZN(new_n390_));
  INV_X1    g189(.A(new_n356_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n283_), .A2(new_n278_), .A3(new_n277_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n281_), .A2(new_n282_), .A3(new_n279_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n254_), .A3(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n391_), .A2(new_n352_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT104), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n293_), .B(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n342_), .A2(KEYINPUT32), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n350_), .A2(new_n351_), .A3(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n348_), .A2(new_n349_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n402_), .A2(new_n335_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n403_), .B2(new_n400_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n395_), .A2(new_n399_), .B1(new_n405_), .B2(new_n294_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n390_), .B1(new_n406_), .B2(new_n380_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n355_), .A2(new_n356_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n284_), .A2(new_n285_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n409_), .A2(new_n253_), .A3(new_n292_), .A4(new_n398_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n293_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n411_));
  AND4_X1   g210(.A1(new_n408_), .A2(new_n410_), .A3(new_n394_), .A4(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n404_), .B1(new_n288_), .B2(new_n293_), .ZN(new_n413_));
  OAI211_X1 g212(.A(KEYINPUT105), .B(new_n381_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n288_), .A2(new_n380_), .A3(new_n293_), .ZN(new_n415_));
  AND4_X1   g214(.A1(new_n385_), .A2(new_n415_), .A3(new_n357_), .A4(new_n353_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n407_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n249_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n389_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT66), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G57gat), .B(G64gat), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(KEYINPUT11), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n422_), .A2(KEYINPUT11), .ZN(new_n425_));
  XOR2_X1   g224(.A(G71gat), .B(G78gat), .Z(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n421_), .A3(KEYINPUT11), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(KEYINPUT11), .B2(new_n422_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n427_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n429_), .B1(new_n430_), .B2(new_n423_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G15gat), .B(G22gat), .ZN(new_n433_));
  INV_X1    g232(.A(G1gat), .ZN(new_n434_));
  INV_X1    g233(.A(G8gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT14), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G1gat), .B(G8gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  XNOR2_X1  g238(.A(new_n432_), .B(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G231gat), .A2(G233gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G127gat), .B(G155gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G183gat), .B(G211gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(KEYINPUT17), .A3(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT79), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n447_), .B(KEYINPUT17), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT80), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n451_), .A2(new_n442_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n449_), .A2(KEYINPUT81), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT81), .B1(new_n449_), .B2(new_n452_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT65), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G85gat), .B(G92gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n458_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT8), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n457_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n458_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n464_), .A2(new_n466_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT7), .ZN(new_n473_));
  INV_X1    g272(.A(G99gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n373_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n459_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n471_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT64), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n462_), .A2(KEYINPUT64), .A3(new_n467_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n458_), .A2(KEYINPUT8), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n470_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G29gat), .B(G36gat), .Z(new_n485_));
  XOR2_X1   g284(.A(G43gat), .B(G50gat), .Z(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n471_), .A2(KEYINPUT9), .ZN(new_n489_));
  XOR2_X1   g288(.A(KEYINPUT10), .B(G99gat), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n373_), .ZN(new_n491_));
  INV_X1    g290(.A(G85gat), .ZN(new_n492_));
  INV_X1    g291(.A(G92gat), .ZN(new_n493_));
  OR3_X1    g292(.A1(new_n492_), .A2(new_n493_), .A3(KEYINPUT9), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n489_), .A2(new_n491_), .A3(new_n494_), .A4(new_n467_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n484_), .A2(new_n488_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G232gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT34), .ZN(new_n498_));
  INV_X1    g297(.A(new_n495_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT69), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n484_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n470_), .A2(new_n478_), .A3(new_n483_), .A4(KEYINPUT69), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n499_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n487_), .B(KEYINPUT15), .ZN(new_n504_));
  OAI221_X1 g303(.A(new_n496_), .B1(KEYINPUT35), .B2(new_n498_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(KEYINPUT35), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G190gat), .B(G218gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT74), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G134gat), .B(G162gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(KEYINPUT36), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT75), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n507_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(KEYINPUT36), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT76), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n507_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT37), .B1(new_n516_), .B2(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n507_), .A2(new_n518_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT37), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n515_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(KEYINPUT77), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT77), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(KEYINPUT37), .C1(new_n516_), .C2(new_n520_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n420_), .A2(new_n456_), .A3(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT5), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n484_), .A2(new_n432_), .A3(new_n495_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G230gat), .A2(G233gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT70), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n539_), .A3(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n501_), .A2(new_n502_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n495_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n432_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n484_), .A2(new_n495_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n432_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n544_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n541_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n535_), .A2(KEYINPUT67), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT67), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n484_), .A2(new_n553_), .A3(new_n432_), .A4(new_n495_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n549_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n556_));
  INV_X1    g355(.A(new_n536_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n556_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n551_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT71), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n534_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n551_), .B(KEYINPUT71), .C1(new_n558_), .C2(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT72), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n558_), .A2(new_n559_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n566_), .A2(KEYINPUT73), .A3(new_n551_), .A4(new_n534_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT73), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n560_), .B2(new_n533_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT72), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n562_), .A2(new_n571_), .A3(new_n563_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT13), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT83), .ZN(new_n577_));
  XOR2_X1   g376(.A(G169gat), .B(G197gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n504_), .A2(new_n439_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n488_), .B2(new_n439_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n488_), .A2(new_n439_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n488_), .A2(new_n439_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n580_), .A2(new_n583_), .B1(new_n586_), .B2(new_n582_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT82), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT84), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n579_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT82), .B1(new_n579_), .B2(new_n590_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n565_), .A2(KEYINPUT13), .A3(new_n570_), .A4(new_n572_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n575_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n529_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(new_n434_), .A3(new_n294_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT38), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n522_), .A2(new_n515_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n420_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT108), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n596_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n575_), .A2(KEYINPUT108), .A3(new_n594_), .A4(new_n595_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n604_), .A2(new_n608_), .A3(new_n456_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n609_), .A2(new_n294_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n600_), .B1(new_n434_), .B2(new_n610_), .ZN(G1324gat));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612_));
  INV_X1    g411(.A(new_n608_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n358_), .A2(new_n385_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n613_), .A2(new_n455_), .A3(new_n614_), .A4(new_n603_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT109), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n615_), .A2(new_n616_), .A3(G8gat), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n615_), .B2(G8gat), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n615_), .A2(G8gat), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(KEYINPUT109), .A3(new_n619_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n614_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(G8gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n598_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n612_), .B1(new_n620_), .B2(new_n626_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n618_), .A2(new_n619_), .B1(new_n598_), .B2(new_n624_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n618_), .A2(new_n619_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n628_), .B(KEYINPUT40), .C1(new_n629_), .C2(new_n617_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(G1325gat));
  INV_X1    g430(.A(G15gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n609_), .B2(new_n249_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT41), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n598_), .A2(new_n632_), .A3(new_n249_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1326gat));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n380_), .B(KEYINPUT110), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n637_), .B1(new_n609_), .B2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT42), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n598_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1327gat));
  NAND2_X1  g442(.A1(new_n456_), .A2(new_n602_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n420_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n597_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n646_), .A2(G29gat), .A3(new_n295_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  INV_X1    g448(.A(new_n528_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n420_), .B2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n381_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n416_), .B1(new_n652_), .B2(new_n390_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n249_), .B1(new_n653_), .B2(new_n414_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT43), .B(new_n528_), .C1(new_n654_), .C2(new_n389_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(new_n655_), .A3(new_n456_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n648_), .B1(new_n656_), .B2(new_n608_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n528_), .B1(new_n654_), .B2(new_n389_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n455_), .B1(new_n658_), .B2(new_n649_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n613_), .A2(new_n659_), .A3(KEYINPUT44), .A4(new_n655_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n660_), .A3(new_n294_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT111), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n661_), .A2(new_n662_), .A3(G29gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n661_), .B2(G29gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n647_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  NAND3_X1  g464(.A1(new_n657_), .A2(new_n660_), .A3(new_n614_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G36gat), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n623_), .A2(G36gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n645_), .A2(new_n597_), .A3(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT45), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT46), .B1(new_n671_), .B2(KEYINPUT112), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT112), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  AOI211_X1 g473(.A(new_n673_), .B(new_n674_), .C1(new_n667_), .C2(new_n670_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n672_), .A2(new_n675_), .ZN(G1329gat));
  NAND4_X1  g475(.A1(new_n657_), .A2(new_n660_), .A3(G43gat), .A4(new_n249_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n646_), .A2(new_n419_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(G43gat), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g479(.A1(new_n657_), .A2(new_n660_), .A3(G50gat), .A4(new_n380_), .ZN(new_n681_));
  INV_X1    g480(.A(G50gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n646_), .B2(new_n638_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1331gat));
  NAND2_X1  g483(.A1(new_n575_), .A2(new_n595_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n594_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n529_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G57gat), .B1(new_n688_), .B2(new_n294_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT113), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n690_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n687_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n693_), .A2(new_n604_), .A3(new_n456_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n294_), .A2(G57gat), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n691_), .A2(new_n692_), .B1(new_n694_), .B2(new_n695_), .ZN(G1332gat));
  INV_X1    g495(.A(G64gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n688_), .A2(new_n697_), .A3(new_n614_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n614_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G64gat), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(KEYINPUT48), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(KEYINPUT48), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(G1333gat));
  INV_X1    g502(.A(G71gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n688_), .A2(new_n704_), .A3(new_n249_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n694_), .A2(new_n249_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G71gat), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT49), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT49), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1334gat));
  NAND3_X1  g509(.A1(new_n688_), .A2(new_n371_), .A3(new_n639_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n687_), .A2(new_n455_), .A3(new_n603_), .A4(new_n639_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT50), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n712_), .A2(new_n713_), .A3(G78gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n712_), .B2(G78gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT114), .Z(G1335gat));
  NAND4_X1  g516(.A1(new_n687_), .A2(new_n651_), .A3(new_n456_), .A4(new_n655_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n295_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n687_), .A2(new_n645_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n492_), .A3(new_n294_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1336gat));
  OAI21_X1  g521(.A(G92gat), .B1(new_n718_), .B2(new_n623_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n493_), .A3(new_n614_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1337gat));
  NAND3_X1  g524(.A1(new_n720_), .A2(new_n490_), .A3(new_n249_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT115), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n718_), .A2(new_n419_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(G99gat), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n727_), .B(G99gat), .C1(new_n718_), .C2(new_n419_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n726_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(KEYINPUT116), .A3(KEYINPUT51), .ZN(new_n733_));
  NAND2_X1  g532(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n734_), .B(new_n726_), .C1(new_n729_), .C2(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1338gat));
  NAND3_X1  g535(.A1(new_n720_), .A2(new_n373_), .A3(new_n380_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n718_), .A2(new_n381_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G106gat), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n738_), .B(G106gat), .C1(new_n718_), .C2(new_n381_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n737_), .B1(new_n740_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT53), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n745_), .B(new_n737_), .C1(new_n740_), .C2(new_n742_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1339gat));
  NAND2_X1  g546(.A1(new_n587_), .A2(new_n579_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n580_), .A2(new_n585_), .A3(new_n582_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n579_), .B1(new_n586_), .B2(new_n581_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT119), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n750_), .A2(new_n751_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT120), .Z(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(new_n570_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n534_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n535_), .A2(new_n539_), .A3(new_n536_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n539_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n545_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n432_), .B1(new_n484_), .B2(new_n495_), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n503_), .A2(new_n763_), .B1(KEYINPUT12), .B2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT55), .B1(new_n762_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n541_), .A2(new_n546_), .A3(new_n767_), .A4(new_n550_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n552_), .A2(new_n554_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n546_), .A2(new_n771_), .A3(new_n550_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n772_), .B2(new_n557_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n552_), .A2(new_n554_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n770_), .B(new_n557_), .C1(new_n765_), .C2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n769_), .B1(new_n773_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT118), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n557_), .B1(new_n765_), .B2(new_n774_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT117), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n775_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(KEYINPUT118), .A3(new_n769_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n759_), .B1(new_n779_), .B2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n534_), .B1(new_n779_), .B2(new_n783_), .ZN(new_n785_));
  OAI22_X1  g584(.A1(KEYINPUT121), .A2(new_n784_), .B1(new_n785_), .B2(KEYINPUT56), .ZN(new_n786_));
  AOI221_X4 g585(.A(new_n778_), .B1(new_n766_), .B2(new_n768_), .C1(new_n781_), .C2(new_n775_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT118), .B1(new_n782_), .B2(new_n769_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n758_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n756_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n650_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n789_), .A2(new_n790_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n784_), .A2(KEYINPUT121), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n795_), .B(new_n796_), .C1(KEYINPUT56), .C2(new_n785_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT122), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(KEYINPUT58), .A4(new_n756_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT58), .B(new_n756_), .C1(new_n786_), .C2(new_n791_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT122), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n799_), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n789_), .B1(new_n785_), .B2(KEYINPUT56), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n570_), .A2(new_n594_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n803_), .A2(new_n805_), .B1(new_n573_), .B2(new_n755_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n602_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n573_), .A2(new_n755_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n533_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n779_), .A2(new_n783_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n810_), .A2(new_n757_), .B1(new_n811_), .B2(new_n758_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n809_), .B1(new_n812_), .B2(new_n804_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT57), .B1(new_n813_), .B2(new_n601_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n808_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n455_), .B1(new_n802_), .B2(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n528_), .A2(new_n456_), .A3(new_n594_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n686_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n816_), .A2(new_n820_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n295_), .B(new_n419_), .C1(new_n386_), .C2(new_n388_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n594_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT59), .B(new_n822_), .C1(new_n816_), .C2(new_n820_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n594_), .A2(G113gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT123), .Z(new_n831_));
  AOI21_X1  g630(.A(new_n825_), .B1(new_n829_), .B2(new_n831_), .ZN(G1340gat));
  XNOR2_X1  g631(.A(KEYINPUT124), .B(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n686_), .B2(KEYINPUT60), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n824_), .B(new_n834_), .C1(KEYINPUT60), .C2(new_n833_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n686_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n833_), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n824_), .A2(new_n838_), .A3(new_n455_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n456_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n838_), .ZN(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n824_), .A2(new_n842_), .A3(new_n602_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n650_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(G1343gat));
  OR2_X1    g644(.A1(new_n816_), .A2(new_n820_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n419_), .A2(new_n380_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n847_), .A2(new_n295_), .A3(new_n614_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n594_), .A3(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g649(.A1(new_n846_), .A2(new_n685_), .A3(new_n848_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g651(.A1(new_n846_), .A2(new_n455_), .A3(new_n848_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1346gat));
  OAI211_X1 g654(.A(new_n528_), .B(new_n848_), .C1(new_n816_), .C2(new_n820_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G162gat), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n601_), .A2(G162gat), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n848_), .B(new_n858_), .C1(new_n816_), .C2(new_n820_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n857_), .A2(KEYINPUT125), .A3(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n623_), .A2(new_n296_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n821_), .A2(new_n639_), .A3(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n594_), .A3(new_n321_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n865_), .A2(new_n594_), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n869_), .B(KEYINPUT126), .Z(new_n870_));
  OAI211_X1 g669(.A(new_n638_), .B(new_n870_), .C1(new_n816_), .C2(new_n820_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n871_), .A2(new_n872_), .A3(G169gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n871_), .B2(G169gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n868_), .B1(new_n873_), .B2(new_n874_), .ZN(G1348gat));
  NAND2_X1  g674(.A1(new_n867_), .A2(new_n685_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n821_), .A2(new_n380_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n686_), .A2(new_n212_), .A3(new_n866_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n876_), .A2(new_n212_), .B1(new_n877_), .B2(new_n878_), .ZN(G1349gat));
  NAND3_X1  g678(.A1(new_n877_), .A2(new_n455_), .A3(new_n865_), .ZN(new_n880_));
  INV_X1    g679(.A(G183gat), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n456_), .A2(new_n318_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n880_), .A2(new_n881_), .B1(new_n867_), .B2(new_n882_), .ZN(G1350gat));
  NOR2_X1   g682(.A1(new_n866_), .A2(new_n639_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n528_), .B(new_n884_), .C1(new_n816_), .C2(new_n820_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G190gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n602_), .A2(new_n217_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n884_), .B(new_n888_), .C1(new_n816_), .C2(new_n820_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT127), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT127), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n886_), .A2(new_n892_), .A3(new_n889_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1351gat));
  NOR3_X1   g693(.A1(new_n847_), .A2(new_n623_), .A3(new_n294_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n846_), .A2(new_n594_), .A3(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g696(.A1(new_n846_), .A2(new_n685_), .A3(new_n895_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g698(.A1(new_n846_), .A2(new_n455_), .A3(new_n895_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT63), .B(G211gat), .Z(new_n903_));
  NAND4_X1  g702(.A1(new_n846_), .A2(new_n455_), .A3(new_n895_), .A4(new_n903_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1354gat));
  NAND2_X1  g704(.A1(new_n846_), .A2(new_n895_), .ZN(new_n906_));
  OAI21_X1  g705(.A(G218gat), .B1(new_n906_), .B2(new_n650_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n601_), .A2(G218gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n906_), .B2(new_n908_), .ZN(G1355gat));
endmodule


