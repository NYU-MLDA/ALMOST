//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n202_), .B1(KEYINPUT11), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT11), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n205_), .B1(new_n203_), .B2(KEYINPUT11), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n204_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT66), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n211_), .A2(new_n212_), .A3(new_n202_), .A4(new_n206_), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  XOR2_X1   g014(.A(G85gat), .B(G92gat), .Z(new_n216_));
  NOR2_X1   g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT6), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n215_), .B(new_n216_), .C1(new_n219_), .C2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G85gat), .B(G92gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n219_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n221_), .A2(new_n223_), .A3(new_n228_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n227_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n226_), .B1(new_n232_), .B2(new_n215_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT9), .ZN(new_n234_));
  INV_X1    g033(.A(G85gat), .ZN(new_n235_));
  INV_X1    g034(.A(G92gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(new_n216_), .B2(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT64), .ZN(new_n239_));
  INV_X1    g038(.A(G106gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT10), .B(G99gat), .Z(new_n241_));
  AOI21_X1  g040(.A(new_n225_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n243_), .B(new_n237_), .C1(new_n216_), .C2(new_n234_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n239_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n214_), .B1(new_n233_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n224_), .A2(KEYINPUT65), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n217_), .B(KEYINPUT7), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(new_n231_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n215_), .B1(new_n249_), .B2(new_n216_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n226_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n245_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n209_), .A2(new_n213_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OR3_X1    g053(.A1(new_n246_), .A2(new_n254_), .A3(KEYINPUT67), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G230gat), .A2(G233gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n252_), .A2(KEYINPUT67), .A3(new_n253_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(KEYINPUT68), .A2(KEYINPUT12), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(new_n253_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n254_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n260_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(KEYINPUT68), .A2(KEYINPUT12), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n263_), .B1(new_n246_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n266_), .A3(new_n256_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G176gat), .B(G204gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT70), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G120gat), .B(G148gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n271_), .B(new_n272_), .Z(new_n273_));
  NAND3_X1  g072(.A1(new_n259_), .A2(new_n267_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n273_), .B1(new_n259_), .B2(new_n267_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n276_), .A2(new_n277_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT13), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G29gat), .B(G36gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G43gat), .B(G50gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT15), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n252_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G232gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT34), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT35), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n284_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n286_), .B(new_n291_), .C1(new_n292_), .C2(new_n252_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n289_), .A2(new_n290_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n294_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G190gat), .B(G218gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G134gat), .B(G162gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  OAI22_X1  g100(.A1(new_n297_), .A2(new_n298_), .B1(KEYINPUT36), .B2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(KEYINPUT36), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n295_), .A2(KEYINPUT72), .A3(new_n296_), .A4(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n301_), .A2(KEYINPUT36), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n297_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT37), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n309_), .A2(KEYINPUT73), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n309_), .A2(KEYINPUT73), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n308_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n302_), .A2(new_n304_), .B1(new_n297_), .B2(new_n306_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(KEYINPUT73), .A3(new_n309_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G15gat), .B(G22gat), .ZN(new_n318_));
  INV_X1    g117(.A(G1gat), .ZN(new_n319_));
  INV_X1    g118(.A(G8gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT14), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G8gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G231gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(new_n253_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G127gat), .B(G155gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT16), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G183gat), .B(G211gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT17), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n334_), .B(KEYINPUT74), .Z(new_n335_));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n331_), .B(new_n332_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n327_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n317_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n281_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT76), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT19), .ZN(new_n345_));
  INV_X1    g144(.A(G169gat), .ZN(new_n346_));
  INV_X1    g145(.A(G176gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT24), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  MUX2_X1   g148(.A(new_n348_), .B(KEYINPUT24), .S(new_n349_), .Z(new_n350_));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT23), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT26), .B(G190gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(KEYINPUT78), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT25), .B(G183gat), .ZN(new_n355_));
  INV_X1    g154(.A(G190gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT78), .B1(new_n356_), .B2(KEYINPUT26), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n350_), .B(new_n352_), .C1(new_n354_), .C2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G183gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n356_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n352_), .A2(new_n361_), .B1(G169gat), .B2(G176gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(KEYINPUT80), .A2(G169gat), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n363_), .B(KEYINPUT22), .C1(KEYINPUT79), .C2(G169gat), .ZN(new_n364_));
  AND2_X1   g163(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n364_), .B(new_n347_), .C1(new_n363_), .C2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n359_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT21), .ZN(new_n369_));
  INV_X1    g168(.A(G197gat), .ZN(new_n370_));
  INV_X1    g169(.A(G204gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT87), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT87), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G204gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n370_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G197gat), .A2(G204gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n369_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G218gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G211gat), .ZN(new_n379_));
  INV_X1    g178(.A(G211gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G218gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n372_), .A2(new_n374_), .A3(new_n370_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n369_), .B1(G197gat), .B2(G204gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n377_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n376_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT87), .B(G204gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n370_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n382_), .A2(KEYINPUT21), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT88), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n372_), .A2(new_n374_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n376_), .B1(new_n393_), .B2(G197gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n369_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT88), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n386_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n391_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(KEYINPUT88), .A3(new_n395_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n400_), .A2(new_n401_), .B1(new_n377_), .B2(new_n385_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT89), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n368_), .B1(new_n399_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT22), .B(G169gat), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n405_), .A2(KEYINPUT93), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(KEYINPUT93), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n347_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n353_), .A2(new_n355_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n409_), .A2(new_n352_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n408_), .A2(new_n362_), .B1(new_n410_), .B2(new_n350_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT20), .B1(new_n411_), .B2(new_n402_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n345_), .B1(new_n404_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT18), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n399_), .A2(new_n403_), .A3(new_n368_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n345_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT20), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n411_), .B2(new_n402_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n413_), .A2(new_n418_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT94), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n419_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n368_), .ZN(new_n427_));
  AOI221_X4 g226(.A(new_n398_), .B1(new_n377_), .B2(new_n385_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n400_), .A2(new_n401_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT89), .B1(new_n429_), .B2(new_n386_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n427_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n411_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n421_), .B1(new_n432_), .B2(new_n397_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n420_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n417_), .B1(new_n426_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT94), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n413_), .A2(new_n436_), .A3(new_n418_), .A4(new_n423_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n425_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT27), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n420_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT97), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n431_), .A2(new_n420_), .A3(new_n433_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n417_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n424_), .A2(KEYINPUT27), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n438_), .A2(new_n439_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G228gat), .A2(G233gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT86), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G155gat), .A2(G162gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT1), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT82), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT82), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT83), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n455_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n453_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G141gat), .ZN(new_n462_));
  INV_X1    g261(.A(G148gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G141gat), .A2(G148gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n458_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n456_), .A2(KEYINPUT83), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n454_), .A2(KEYINPUT82), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n455_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT3), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n465_), .A2(KEYINPUT84), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT2), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n476_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478_));
  OAI22_X1  g277(.A1(new_n478_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n475_), .A2(new_n477_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n473_), .A2(new_n451_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n467_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n450_), .B1(new_n483_), .B2(KEYINPUT29), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(new_n399_), .A3(new_n403_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n451_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n481_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n466_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n473_), .B2(new_n453_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT29), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n397_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n450_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n485_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G78gat), .B(G106gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n495_), .B(KEYINPUT90), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT91), .ZN(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(new_n483_), .B2(KEYINPUT29), .ZN(new_n501_));
  XOR2_X1   g300(.A(G22gat), .B(G50gat), .Z(new_n502_));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n503_));
  INV_X1    g302(.A(new_n500_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n467_), .A2(new_n482_), .A3(new_n503_), .A4(new_n504_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n501_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n502_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n485_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n498_), .A2(new_n499_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n428_), .A2(new_n430_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n511_), .A2(new_n484_), .B1(new_n450_), .B2(new_n492_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n501_), .A2(new_n505_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n502_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n501_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n496_), .B(new_n512_), .C1(new_n517_), .C2(KEYINPUT91), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n510_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n520_), .B1(new_n512_), .B2(new_n496_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n494_), .A2(KEYINPUT92), .A3(new_n497_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n508_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n519_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n448_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT98), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT4), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G127gat), .B(G134gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G113gat), .B(G120gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  OAI211_X1 g330(.A(KEYINPUT95), .B(new_n531_), .C1(new_n488_), .C2(new_n490_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n529_), .B(new_n530_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n467_), .A2(new_n482_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n528_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n467_), .B2(new_n482_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT4), .B1(new_n536_), .B2(KEYINPUT95), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G225gat), .A2(G233gat), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n535_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G1gat), .B(G29gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT96), .B(G85gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT0), .B(G57gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n534_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n538_), .B1(new_n545_), .B2(new_n536_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n539_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n544_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550_));
  AOI211_X1 g349(.A(new_n550_), .B(new_n533_), .C1(new_n467_), .C2(new_n482_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT4), .B1(new_n551_), .B2(new_n545_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n537_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n538_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n549_), .B1(new_n555_), .B2(new_n546_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n527_), .B1(new_n548_), .B2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n544_), .B1(new_n539_), .B2(new_n547_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n555_), .A2(new_n549_), .A3(new_n546_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(KEYINPUT98), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G227gat), .A2(G233gat), .ZN(new_n563_));
  INV_X1    g362(.A(G15gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(G71gat), .ZN(new_n566_));
  INV_X1    g365(.A(G99gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n427_), .A2(KEYINPUT30), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n427_), .A2(KEYINPUT30), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n568_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n568_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n569_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n531_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT81), .B(G43gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT31), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n572_), .A2(new_n575_), .A3(new_n533_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n577_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n526_), .A2(new_n562_), .A3(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n424_), .A2(KEYINPUT94), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n435_), .A2(new_n437_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n439_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n446_), .A2(new_n447_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n587_), .A2(new_n524_), .A3(new_n588_), .A4(new_n561_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n448_), .A2(KEYINPUT99), .A3(new_n524_), .A4(new_n561_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT33), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n558_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n556_), .A2(KEYINPUT33), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n538_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n545_), .A2(new_n536_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n596_), .B(new_n549_), .C1(new_n597_), .C2(new_n538_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n594_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n418_), .A2(KEYINPUT32), .ZN(new_n600_));
  INV_X1    g399(.A(new_n445_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n601_), .B2(new_n442_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n413_), .A2(new_n423_), .A3(new_n600_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n548_), .B2(new_n556_), .ZN(new_n604_));
  OAI22_X1  g403(.A1(new_n599_), .A2(new_n438_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n525_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n591_), .A2(new_n592_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n584_), .B1(new_n607_), .B2(new_n583_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n324_), .A2(new_n292_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G229gat), .A2(G233gat), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n285_), .A2(new_n324_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n324_), .B(new_n292_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n610_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n611_), .A2(new_n612_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G169gat), .B(G197gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n619_), .A2(KEYINPUT77), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(KEYINPUT77), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n615_), .A2(new_n618_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n608_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n343_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n561_), .A2(G1gat), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT100), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n627_), .A2(new_n631_), .A3(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n281_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n636_), .A2(new_n625_), .A3(new_n340_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n308_), .B(KEYINPUT101), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n608_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT102), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n637_), .A2(new_n642_), .A3(new_n639_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n561_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(new_n319_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n630_), .A2(KEYINPUT38), .A3(new_n632_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n635_), .A2(new_n645_), .A3(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(new_n448_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n627_), .A2(new_n320_), .A3(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n637_), .A2(new_n648_), .A3(new_n639_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(G8gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(new_n650_), .B2(G8gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n649_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(G1325gat));
  INV_X1    g456(.A(new_n583_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n627_), .A2(new_n564_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n641_), .A2(new_n643_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n564_), .B1(new_n660_), .B2(new_n658_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(KEYINPUT41), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(KEYINPUT41), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n627_), .A2(new_n665_), .A3(new_n524_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n525_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n665_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n667_), .A2(KEYINPUT42), .A3(new_n665_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n670_), .B2(new_n671_), .ZN(G1327gat));
  INV_X1    g471(.A(new_n340_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(new_n315_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n281_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n626_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n562_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679_));
  INV_X1    g478(.A(new_n317_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n608_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT104), .ZN(new_n682_));
  AOI22_X1  g481(.A1(new_n589_), .A2(new_n590_), .B1(new_n605_), .B2(new_n525_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n658_), .B1(new_n683_), .B2(new_n592_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n317_), .B1(new_n684_), .B2(new_n584_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT43), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n682_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n681_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n636_), .A2(new_n625_), .A3(new_n673_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n688_), .A2(KEYINPUT44), .A3(new_n689_), .A4(new_n690_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n691_), .A2(G29gat), .A3(new_n562_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n678_), .B1(new_n692_), .B2(new_n695_), .ZN(G1328gat));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n691_), .A2(new_n648_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n695_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n648_), .A2(KEYINPUT105), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n648_), .A2(KEYINPUT105), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n698_), .ZN(new_n704_));
  OR3_X1    g503(.A1(new_n676_), .A2(KEYINPUT45), .A3(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT45), .B1(new_n676_), .B2(new_n704_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n697_), .B1(new_n700_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n695_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n691_), .A2(new_n648_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G36gat), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(KEYINPUT46), .A3(new_n707_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n709_), .A2(new_n713_), .ZN(G1329gat));
  NAND3_X1  g513(.A1(new_n691_), .A2(G43gat), .A3(new_n658_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n676_), .A2(new_n583_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT106), .B(G43gat), .ZN(new_n717_));
  OAI22_X1  g516(.A1(new_n710_), .A2(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT47), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720_));
  OAI221_X1 g519(.A(new_n720_), .B1(new_n716_), .B2(new_n717_), .C1(new_n710_), .C2(new_n715_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1330gat));
  AOI21_X1  g521(.A(G50gat), .B1(new_n677_), .B2(new_n524_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n691_), .A2(G50gat), .A3(new_n524_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n695_), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n281_), .A2(new_n624_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n608_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n341_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n562_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n281_), .A2(new_n624_), .A3(new_n340_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(new_n639_), .ZN(new_n731_));
  INV_X1    g530(.A(G57gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n562_), .B2(KEYINPUT107), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(KEYINPUT107), .B2(new_n732_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n729_), .B1(new_n731_), .B2(new_n734_), .ZN(G1332gat));
  INV_X1    g534(.A(G64gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n731_), .B2(new_n703_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT48), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n728_), .A2(new_n736_), .A3(new_n703_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n728_), .A2(new_n741_), .A3(new_n658_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n731_), .A2(new_n658_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT49), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(G71gat), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n743_), .B2(G71gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n742_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(G1334gat));
  INV_X1    g549(.A(G78gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n731_), .B2(new_n524_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT50), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n728_), .A2(new_n751_), .A3(new_n524_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1335gat));
  NAND2_X1  g554(.A1(new_n562_), .A2(G85gat), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT111), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n281_), .A2(new_n624_), .A3(new_n673_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n686_), .B1(new_n608_), .B2(new_n680_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n686_), .B1(new_n685_), .B2(new_n679_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n689_), .B(new_n759_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n688_), .A2(KEYINPUT110), .A3(new_n689_), .A4(new_n759_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n758_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n726_), .A2(new_n727_), .A3(new_n674_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n562_), .ZN(new_n773_));
  OR3_X1    g572(.A1(new_n768_), .A2(new_n769_), .A3(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n769_), .B1(new_n768_), .B2(new_n773_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1336gat));
  NAND3_X1  g575(.A1(new_n772_), .A2(new_n236_), .A3(new_n648_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n703_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n779_), .B2(new_n236_), .ZN(G1337gat));
  NAND3_X1  g579(.A1(new_n772_), .A2(new_n658_), .A3(new_n241_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n583_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(new_n567_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n781_), .B(new_n784_), .C1(new_n782_), .C2(new_n567_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n772_), .A2(new_n240_), .A3(new_n524_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n688_), .A2(new_n524_), .A3(new_n689_), .A4(new_n759_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(G106gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(G106gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n789_), .B(new_n795_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1339gat));
  NAND3_X1  g598(.A1(new_n233_), .A2(new_n214_), .A3(new_n245_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n246_), .B2(new_n263_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n260_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n257_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT115), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n267_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n262_), .A2(new_n266_), .A3(KEYINPUT55), .A4(new_n256_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n808_), .B(new_n257_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n804_), .A2(new_n806_), .A3(new_n807_), .A4(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n273_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n811_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AOI211_X1 g614(.A(KEYINPUT116), .B(KEYINPUT56), .C1(new_n810_), .C2(new_n811_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n812_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n624_), .A2(new_n274_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n612_), .A2(new_n609_), .A3(new_n614_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n618_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n613_), .A2(new_n610_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT117), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n278_), .A2(new_n279_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n308_), .B1(new_n819_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n813_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n812_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n825_), .A2(new_n274_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT58), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n680_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n812_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n832_), .B(KEYINPUT58), .C1(new_n835_), .C2(new_n813_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n831_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n832_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n829_), .A2(KEYINPUT57), .B1(new_n834_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n827_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n308_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n340_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n281_), .A2(new_n341_), .A3(new_n625_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n658_), .A2(new_n562_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n526_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(KEYINPUT59), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n844_), .A2(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT118), .B(new_n842_), .C1(new_n843_), .C2(new_n308_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n841_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n849_), .B1(new_n860_), .B2(new_n340_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n854_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n624_), .B(new_n856_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G113gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n340_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n850_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n853_), .ZN(new_n868_));
  OR3_X1    g667(.A1(new_n868_), .A2(G113gat), .A3(new_n625_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n865_), .A2(new_n869_), .ZN(G1340gat));
  OAI211_X1 g669(.A(new_n636_), .B(new_n856_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G120gat), .ZN(new_n872_));
  INV_X1    g671(.A(G120gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n281_), .B2(KEYINPUT60), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n862_), .B(new_n874_), .C1(KEYINPUT60), .C2(new_n873_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(G1341gat));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n861_), .A2(new_n340_), .A3(new_n854_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(G127gat), .ZN(new_n879_));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT120), .B(new_n880_), .C1(new_n868_), .C2(new_n340_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n868_), .A2(KEYINPUT59), .B1(new_n851_), .B2(new_n855_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n340_), .A2(new_n880_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n879_), .A2(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(G1342gat));
  INV_X1    g683(.A(new_n638_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n861_), .A2(new_n885_), .A3(new_n854_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT121), .B1(new_n886_), .B2(G134gat), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888_));
  INV_X1    g687(.A(G134gat), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n888_), .B(new_n889_), .C1(new_n868_), .C2(new_n885_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n317_), .A2(G134gat), .ZN(new_n891_));
  XOR2_X1   g690(.A(new_n891_), .B(KEYINPUT122), .Z(new_n892_));
  AOI22_X1  g691(.A1(new_n887_), .A2(new_n890_), .B1(new_n882_), .B2(new_n892_), .ZN(G1343gat));
  NOR4_X1   g692(.A1(new_n703_), .A2(new_n525_), .A3(new_n561_), .A4(new_n658_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT123), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n866_), .B2(new_n850_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n624_), .ZN(new_n897_));
  XOR2_X1   g696(.A(KEYINPUT124), .B(G141gat), .Z(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n636_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g700(.A1(new_n896_), .A2(new_n673_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  INV_X1    g703(.A(G162gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n896_), .B2(new_n317_), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n861_), .A2(G162gat), .A3(new_n895_), .A4(new_n885_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT125), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n896_), .A2(new_n905_), .A3(new_n638_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n861_), .A2(new_n680_), .A3(new_n895_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n909_), .B(new_n910_), .C1(new_n911_), .C2(new_n905_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n912_), .ZN(G1347gat));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n778_), .A2(new_n562_), .A3(new_n583_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n525_), .ZN(new_n916_));
  AOI211_X1 g715(.A(new_n625_), .B(new_n916_), .C1(new_n846_), .C2(new_n850_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n914_), .B1(new_n917_), .B2(new_n346_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n916_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n851_), .A2(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(KEYINPUT62), .B(G169gat), .C1(new_n921_), .C2(new_n625_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n918_), .A2(new_n919_), .A3(new_n922_), .ZN(G1348gat));
  OAI21_X1  g722(.A(new_n347_), .B1(new_n921_), .B2(new_n281_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n861_), .A2(new_n524_), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n915_), .A2(G176gat), .A3(new_n636_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n924_), .A2(new_n925_), .A3(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n916_), .B1(new_n846_), .B2(new_n850_), .ZN(new_n930_));
  AOI21_X1  g729(.A(G176gat), .B1(new_n930_), .B2(new_n636_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n867_), .A2(new_n525_), .A3(new_n927_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT126), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n929_), .A2(new_n933_), .ZN(G1349gat));
  NOR3_X1   g733(.A1(new_n921_), .A2(new_n355_), .A3(new_n340_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n926_), .A2(new_n673_), .A3(new_n915_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n360_), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n921_), .B2(new_n680_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n930_), .A2(new_n353_), .A3(new_n638_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1351gat));
  NOR4_X1   g739(.A1(new_n778_), .A2(new_n525_), .A3(new_n562_), .A4(new_n658_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n861_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n624_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g744(.A1(new_n867_), .A2(new_n941_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n946_), .A2(new_n388_), .A3(new_n281_), .ZN(new_n947_));
  AOI21_X1  g746(.A(G204gat), .B1(new_n943_), .B2(new_n636_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1353gat));
  NOR2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n340_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n867_), .A2(new_n941_), .A3(new_n951_), .A4(new_n952_), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n953_), .A2(KEYINPUT127), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n953_), .A2(KEYINPUT127), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n951_), .B1(new_n943_), .B2(new_n952_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n954_), .A2(new_n955_), .A3(new_n956_), .ZN(G1354gat));
  OAI21_X1  g756(.A(G218gat), .B1(new_n946_), .B2(new_n680_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n943_), .A2(new_n378_), .A3(new_n638_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1355gat));
endmodule


